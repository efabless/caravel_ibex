* NGSPICE file created from DMC_32x16HC.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_2 abstract view
.subckt sky130_fd_sc_hd__ebufn_2 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlclkp_1 abstract view
.subckt sky130_fd_sc_hd__dlclkp_1 CLK GATE VGND VNB VPB VPWR GCLK
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_4 abstract view
.subckt sky130_fd_sc_hd__nor4b_4 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

.subckt DMC_32x16HC A[0] A[10] A[11] A[12] A[13] A[14] A[15] A[16] A[17] A[18] A[19]
+ A[1] A[20] A[21] A[2] A[3] A[4] A[5] A[6] A[7] A[8] A[9] A_h[0] A_h[10] A_h[11]
+ A_h[12] A_h[13] A_h[14] A_h[15] A_h[16] A_h[17] A_h[18] A_h[19] A_h[1] A_h[2] A_h[3]
+ A_h[4] A_h[5] A_h[6] A_h[7] A_h[8] A_h[9] Do[0] Do[10] Do[11] Do[12] Do[13] Do[14]
+ Do[15] Do[16] Do[17] Do[18] Do[19] Do[1] Do[20] Do[21] Do[22] Do[23] Do[24] Do[25]
+ Do[26] Do[27] Do[28] Do[29] Do[2] Do[30] Do[31] Do[3] Do[4] Do[5] Do[6] Do[7] Do[8]
+ Do[9] clk hit line[0] line[100] line[101] line[102] line[103] line[104] line[105]
+ line[106] line[107] line[108] line[109] line[10] line[110] line[111] line[112] line[113]
+ line[114] line[115] line[116] line[117] line[118] line[119] line[11] line[120] line[121]
+ line[122] line[123] line[124] line[125] line[126] line[127] line[12] line[13] line[14]
+ line[15] line[16] line[17] line[18] line[19] line[1] line[20] line[21] line[22]
+ line[23] line[24] line[25] line[26] line[27] line[28] line[29] line[2] line[30]
+ line[31] line[32] line[33] line[34] line[35] line[36] line[37] line[38] line[39]
+ line[3] line[40] line[41] line[42] line[43] line[44] line[45] line[46] line[47]
+ line[48] line[49] line[4] line[50] line[51] line[52] line[53] line[54] line[55]
+ line[56] line[57] line[58] line[59] line[5] line[60] line[61] line[62] line[63]
+ line[64] line[65] line[66] line[67] line[68] line[69] line[6] line[70] line[71]
+ line[72] line[73] line[74] line[75] line[76] line[77] line[78] line[79] line[7]
+ line[80] line[81] line[82] line[83] line[84] line[85] line[86] line[87] line[88]
+ line[89] line[8] line[90] line[91] line[92] line[93] line[94] line[95] line[96]
+ line[97] line[98] line[99] line[9] rst_n wr vccd1 vssd1
XOVHB\[16\].VALID\[10\].TOBUF OVHB\[16\].VALID\[10\].FF/Q OVHB\[16\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04932_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__09515__D line[41] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05903_ _05903_/A _05914_/Y vssd1 vssd1 vccd1 vccd1 _13743_/Z sky130_fd_sc_hd__ebufn_2
X_09671_ _09671_/A _09694_/Y vssd1 vssd1 vccd1 vccd1 _13871_/Z sky130_fd_sc_hd__ebufn_2
X_06883_ _06883_/A _06894_/Y vssd1 vssd1 vccd1 vccd1 _13883_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_94_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08622_ _08640_/CLK line[31] vssd1 vssd1 vccd1 vccd1 _08623_/A sky130_fd_sc_hd__dfxtp_1
X_05834_ _05840_/CLK line[22] vssd1 vssd1 vccd1 vccd1 _05835_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.M\[1\].MUX\[1\]_A1 _13716_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07035__D line[64] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08553_ _08553_/A _08574_/Y vssd1 vssd1 vccd1 vccd1 _13873_/Z sky130_fd_sc_hd__ebufn_2
X_05765_ _05765_/A _05774_/Y vssd1 vssd1 vccd1 vccd1 _13885_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11780__D line[52] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06874__D line[113] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07504_ _07520_/CLK line[17] vssd1 vssd1 vccd1 vccd1 _07505_/A sky130_fd_sc_hd__dfxtp_1
X_08484_ _08500_/CLK line[81] vssd1 vssd1 vccd1 vccd1 _08485_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05696_ _05700_/CLK line[87] vssd1 vssd1 vccd1 vccd1 _05697_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06229__A _13903_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09250__D line[62] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07435_ _07435_/A _07454_/Y vssd1 vssd1 vccd1 vccd1 _13875_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_22_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07366_ _07380_/CLK line[82] vssd1 vssd1 vccd1 vccd1 _07367_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[9\].VALID\[9\].FF_D A[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06317_ _06317_/A _06334_/Y vssd1 vssd1 vccd1 vccd1 _13877_/Z sky130_fd_sc_hd__ebufn_2
X_09105_ _09105_/A _09134_/Y vssd1 vssd1 vccd1 vccd1 _13865_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_148_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07297_ _07297_/A _07314_/Y vssd1 vssd1 vccd1 vccd1 _13737_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_136_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09036_ _09060_/CLK line[92] vssd1 vssd1 vccd1 vccd1 _09037_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_108_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06248_ _06260_/CLK line[83] vssd1 vssd1 vccd1 vccd1 _06249_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_184_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12116__D line[92] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06179_ _06179_/A _06194_/Y vssd1 vssd1 vccd1 vccd1 _13739_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[27\].CLKBUF\[2\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11020__D line[89] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06114__D line[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11955__D line[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__04929__A1_N A_h[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09938_ _13921_/X wr vssd1 vssd1 vccd1 vccd1 _09938_/X sky130_fd_sc_hd__and2_1
XFILLER_77_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09425__D line[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09869_ _13921_/X vssd1 vssd1 vccd1 vccd1 _09869_/Y sky130_fd_sc_hd__inv_2
X_11900_ _11930_/CLK line[112] vssd1 vssd1 vccd1 vccd1 _11901_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_45_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12880_ _12910_/CLK line[48] vssd1 vssd1 vccd1 vccd1 _12881_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_172_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07523__A _13911_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11831_ _11831_/A _11864_/Y vssd1 vssd1 vccd1 vccd1 _13791_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_45_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11690__D line[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11762_ _11790_/CLK line[58] vssd1 vssd1 vccd1 vccd1 _11763_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13501_ _13505_/CLK line[71] vssd1 vssd1 vccd1 vccd1 _13502_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10713_ _10713_/A _10744_/Y vssd1 vssd1 vccd1 vccd1 _13793_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_159_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[9\].VALID\[11\].FF_D A[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10884__A _13925_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11693_ _11693_/A _11724_/Y vssd1 vssd1 vccd1 vccd1 _13653_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13432_ _13432_/A _13439_/Y vssd1 vssd1 vccd1 vccd1 _13712_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10644_ _10670_/CLK line[59] vssd1 vssd1 vccd1 vccd1 _10645_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13363_ _13365_/CLK line[8] vssd1 vssd1 vccd1 vccd1 _13364_/A sky130_fd_sc_hd__dfxtp_1
X_10575_ _10575_/A _10604_/Y vssd1 vssd1 vccd1 vccd1 _13655_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_154_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12314_ _12314_/A _12319_/Y vssd1 vssd1 vccd1 vccd1 _13714_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_127_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13294_ _13294_/A _13299_/Y vssd1 vssd1 vccd1 vccd1 _13854_/Z sky130_fd_sc_hd__ebufn_2
X_12245_ _12245_/CLK line[9] vssd1 vssd1 vccd1 vccd1 _12246_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06024__D line[123] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12176_ _12176_/A _12179_/Y vssd1 vssd1 vccd1 vccd1 _13856_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_96_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11865__D line[96] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_DATA\[0\].CLKBUF\[1\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11127_ _11127_/CLK _11128_/X vssd1 vssd1 vccd1 vccd1 _11125_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_49_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05863__D line[35] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11058_ _13925_/X wr vssd1 vssd1 vccd1 vccd1 _11058_/X sky130_fd_sc_hd__and2_1
XFILLER_92_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10009_ _13922_/X vssd1 vssd1 vccd1 vccd1 _10009_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10778__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12696__D line[87] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XOVHB\[22\].CGAND _13915_/X wr vssd1 vssd1 vccd1 vccd1 OVHB\[22\].CGAND/X sky130_fd_sc_hd__and2_4
X_05550_ _05560_/CLK line[20] vssd1 vssd1 vccd1 vccd1 _05551_/A sky130_fd_sc_hd__dfxtp_1
X_05481_ _05481_/A _05494_/Y vssd1 vssd1 vccd1 vccd1 _13881_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_60_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11105__D line[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07220_ _07240_/CLK line[30] vssd1 vssd1 vccd1 vccd1 _07221_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_20_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05103__D line[72] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07151_ _07151_/A _07174_/Y vssd1 vssd1 vccd1 vccd1 _13871_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10944__D line[54] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13320__D line[116] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06102_ _06120_/CLK line[31] vssd1 vssd1 vccd1 vccd1 _06103_/A sky130_fd_sc_hd__dfxtp_1
X_07082_ _07100_/CLK line[95] vssd1 vssd1 vccd1 vccd1 _07083_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08414__D line[49] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06033_ _06033_/A _06054_/Y vssd1 vssd1 vccd1 vccd1 _13873_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[18\].VALID\[4\].TOBUF OVHB\[18\].VALID\[4\].FF/Q OVHB\[18\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04925_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_114_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07984_ _08010_/CLK line[123] vssd1 vssd1 vccd1 vccd1 _07985_/A sky130_fd_sc_hd__dfxtp_1
X_09723_ _09725_/CLK line[8] vssd1 vssd1 vccd1 vccd1 _09724_/A sky130_fd_sc_hd__dfxtp_1
X_06935_ _06935_/A _06964_/Y vssd1 vssd1 vccd1 vccd1 _13655_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_95_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09654_ _09654_/A _09659_/Y vssd1 vssd1 vccd1 vccd1 _13854_/Z sky130_fd_sc_hd__ebufn_2
X_06866_ _06890_/CLK line[124] vssd1 vssd1 vccd1 vccd1 _06867_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_55_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08605_ _08605_/CLK line[9] vssd1 vssd1 vccd1 vccd1 _08606_/A sky130_fd_sc_hd__dfxtp_1
X_05817_ _05817_/A _05844_/Y vssd1 vssd1 vccd1 vccd1 _13657_/Z sky130_fd_sc_hd__ebufn_2
X_09585_ _09585_/CLK line[73] vssd1 vssd1 vccd1 vccd1 _09586_/A sky130_fd_sc_hd__dfxtp_1
X_06797_ _06797_/A _06824_/Y vssd1 vssd1 vccd1 vccd1 _13797_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_63_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08536_ _08536_/A _08539_/Y vssd1 vssd1 vccd1 vccd1 _13856_/Z sky130_fd_sc_hd__ebufn_2
X_05748_ _05770_/CLK line[125] vssd1 vssd1 vccd1 vccd1 _05749_/A sky130_fd_sc_hd__dfxtp_1
XPHY_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08467_ _08467_/CLK _08468_/X vssd1 vssd1 vccd1 vccd1 _08465_/CLK sky130_fd_sc_hd__dlclkp_1
XPHY_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05679_ _05679_/A _05704_/Y vssd1 vssd1 vccd1 vccd1 _13799_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_23_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07418_ _13910_/X wr vssd1 vssd1 vccd1 vccd1 _07418_/X sky130_fd_sc_hd__and2_1
X_08398_ _13913_/X wr vssd1 vssd1 vccd1 vccd1 _08398_/X sky130_fd_sc_hd__and2_1
XPHY_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05013__D line[45] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10854__D line[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07349_ _13910_/X vssd1 vssd1 vccd1 vccd1 _07349_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[9\].VALID\[9\].FF OVHB\[9\].V/CLK A[16] vssd1 vssd1 vccd1 vccd1 OVHB\[9\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13230__D line[80] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10360_ _10390_/CLK line[48] vssd1 vssd1 vccd1 vccd1 _10361_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_109_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09019_ _09025_/CLK line[70] vssd1 vssd1 vccd1 vccd1 _09020_/A sky130_fd_sc_hd__dfxtp_1
X_10291_ _10291_/A _10324_/Y vssd1 vssd1 vccd1 vccd1 _13651_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_124_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12424__A _13935_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12030_ _12030_/A _12039_/Y vssd1 vssd1 vccd1 vccd1 _13710_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12143__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11685__D line[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06779__D line[70] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09155__D line[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05038__A _13931_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13981_ _13982_/A _13982_/B _13982_/C _13982_/D vssd1 vssd1 vccd1 vccd1 _13981_/X
+ sky130_fd_sc_hd__and4b_4
XANTENNA_DATA\[25\].CLKBUF\[4\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12932_ _12932_/A _12949_/Y vssd1 vssd1 vccd1 vccd1 _13772_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_37_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XOVHB\[24\].VALID\[3\].TOBUF OVHB\[24\].VALID\[3\].FF/Q OVHB\[24\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04919_/B2 sky130_fd_sc_hd__ebufn_2
X_12863_ _12875_/CLK line[35] vssd1 vssd1 vccd1 vccd1 _12864_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13405__D line[32] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[21\].VALID\[1\].FF_D A[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11814_ _11814_/A _11829_/Y vssd1 vssd1 vccd1 vccd1 _13774_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12794_ _12794_/A _12809_/Y vssd1 vssd1 vccd1 vccd1 _13634_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07403__D line[99] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11745_ _11755_/CLK line[36] vssd1 vssd1 vccd1 vccd1 _11746_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08084__A _13932_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11676_ _11676_/A _11689_/Y vssd1 vssd1 vccd1 vccd1 _13636_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12318__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13415_ _13435_/CLK line[46] vssd1 vssd1 vccd1 vccd1 _13416_/A sky130_fd_sc_hd__dfxtp_1
X_10627_ _10635_/CLK line[37] vssd1 vssd1 vccd1 vccd1 _10628_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[14\].VALID\[5\].FF_D A[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13346_ _13346_/A _13369_/Y vssd1 vssd1 vccd1 vccd1 _13626_/Z sky130_fd_sc_hd__ebufn_2
X_10558_ _10558_/A _10569_/Y vssd1 vssd1 vccd1 vccd1 _13638_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.M\[3\].MUX\[2\]_A3 _13863_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13277_ _13295_/CLK line[111] vssd1 vssd1 vccd1 vccd1 _13278_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_154_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10489_ _10495_/CLK line[102] vssd1 vssd1 vccd1 vccd1 _10490_/A sky130_fd_sc_hd__dfxtp_1
X_12228_ _12228_/A _12249_/Y vssd1 vssd1 vccd1 vccd1 _13628_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11595__D line[110] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06689__D line[43] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12159_ _12175_/CLK line[97] vssd1 vssd1 vccd1 vccd1 _12160_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05593__D line[40] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09065__D line[96] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_04981_ _04981_/A _05004_/Y vssd1 vssd1 vccd1 vccd1 _13661_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_111_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06720_ _06750_/CLK line[48] vssd1 vssd1 vccd1 vccd1 _06721_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08259__A _13932_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06651_ _06651_/A _06684_/Y vssd1 vssd1 vccd1 vccd1 _13651_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_37_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05602_ _05630_/CLK line[58] vssd1 vssd1 vccd1 vccd1 _05603_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_91_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09370_ _09370_/A _09379_/Y vssd1 vssd1 vccd1 vccd1 _13850_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__04937__D line[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06582_ _06610_/CLK line[122] vssd1 vssd1 vccd1 vccd1 _06583_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[16\].VALID\[9\].TOBUF OVHB\[16\].VALID\[9\].FF/Q OVHB\[16\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04914_/B2 sky130_fd_sc_hd__ebufn_2
X_08321_ _08325_/CLK line[7] vssd1 vssd1 vccd1 vccd1 _08322_/A sky130_fd_sc_hd__dfxtp_1
X_05533_ _05533_/A _05564_/Y vssd1 vssd1 vccd1 vccd1 _13653_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_177_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08252_ _08252_/A _08259_/Y vssd1 vssd1 vccd1 vccd1 _13852_/Z sky130_fd_sc_hd__ebufn_2
X_05464_ _05490_/CLK line[123] vssd1 vssd1 vccd1 vccd1 _05465_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[30\].VALID\[2\].TOBUF OVHB\[30\].VALID\[2\].FF/Q OVHB\[30\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04930_/B2 sky130_fd_sc_hd__ebufn_2
X_07203_ _07205_/CLK line[8] vssd1 vssd1 vccd1 vccd1 _07204_/A sky130_fd_sc_hd__dfxtp_1
X_08183_ _08185_/CLK line[72] vssd1 vssd1 vccd1 vccd1 _08184_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[20\].V_D TIE/HI vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05395_ _05395_/A _05424_/Y vssd1 vssd1 vccd1 vccd1 _13795_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13050__D line[121] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05768__D line[120] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07134_ _07134_/A _07139_/Y vssd1 vssd1 vccd1 vccd1 _13854_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08144__D line[54] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[18\].VALID\[1\].FF OVHB\[18\].V/CLK A[8] vssd1 vssd1 vccd1 vccd1 OVHB\[18\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_07065_ _07065_/CLK line[73] vssd1 vssd1 vccd1 vccd1 _07066_/A sky130_fd_sc_hd__dfxtp_1
X_06016_ _06016_/A _06019_/Y vssd1 vssd1 vccd1 vccd1 _13856_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[12\].CGAND_B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09553__A _13920_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07967_ _07975_/CLK line[101] vssd1 vssd1 vccd1 vccd1 _07968_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[16\].CGAND_A _13909_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09706_ _09706_/A _09729_/Y vssd1 vssd1 vccd1 vccd1 _13626_/Z sky130_fd_sc_hd__ebufn_2
X_06918_ _06918_/A _06929_/Y vssd1 vssd1 vccd1 vccd1 _13638_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07898_ _07898_/A _07909_/Y vssd1 vssd1 vccd1 vccd1 _13778_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09703__D line[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09637_ _09655_/CLK line[111] vssd1 vssd1 vccd1 vccd1 _09638_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_16_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06849_ _06855_/CLK line[102] vssd1 vssd1 vccd1 vccd1 _06850_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13225__D line[73] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08319__D line[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09568_ _09568_/A _09589_/Y vssd1 vssd1 vccd1 vccd1 _13768_/Z sky130_fd_sc_hd__ebufn_2
XPHY_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08519_ _08535_/CLK line[97] vssd1 vssd1 vccd1 vccd1 _08520_/A sky130_fd_sc_hd__dfxtp_1
XPHY_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09499_ _09515_/CLK line[33] vssd1 vssd1 vccd1 vccd1 _09500_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_168_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[27\].VALID\[5\].FF_D A[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11530_ _11530_/A _11549_/Y vssd1 vssd1 vccd1 vccd1 _13770_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10584__D line[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11461_ _11475_/CLK line[34] vssd1 vssd1 vccd1 vccd1 _11462_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05678__D line[93] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13200_ _13200_/A _13229_/Y vssd1 vssd1 vccd1 vccd1 _13760_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08054__D line[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10412_ _10412_/A _10429_/Y vssd1 vssd1 vccd1 vccd1 _13772_/Z sky130_fd_sc_hd__ebufn_2
X_11392_ _11392_/A _11409_/Y vssd1 vssd1 vccd1 vccd1 _13632_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09728__A _13921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XOVHB\[22\].VALID\[8\].TOBUF OVHB\[22\].VALID\[8\].FF/Q OVHB\[22\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04931_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_99_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13131_ _13155_/CLK line[44] vssd1 vssd1 vccd1 vccd1 _13132_/A sky130_fd_sc_hd__dfxtp_1
X_10343_ _10355_/CLK line[35] vssd1 vssd1 vccd1 vccd1 _10344_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07893__D line[67] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10274_ _10274_/A _10289_/Y vssd1 vssd1 vccd1 vccd1 _13634_/Z sky130_fd_sc_hd__ebufn_2
X_13062_ _13062_/A _13089_/Y vssd1 vssd1 vccd1 vccd1 _13622_/Z sky130_fd_sc_hd__ebufn_2
X_12013_ _12035_/CLK line[45] vssd1 vssd1 vccd1 vccd1 _12014_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_105_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XOVHB\[6\].VALID\[12\].TOBUF OVHB\[6\].VALID\[12\].FF/Q OVHB\[6\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04929_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__06302__D line[122] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[16\].VALID\[3\].FF OVHB\[16\].V/CLK A[10] vssd1 vssd1 vccd1 vccd1 OVHB\[16\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_93_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13964_ _13971_/A _13971_/B _13971_/C _13971_/D vssd1 vssd1 vccd1 vccd1 _13964_/Y
+ sky130_fd_sc_hd__nor4b_4
XFILLER_74_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10759__D line[97] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12915_ _12945_/CLK line[64] vssd1 vssd1 vccd1 vccd1 _12916_/A sky130_fd_sc_hd__dfxtp_1
X_13895_ A[2] vssd1 vssd1 vccd1 vccd1 _13905_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__13135__D line[46] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12846_ _12846_/A _12879_/Y vssd1 vssd1 vccd1 vccd1 _13686_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08229__D line[107] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07133__D line[104] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[23\].CLKBUF\[6\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12974__D line[86] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12777_ _12805_/CLK line[10] vssd1 vssd1 vccd1 vccd1 _12778_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11233__A _13933_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11728_ _11728_/A _11759_/Y vssd1 vssd1 vccd1 vccd1 _13688_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11659_ _11685_/CLK line[11] vssd1 vssd1 vccd1 vccd1 _11660_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05180_ _05210_/CLK line[112] vssd1 vssd1 vccd1 vccd1 _05181_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_116_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13329_ _13329_/A _13334_/Y vssd1 vssd1 vccd1 vccd1 _13889_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[16\].VALID\[13\].FF_D A[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MUX.M\[2\].MUX\[3\]_A1 _13739_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[8\].VALID\[0\].FF_D A[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08870_ _08870_/A _08889_/Y vssd1 vssd1 vccd1 vccd1 _13630_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07308__D line[56] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07821_ _07835_/CLK line[34] vssd1 vssd1 vccd1 vccd1 _07822_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_96_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11408__A _13926_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_04964_ _04964_/A _04969_/Y vssd1 vssd1 vccd1 vccd1 _13644_/Z sky130_fd_sc_hd__ebufn_2
X_07752_ _07752_/A _07769_/Y vssd1 vssd1 vccd1 vccd1 _13632_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[5\].V_D TIE/HI vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06703_ _06715_/CLK line[35] vssd1 vssd1 vccd1 vccd1 _06704_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[6\].VALID\[0\].TOBUF OVHB\[6\].VALID\[0\].FF/Q OVHB\[6\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04924_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[26\].VALID\[12\].FF_D A[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07683_ _07695_/CLK line[99] vssd1 vssd1 vccd1 vccd1 _07684_/A sky130_fd_sc_hd__dfxtp_1
X_09422_ _09422_/A _09449_/Y vssd1 vssd1 vccd1 vccd1 _13622_/Z sky130_fd_sc_hd__ebufn_2
X_06634_ _06634_/A _06649_/Y vssd1 vssd1 vccd1 vccd1 _13634_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[14\].VALID\[5\].FF OVHB\[14\].V/CLK A[12] vssd1 vssd1 vccd1 vccd1 OVHB\[14\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07043__D line[77] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09353_ _09375_/CLK line[109] vssd1 vssd1 vccd1 vccd1 _09354_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12884__D line[59] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06565_ _06575_/CLK line[100] vssd1 vssd1 vccd1 vccd1 _06566_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[31\].VALID\[9\].FF OVHB\[31\].V/CLK A[16] vssd1 vssd1 vccd1 vccd1 OVHB\[31\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_08304_ _08304_/A _08329_/Y vssd1 vssd1 vccd1 vccd1 _13624_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06882__D line[117] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05516_ _05516_/A _05529_/Y vssd1 vssd1 vccd1 vccd1 _13636_/Z sky130_fd_sc_hd__ebufn_2
X_06496_ _06496_/A _06509_/Y vssd1 vssd1 vccd1 vccd1 _13776_/Z sky130_fd_sc_hd__ebufn_2
X_09284_ _09284_/A _09309_/Y vssd1 vssd1 vccd1 vccd1 _13764_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_166_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05447_ _05455_/CLK line[101] vssd1 vssd1 vccd1 vccd1 _05448_/A sky130_fd_sc_hd__dfxtp_1
X_08235_ _08255_/CLK line[110] vssd1 vssd1 vccd1 vccd1 _08236_/A sky130_fd_sc_hd__dfxtp_1
X_05378_ _05378_/A _05389_/Y vssd1 vssd1 vccd1 vccd1 _13778_/Z sky130_fd_sc_hd__ebufn_2
X_08166_ _08166_/A _08189_/Y vssd1 vssd1 vccd1 vccd1 _13766_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_118_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07117_ _07135_/CLK line[111] vssd1 vssd1 vccd1 vccd1 _07118_/A sky130_fd_sc_hd__dfxtp_1
X_08097_ _08115_/CLK line[47] vssd1 vssd1 vccd1 vccd1 _08098_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_161_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07048_ _07048_/A _07069_/Y vssd1 vssd1 vccd1 vccd1 _13768_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07068__A _13909_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12124__D line[81] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07218__D line[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11963__D line[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08999_ _09025_/CLK line[75] vssd1 vssd1 vccd1 vccd1 _09000_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_87_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[29\].VALID\[14\].TOBUF OVHB\[29\].VALID\[14\].FF/Q OVHB\[29\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_47_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09433__D line[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10961_ _10985_/CLK line[76] vssd1 vssd1 vccd1 vccd1 _10962_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_90_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12700_ _12700_/CLK line[89] vssd1 vssd1 vccd1 vccd1 _12701_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_55_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13680_ _13680_/CLK line[25] vssd1 vssd1 vccd1 vccd1 _13681_/A sky130_fd_sc_hd__dfxtp_1
X_10892_ _10892_/A _10919_/Y vssd1 vssd1 vccd1 vccd1 _13692_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_203_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12631_ _12631_/A _12634_/Y vssd1 vssd1 vccd1 vccd1 _13751_/Z sky130_fd_sc_hd__ebufn_2
XPHY_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[10\].VALID\[8\].FF_D A[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06792__D line[90] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12562_ _12562_/CLK _12563_/X vssd1 vssd1 vccd1 vccd1 _12560_/CLK sky130_fd_sc_hd__dlclkp_1
XPHY_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11513_ _13926_/X wr vssd1 vssd1 vccd1 vccd1 _11513_/X sky130_fd_sc_hd__and2_1
XPHY_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12493_ _13935_/X wr vssd1 vssd1 vccd1 vccd1 _12493_/X sky130_fd_sc_hd__and2_1
XOVHB\[24\].INV _13964_/Y vssd1 vssd1 vccd1 vccd1 OVHB\[24\].INV/Y sky130_fd_sc_hd__inv_2
XFILLER_184_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[12\].VALID\[7\].FF OVHB\[12\].V/CLK A[14] vssd1 vssd1 vccd1 vccd1 OVHB\[12\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11444_ _13926_/X vssd1 vssd1 vccd1 vccd1 _11444_/Y sky130_fd_sc_hd__inv_2
XFILLER_144_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11375_ _11405_/CLK line[0] vssd1 vssd1 vccd1 vccd1 _11376_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09608__D line[83] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13114_ _13120_/CLK line[22] vssd1 vssd1 vccd1 vccd1 _13115_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[22\].VALID\[13\].TOBUF OVHB\[22\].VALID\[13\].FF/Q OVHB\[22\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04916_/B2 sky130_fd_sc_hd__ebufn_2
X_10326_ _10326_/A _10359_/Y vssd1 vssd1 vccd1 vccd1 _13686_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_140_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13045_ _13045_/A _13054_/Y vssd1 vssd1 vccd1 vccd1 _13885_/Z sky130_fd_sc_hd__ebufn_2
X_10257_ _10285_/CLK line[10] vssd1 vssd1 vccd1 vccd1 _10258_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[24\].V OVHB\[24\].V/CLK TIE/HI rst_n vssd1 vssd1 vccd1 vccd1 OVHB\[24\].V/Q
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_59_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06032__D line[127] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10188_ _10188_/A _10219_/Y vssd1 vssd1 vccd1 vccd1 _13828_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11873__D line[109] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06967__D line[42] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__04926__B2 _04926_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05871__D line[39] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10489__D line[102] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13947_ _13949_/B _13949_/A _13949_/C _13949_/D vssd1 vssd1 vccd1 vccd1 _13947_/X
+ sky130_fd_sc_hd__and4b_4
XFILLER_46_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13878_ _13890_/CLK line[115] vssd1 vssd1 vccd1 vccd1 _13879_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_62_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12829_ _12829_/A _12844_/Y vssd1 vssd1 vccd1 vccd1 _13669_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_188_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07798__D line[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06350_ _06350_/A _06369_/Y vssd1 vssd1 vccd1 vccd1 _13630_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_203_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05301_ _05315_/CLK line[34] vssd1 vssd1 vccd1 vccd1 _05302_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11898__A _13927_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06281_ _06295_/CLK line[98] vssd1 vssd1 vccd1 vccd1 _06282_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11113__D line[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDATA\[29\].CLKBUF\[3\] clk vssd1 vssd1 vccd1 vccd1 _10952_/CLK sky130_fd_sc_hd__clkbuf_4
X_08020_ _08020_/A _08049_/Y vssd1 vssd1 vccd1 vccd1 _13620_/Z sky130_fd_sc_hd__ebufn_2
X_05232_ _05232_/A _05249_/Y vssd1 vssd1 vccd1 vccd1 _13632_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06207__D line[79] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05163_ _05175_/CLK line[99] vssd1 vssd1 vccd1 vccd1 _05164_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[4\].VALID\[5\].TOBUF OVHB\[4\].VALID\[5\].FF/Q OVHB\[4\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04927_/B2 sky130_fd_sc_hd__ebufn_2
XOVHB\[10\].VOBUF OVHB\[10\].V/Q OVHB\[10\].INV/Y vssd1 vssd1 vccd1 vccd1 _04912_/B1
+ sky130_fd_sc_hd__ebufn_2
XANTENNA__08422__D line[53] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09971_ _09971_/A _09974_/Y vssd1 vssd1 vccd1 vccd1 _13891_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_89_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05094_ _05094_/A _05109_/Y vssd1 vssd1 vccd1 vccd1 _13774_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_131_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XOVHB\[29\].VALID\[8\].TOBUF OVHB\[29\].VALID\[8\].FF/Q OVHB\[29\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04931_/B2 sky130_fd_sc_hd__ebufn_2
X_08922_ _08922_/CLK _08923_/X vssd1 vssd1 vccd1 vccd1 _08920_/CLK sky130_fd_sc_hd__dlclkp_1
XOVHB\[10\].VALID\[9\].FF OVHB\[10\].V/CLK A[16] vssd1 vssd1 vccd1 vccd1 OVHB\[10\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_112_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XOVHB\[15\].V OVHB\[15\].V/CLK TIE/HI rst_n vssd1 vssd1 vccd1 vccd1 OVHB\[15\].V/Q
+ sky130_fd_sc_hd__dfrtp_1
X_08853_ _13914_/X wr vssd1 vssd1 vccd1 vccd1 _08853_/X sky130_fd_sc_hd__and2_1
XFILLER_29_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_OVHB\[30\].VALID\[4\].FF_D A[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07804_ _13912_/X vssd1 vssd1 vccd1 vccd1 _07804_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08784_ _13914_/X vssd1 vssd1 vccd1 vccd1 _08784_/Y sky130_fd_sc_hd__inv_2
XANTENNA__05781__D line[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05996_ _05996_/A _06019_/Y vssd1 vssd1 vccd1 vccd1 _13836_/Z sky130_fd_sc_hd__ebufn_2
X_07735_ _07765_/CLK line[0] vssd1 vssd1 vccd1 vccd1 _07736_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10399__D line[75] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_04947_ _04965_/CLK line[15] vssd1 vssd1 vccd1 vccd1 _04948_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_37_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07666_ _07666_/A _07699_/Y vssd1 vssd1 vccd1 vccd1 _13826_/Z sky130_fd_sc_hd__ebufn_2
X_09405_ _09405_/A _09414_/Y vssd1 vssd1 vccd1 vccd1 _13885_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[23\].VALID\[8\].FF_D A[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06617_ _06645_/CLK line[10] vssd1 vssd1 vccd1 vccd1 _06618_/A sky130_fd_sc_hd__dfxtp_1
X_07597_ _07625_/CLK line[74] vssd1 vssd1 vccd1 vccd1 _07598_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13503__D line[72] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09336_ _09340_/CLK line[87] vssd1 vssd1 vccd1 vccd1 _09337_/A sky130_fd_sc_hd__dfxtp_1
X_06548_ _06548_/A _06579_/Y vssd1 vssd1 vccd1 vccd1 _13828_/Z sky130_fd_sc_hd__ebufn_2
X_09267_ _09267_/A _09274_/Y vssd1 vssd1 vccd1 vccd1 _13747_/Z sky130_fd_sc_hd__ebufn_2
X_06479_ _06505_/CLK line[75] vssd1 vssd1 vccd1 vccd1 _06480_/A sky130_fd_sc_hd__dfxtp_1
X_08218_ _08220_/CLK line[88] vssd1 vssd1 vccd1 vccd1 _08219_/A sky130_fd_sc_hd__dfxtp_1
X_09198_ _09200_/CLK line[24] vssd1 vssd1 vccd1 vccd1 _09199_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05021__D line[34] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10862__D line[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08149_ _08149_/A _08154_/Y vssd1 vssd1 vccd1 vccd1 _13749_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05956__D line[92] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08332__D line[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDATA\[28\].CLKBUF\[0\] clk vssd1 vssd1 vccd1 vccd1 _10567_/CLK sky130_fd_sc_hd__clkbuf_4
X_11160_ _11160_/CLK line[25] vssd1 vssd1 vccd1 vccd1 _11161_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_136_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10111_ _10111_/A _10114_/Y vssd1 vssd1 vccd1 vccd1 _13751_/Z sky130_fd_sc_hd__ebufn_2
X_11091_ _11091_/A _11094_/Y vssd1 vssd1 vccd1 vccd1 _13891_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[18\].CLKBUF\[6\] clk vssd1 vssd1 vccd1 vccd1 _07697_/CLK sky130_fd_sc_hd__clkbuf_4
X_10042_ _10042_/CLK _10043_/X vssd1 vssd1 vccd1 vccd1 _10040_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__12789__D line[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09163__D line[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XOVHB\[11\].VALID\[0\].TOBUF OVHB\[11\].VALID\[0\].FF/Q OVHB\[11\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04924_/B2 sky130_fd_sc_hd__ebufn_2
X_13801_ _13801_/A _13824_/Y vssd1 vssd1 vccd1 vccd1 _13801_/Z sky130_fd_sc_hd__ebufn_2
X_11993_ _11993_/A _12004_/Y vssd1 vssd1 vccd1 vccd1 _13673_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13263__A _13938_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13732_ _13750_/CLK line[63] vssd1 vssd1 vccd1 vccd1 _13733_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10102__D line[53] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10944_ _10950_/CLK line[54] vssd1 vssd1 vccd1 vccd1 _10945_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_204_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13663_ _13663_/A _13684_/Y vssd1 vssd1 vccd1 vccd1 _13663_/Z sky130_fd_sc_hd__ebufn_2
X_10875_ _10875_/A _10884_/Y vssd1 vssd1 vccd1 vccd1 _13675_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13413__D line[45] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12614_ _12630_/CLK line[49] vssd1 vssd1 vccd1 vccd1 _12615_/A sky130_fd_sc_hd__dfxtp_1
XPHY_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08507__D line[106] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13594_ _13610_/CLK line[113] vssd1 vssd1 vccd1 vccd1 _13595_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07411__D line[103] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12545_ _12545_/A _12564_/Y vssd1 vssd1 vccd1 vccd1 _13665_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12029__D line[38] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12476_ _12490_/CLK line[114] vssd1 vssd1 vccd1 vccd1 _12477_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[5\].VALID\[0\].FF OVHB\[5\].V/CLK A[7] vssd1 vssd1 vccd1 vccd1 OVHB\[5\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_11427_ _11427_/A _11444_/Y vssd1 vssd1 vccd1 vccd1 _13667_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[18\].CG_CLK clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[16\].CLKBUF\[0\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[4\].VALID\[3\].FF_D A[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09338__D line[88] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11358_ _11370_/CLK line[115] vssd1 vssd1 vccd1 vccd1 _11359_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_98_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10309_ _10309_/A _10324_/Y vssd1 vssd1 vccd1 vccd1 _13669_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_112_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13438__A _13898_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11289_ _11289_/A _11304_/Y vssd1 vssd1 vccd1 vccd1 _13809_/Z sky130_fd_sc_hd__ebufn_2
X_13028_ _13050_/CLK line[125] vssd1 vssd1 vccd1 vccd1 _13029_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_67_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06697__D line[47] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05850_ _05850_/A _05879_/Y vssd1 vssd1 vccd1 vccd1 _13690_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09073__D line[109] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDATA\[17\].CLKBUF\[3\] clk vssd1 vssd1 vccd1 vccd1 _07312_/CLK sky130_fd_sc_hd__clkbuf_4
X_05781_ _05805_/CLK line[12] vssd1 vssd1 vccd1 vccd1 _05782_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_19_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10012__D line[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07520_ _07520_/CLK line[25] vssd1 vssd1 vccd1 vccd1 _07521_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[9\].CLKBUF\[0\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07451_ _07451_/A _07454_/Y vssd1 vssd1 vccd1 vccd1 _13891_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_210_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06402_ _06402_/CLK _06403_/X vssd1 vssd1 vccd1 vccd1 _06400_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__04945__D line[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07382_ _07382_/CLK _07383_/X vssd1 vssd1 vccd1 vccd1 _07380_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__07321__D line[76] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09121_ _09121_/A _09134_/Y vssd1 vssd1 vccd1 vccd1 _13881_/Z sky130_fd_sc_hd__ebufn_2
X_06333_ _13903_/X wr vssd1 vssd1 vccd1 vccd1 _06333_/X sky130_fd_sc_hd__and2_1
XFILLER_175_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09052_ _09060_/CLK line[85] vssd1 vssd1 vccd1 vccd1 _09053_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09098__A _13915_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06264_ _13903_/X vssd1 vssd1 vccd1 vccd1 _06264_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11778__D line[51] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05215_ _05245_/CLK line[0] vssd1 vssd1 vccd1 vccd1 _05216_/A sky130_fd_sc_hd__dfxtp_1
X_08003_ _08003_/A _08014_/Y vssd1 vssd1 vccd1 vccd1 _13883_/Z sky130_fd_sc_hd__ebufn_2
X_06195_ _06225_/CLK line[64] vssd1 vssd1 vccd1 vccd1 _06196_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_128_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09248__D line[61] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05146_ _05146_/A _05179_/Y vssd1 vssd1 vccd1 vccd1 _13826_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[17\].CGAND _13910_/X wr vssd1 vssd1 vccd1 vccd1 OVHB\[17\].CGAND/X sky130_fd_sc_hd__and2_4
X_09954_ _09970_/CLK line[113] vssd1 vssd1 vccd1 vccd1 _09955_/A sky130_fd_sc_hd__dfxtp_1
X_05077_ _05105_/CLK line[74] vssd1 vssd1 vccd1 vccd1 _05078_/A sky130_fd_sc_hd__dfxtp_1
X_08905_ _08905_/A _08924_/Y vssd1 vssd1 vccd1 vccd1 _13665_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[3\].VALID\[2\].FF OVHB\[3\].V/CLK A[9] vssd1 vssd1 vccd1 vccd1 OVHB\[3\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_09885_ _09885_/A _09904_/Y vssd1 vssd1 vccd1 vccd1 _13805_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_112_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12402__D line[95] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08836_ _08850_/CLK line[114] vssd1 vssd1 vccd1 vccd1 _08837_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[19\].VALID\[0\].FF_D A[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06400__D line[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08767_ _08767_/A _08784_/Y vssd1 vssd1 vccd1 vccd1 _13807_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_72_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05979_ _05979_/A _05984_/Y vssd1 vssd1 vccd1 vccd1 _13819_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11018__D line[88] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07718_ _07730_/CLK line[115] vssd1 vssd1 vccd1 vccd1 _07719_/A sky130_fd_sc_hd__dfxtp_1
X_08698_ _08710_/CLK line[51] vssd1 vssd1 vccd1 vccd1 _08699_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09711__D line[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07649_ _07649_/A _07664_/Y vssd1 vssd1 vccd1 vccd1 _13809_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[16\].CLKBUF\[0\] clk vssd1 vssd1 vccd1 vccd1 _06927_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_186_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10660_ _10670_/CLK line[52] vssd1 vssd1 vccd1 vccd1 _10661_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_41_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[9\].INV _13943_/X vssd1 vssd1 vccd1 vccd1 OVHB\[9\].INV/Y sky130_fd_sc_hd__inv_2
XMUX.M\[2\].MUX\[0\] _13651_/Z _13721_/Z _13791_/Z _13861_/Z MUX.SEL0BUF\[2\]/X MUX.SEL1BUF\[2\]/X
+ vssd1 vssd1 vccd1 vccd1 Do[16] sky130_fd_sc_hd__mux4_1
XFILLER_139_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09319_ _09319_/A _09344_/Y vssd1 vssd1 vccd1 vccd1 _13799_/Z sky130_fd_sc_hd__ebufn_2
X_10591_ _10591_/A _10604_/Y vssd1 vssd1 vccd1 vccd1 _13671_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_21_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12330_ _12350_/CLK line[62] vssd1 vssd1 vccd1 vccd1 _12331_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_193_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10592__D line[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12261_ _12261_/A _12284_/Y vssd1 vssd1 vccd1 vccd1 _13661_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05686__D line[82] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08062__D line[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11212_ _11230_/CLK line[63] vssd1 vssd1 vccd1 vccd1 _11213_/A sky130_fd_sc_hd__dfxtp_1
X_12192_ _12210_/CLK line[127] vssd1 vssd1 vccd1 vccd1 _12193_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_162_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11143_ _11143_/A _11164_/Y vssd1 vssd1 vccd1 vccd1 _13663_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08997__D line[74] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05983__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11074_ _11090_/CLK line[113] vssd1 vssd1 vccd1 vccd1 _11075_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_1_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[19\].VALID\[12\].TOBUF OVHB\[19\].VALID\[12\].FF/Q OVHB\[19\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04929_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_163_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10025_ _10025_/A _10044_/Y vssd1 vssd1 vccd1 vccd1 _13665_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_76_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06310__D line[126] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11976_ _12000_/CLK line[28] vssd1 vssd1 vccd1 vccd1 _11977_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[1\].VALID\[4\].FF OVHB\[1\].V/CLK A[11] vssd1 vssd1 vccd1 vccd1 OVHB\[1\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_13715_ _13715_/CLK line[41] vssd1 vssd1 vccd1 vccd1 _13716_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_72_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10767__D line[101] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10927_ _10927_/A _10954_/Y vssd1 vssd1 vccd1 vccd1 _13727_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13143__D line[35] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13646_ _13646_/A _13649_/Y vssd1 vssd1 vccd1 vccd1 _13646_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08237__D line[111] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10858_ _10880_/CLK line[29] vssd1 vssd1 vccd1 vccd1 _10859_/A sky130_fd_sc_hd__dfxtp_1
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13577_ _13577_/CLK _13578_/X vssd1 vssd1 vccd1 vccd1 _13575_/CLK sky130_fd_sc_hd__dlclkp_1
X_10789_ _10789_/A _10814_/Y vssd1 vssd1 vccd1 vccd1 _13869_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_12_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12528_ _13936_/X wr vssd1 vssd1 vccd1 vccd1 _12528_/X sky130_fd_sc_hd__and2_1
XFILLER_157_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_MUX.M\[3\].MUX\[5\]_A1 _13729_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12459_ _13935_/X vssd1 vssd1 vccd1 vccd1 _12459_/Y sky130_fd_sc_hd__inv_2
XOVHB\[12\].VALID\[11\].TOBUF OVHB\[12\].VALID\[11\].FF/Q OVHB\[12\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04915_/B2 sky130_fd_sc_hd__ebufn_2
X_05000_ _05000_/CLK line[25] vssd1 vssd1 vccd1 vccd1 _05001_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_125_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08700__D line[52] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06951_ _06951_/A _06964_/Y vssd1 vssd1 vccd1 vccd1 _13671_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_100_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMUX.M\[1\].MUX\[2\] _13618_/Z _13688_/Z _13758_/Z _13828_/Z MUX.SEL0BUF\[1\]/X MUX.SEL1BUF\[1\]/X
+ vssd1 vssd1 vccd1 vccd1 Do[10] sky130_fd_sc_hd__mux4_1
XANTENNA_DATA\[14\].CLKBUF\[2\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13318__D line[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05902_ _05910_/CLK line[53] vssd1 vssd1 vccd1 vccd1 _05903_/A sky130_fd_sc_hd__dfxtp_1
X_09670_ _09690_/CLK line[126] vssd1 vssd1 vccd1 vccd1 _09671_/A sky130_fd_sc_hd__dfxtp_1
X_06882_ _06890_/CLK line[117] vssd1 vssd1 vccd1 vccd1 _06883_/A sky130_fd_sc_hd__dfxtp_1
X_08621_ _08621_/A _08644_/Y vssd1 vssd1 vccd1 vccd1 _13661_/Z sky130_fd_sc_hd__ebufn_2
X_05833_ _05833_/A _05844_/Y vssd1 vssd1 vccd1 vccd1 _13673_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_54_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MUX.M\[1\].MUX\[1\]_A2 _13786_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08552_ _08570_/CLK line[127] vssd1 vssd1 vccd1 vccd1 _08553_/A sky130_fd_sc_hd__dfxtp_1
X_05764_ _05770_/CLK line[118] vssd1 vssd1 vccd1 vccd1 _05765_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[18\].VALID\[0\].TOBUF OVHB\[18\].VALID\[0\].FF/Q OVHB\[18\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04924_/B2 sky130_fd_sc_hd__ebufn_2
X_07503_ _07503_/A _07524_/Y vssd1 vssd1 vccd1 vccd1 _13663_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10677__D line[74] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08483_ _08483_/A _08504_/Y vssd1 vssd1 vccd1 vccd1 _13803_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05695_ _05695_/A _05704_/Y vssd1 vssd1 vccd1 vccd1 _13815_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_22_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07434_ _07450_/CLK line[113] vssd1 vssd1 vccd1 vccd1 _07435_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07051__D line[66] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12892__D line[63] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07365_ _07365_/A _07384_/Y vssd1 vssd1 vccd1 vccd1 _13805_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07986__D line[124] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09104_ _09130_/CLK line[123] vssd1 vssd1 vccd1 vccd1 _09105_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06890__D line[121] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06316_ _06330_/CLK line[114] vssd1 vssd1 vccd1 vccd1 _06317_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[7\].CLKBUF\[2\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07296_ _07310_/CLK line[50] vssd1 vssd1 vccd1 vccd1 _07297_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_175_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09035_ _09035_/A _09064_/Y vssd1 vssd1 vccd1 vccd1 _13795_/Z sky130_fd_sc_hd__ebufn_2
X_06247_ _06247_/A _06264_/Y vssd1 vssd1 vccd1 vccd1 _13807_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_117_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06178_ _06190_/CLK line[51] vssd1 vssd1 vccd1 vccd1 _06179_/A sky130_fd_sc_hd__dfxtp_1
X_05129_ _05129_/A _05144_/Y vssd1 vssd1 vccd1 vccd1 _13809_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_77_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08610__D line[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09937_ _09937_/CLK _09938_/X vssd1 vssd1 vccd1 vccd1 _09935_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_131_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12132__D line[85] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09868_ _13921_/X wr vssd1 vssd1 vccd1 vccd1 _09868_/X sky130_fd_sc_hd__and2_1
XANTENNA__07226__D line[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07804__A _13912_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08819_ _13914_/X vssd1 vssd1 vccd1 vccd1 _08819_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09799_ _13921_/X vssd1 vssd1 vccd1 vccd1 _09799_/Y sky130_fd_sc_hd__inv_2
X_11830_ _11860_/CLK line[80] vssd1 vssd1 vccd1 vccd1 _11831_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07523__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09441__D line[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11761_ _11761_/A _11794_/Y vssd1 vssd1 vccd1 vccd1 _13721_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13500_ _13500_/A _13509_/Y vssd1 vssd1 vccd1 vccd1 _13780_/Z sky130_fd_sc_hd__ebufn_2
X_10712_ _10740_/CLK line[90] vssd1 vssd1 vccd1 vccd1 _10713_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11692_ _11720_/CLK line[26] vssd1 vssd1 vccd1 vccd1 _11693_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMUX.M\[0\].MUX\[4\] _13636_/Z _13706_/Z _13776_/Z _13846_/Z MUX.SEL0BUF\[0\]/X MUX.SEL1BUF\[0\]/X
+ vssd1 vssd1 vccd1 vccd1 Do[4] sky130_fd_sc_hd__mux4_1
XPHY_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13431_ _13435_/CLK line[39] vssd1 vssd1 vccd1 vccd1 _13432_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_9_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10643_ _10643_/A _10674_/Y vssd1 vssd1 vccd1 vccd1 _13723_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13362_ _13362_/A _13369_/Y vssd1 vssd1 vccd1 vccd1 _13642_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[0\].VALID\[6\].FF_D A[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10574_ _10600_/CLK line[27] vssd1 vssd1 vccd1 vccd1 _10575_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_194_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12313_ _12315_/CLK line[40] vssd1 vssd1 vccd1 vccd1 _12314_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12307__D line[37] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13293_ _13295_/CLK line[104] vssd1 vssd1 vccd1 vccd1 _13294_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_108_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12244_ _12244_/A _12249_/Y vssd1 vssd1 vccd1 vccd1 _13644_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_154_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12175_ _12175_/CLK line[105] vssd1 vssd1 vccd1 vccd1 _12176_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_69_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09616__D line[87] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11126_ _11126_/A _11129_/Y vssd1 vssd1 vccd1 vccd1 _13646_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_150_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12042__D line[58] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11057_ _11057_/CLK _11058_/X vssd1 vssd1 vccd1 vccd1 _11055_/CLK sky130_fd_sc_hd__dlclkp_1
X_10008_ _13922_/X wr vssd1 vssd1 vccd1 vccd1 _10008_/X sky130_fd_sc_hd__and2_1
XANTENNA__06040__D line[116] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[24\].VALID\[14\].FF OVHB\[24\].V/CLK A[21] vssd1 vssd1 vccd1 vccd1 OVHB\[24\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11881__D line[98] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06975__D line[46] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09351__D line[108] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11959_ _11965_/CLK line[6] vssd1 vssd1 vccd1 vccd1 _11960_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_17_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_OVHB\[3\].VALID\[12\].FF_D A[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05480_ _05490_/CLK line[116] vssd1 vssd1 vccd1 vccd1 _05481_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[26\].VALID\[1\].FF OVHB\[26\].V/CLK A[8] vssd1 vssd1 vccd1 vccd1 OVHB\[26\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_13629_ _13645_/CLK line[1] vssd1 vssd1 vccd1 vccd1 _13630_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07150_ _07170_/CLK line[126] vssd1 vssd1 vccd1 vccd1 _07151_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_157_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06101_ _06101_/A _06124_/Y vssd1 vssd1 vccd1 vccd1 _13661_/Z sky130_fd_sc_hd__ebufn_2
X_07081_ _07081_/A _07104_/Y vssd1 vssd1 vccd1 vccd1 _13801_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12217__D line[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11121__D line[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06215__D line[68] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06032_ _06050_/CLK line[127] vssd1 vssd1 vccd1 vccd1 _06033_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_160_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XOVHB\[16\].VALID\[5\].TOBUF OVHB\[16\].VALID\[5\].FF/Q OVHB\[16\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04927_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__09526__D line[60] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08430__D line[57] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07983_ _07983_/A _08014_/Y vssd1 vssd1 vccd1 vccd1 _13863_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[15\].VALID\[3\].FF_D A[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13048__D line[120] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09722_ _09722_/A _09729_/Y vssd1 vssd1 vccd1 vccd1 _13642_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_68_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XDATA\[8\].CLKBUF\[7\] clk vssd1 vssd1 vccd1 vccd1 _13612_/CLK sky130_fd_sc_hd__clkbuf_4
X_06934_ _06960_/CLK line[27] vssd1 vssd1 vccd1 vccd1 _06935_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_86_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09653_ _09655_/CLK line[104] vssd1 vssd1 vccd1 vccd1 _09654_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_67_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06865_ _06865_/A _06894_/Y vssd1 vssd1 vccd1 vccd1 _13865_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_28_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08604_ _08604_/A _08609_/Y vssd1 vssd1 vccd1 vccd1 _13644_/Z sky130_fd_sc_hd__ebufn_2
X_05816_ _05840_/CLK line[28] vssd1 vssd1 vccd1 vccd1 _05817_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_103_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09584_ _09584_/A _09589_/Y vssd1 vssd1 vccd1 vccd1 _13784_/Z sky130_fd_sc_hd__ebufn_2
X_06796_ _06820_/CLK line[92] vssd1 vssd1 vccd1 vccd1 _06797_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05144__A _13931_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08535_ _08535_/CLK line[105] vssd1 vssd1 vccd1 vccd1 _08536_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[12\].CLKBUF\[4\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05747_ _05747_/A _05774_/Y vssd1 vssd1 vccd1 vccd1 _13867_/Z sky130_fd_sc_hd__ebufn_2
XPHY_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MUX.M\[0\].MUX\[2\]_A0 _13632_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08466_ _08466_/A _08469_/Y vssd1 vssd1 vccd1 vccd1 _13786_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05678_ _05700_/CLK line[93] vssd1 vssd1 vccd1 vccd1 _05679_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_50_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07417_ _07417_/CLK _07418_/X vssd1 vssd1 vccd1 vccd1 _07415_/CLK sky130_fd_sc_hd__dlclkp_1
XPHY_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08397_ _08397_/CLK _08398_/X vssd1 vssd1 vccd1 vccd1 _08395_/CLK sky130_fd_sc_hd__dlclkp_1
XPHY_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08605__D line[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07348_ _13910_/X wr vssd1 vssd1 vccd1 vccd1 _07348_/X sky130_fd_sc_hd__and2_1
XFILLER_12_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07279_ _13910_/X vssd1 vssd1 vccd1 vccd1 _07279_/Y sky130_fd_sc_hd__inv_2
XFILLER_164_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11031__D line[108] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XOVHB\[24\].VALID\[3\].FF OVHB\[24\].V/CLK A[10] vssd1 vssd1 vccd1 vccd1 OVHB\[24\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09018_ _09018_/A _09029_/Y vssd1 vssd1 vccd1 vccd1 _13778_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06125__D line[32] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10290_ _10320_/CLK line[16] vssd1 vssd1 vccd1 vccd1 _10291_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_117_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10870__D line[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[5\].CLKBUF\[4\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05964__D line[81] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08340__D line[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05319__A _13900_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05038__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13980_ _13982_/B _13982_/A _13982_/C _13982_/D vssd1 vssd1 vccd1 vccd1 _13980_/X
+ sky130_fd_sc_hd__and4b_4
XANTENNA_DATA\[31\].CLKBUF\[6\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12931_ _12945_/CLK line[66] vssd1 vssd1 vccd1 vccd1 _12932_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12797__D line[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12862_ _12862_/A _12879_/Y vssd1 vssd1 vccd1 vccd1 _13702_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[22\].VALID\[4\].TOBUF OVHB\[22\].VALID\[4\].FF/Q OVHB\[22\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04925_/B2 sky130_fd_sc_hd__ebufn_2
XDATA\[7\].CLKBUF\[4\] clk vssd1 vssd1 vccd1 vccd1 _13227_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_73_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11813_ _11825_/CLK line[67] vssd1 vssd1 vccd1 vccd1 _11814_/A sky130_fd_sc_hd__dfxtp_1
X_12793_ _12805_/CLK line[3] vssd1 vssd1 vccd1 vccd1 _12794_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_27_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11206__D line[60] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10110__D line[57] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11744_ _11744_/A _11759_/Y vssd1 vssd1 vccd1 vccd1 _13704_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_186_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05204__D line[118] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11675_ _11685_/CLK line[4] vssd1 vssd1 vccd1 vccd1 _11676_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13421__D line[34] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13414_ _13414_/A _13439_/Y vssd1 vssd1 vccd1 vccd1 _13694_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10626_ _10626_/A _10639_/Y vssd1 vssd1 vccd1 vccd1 _13706_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08515__D line[110] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13345_ _13365_/CLK line[14] vssd1 vssd1 vccd1 vccd1 _13346_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_10_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10557_ _10565_/CLK line[5] vssd1 vssd1 vccd1 vccd1 _10558_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_127_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13276_ _13276_/A _13299_/Y vssd1 vssd1 vccd1 vccd1 _13836_/Z sky130_fd_sc_hd__ebufn_2
X_10488_ _10488_/A _10499_/Y vssd1 vssd1 vccd1 vccd1 _13848_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06613__A _13904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10780__D line[112] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12227_ _12245_/CLK line[15] vssd1 vssd1 vccd1 vccd1 _12228_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_170_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_OVHB\[28\].VALID\[3\].FF_D A[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12158_ _12158_/A _12179_/Y vssd1 vssd1 vccd1 vccd1 _13838_/Z sky130_fd_sc_hd__ebufn_2
X_11109_ _11125_/CLK line[1] vssd1 vssd1 vccd1 vccd1 _11110_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_111_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_04980_ _05000_/CLK line[30] vssd1 vssd1 vccd1 vccd1 _04981_/A sky130_fd_sc_hd__dfxtp_1
X_12089_ _12105_/CLK line[65] vssd1 vssd1 vccd1 vccd1 _12090_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[22\].VALID\[5\].FF OVHB\[22\].V/CLK A[12] vssd1 vssd1 vccd1 vccd1 OVHB\[22\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_209_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[30\].VALID\[10\].FF OVHB\[30\].V/CLK A[17] vssd1 vssd1 vccd1 vccd1 OVHB\[30\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_06650_ _06680_/CLK line[16] vssd1 vssd1 vccd1 vccd1 _06651_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_25_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09081__D line[98] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05601_ _05601_/A _05634_/Y vssd1 vssd1 vccd1 vccd1 _13721_/Z sky130_fd_sc_hd__ebufn_2
X_06581_ _06581_/A _06614_/Y vssd1 vssd1 vccd1 vccd1 _13861_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10020__D line[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08320_ _08320_/A _08329_/Y vssd1 vssd1 vccd1 vccd1 _13640_/Z sky130_fd_sc_hd__ebufn_2
X_05532_ _05560_/CLK line[26] vssd1 vssd1 vccd1 vccd1 _05533_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05114__D line[91] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XDATA\[6\].CLKBUF\[1\] clk vssd1 vssd1 vccd1 vccd1 _12842_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__10955__D line[64] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08251_ _08255_/CLK line[103] vssd1 vssd1 vccd1 vccd1 _08252_/A sky130_fd_sc_hd__dfxtp_1
X_05463_ _05463_/A _05494_/Y vssd1 vssd1 vccd1 vccd1 _13863_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_20_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07202_ _07202_/A _07209_/Y vssd1 vssd1 vccd1 vccd1 _13642_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__04953__D line[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08182_ _08182_/A _08189_/Y vssd1 vssd1 vccd1 vccd1 _13782_/Z sky130_fd_sc_hd__ebufn_2
X_05394_ _05420_/CLK line[91] vssd1 vssd1 vccd1 vccd1 _05395_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_192_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07133_ _07135_/CLK line[104] vssd1 vssd1 vccd1 vccd1 _07134_/A sky130_fd_sc_hd__dfxtp_1
X_07064_ _07064_/A _07069_/Y vssd1 vssd1 vccd1 vccd1 _13784_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11786__D line[55] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06015_ _06015_/CLK line[105] vssd1 vssd1 vccd1 vccd1 _06016_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[20\].VALID\[12\].FF OVHB\[20\].V/CLK A[19] vssd1 vssd1 vccd1 vccd1 OVHB\[20\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_161_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09256__D line[50] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09834__A _13921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XOVHB\[9\].VALID\[14\].TOBUF OVHB\[9\].VALID\[14\].FF/Q OVHB\[9\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_199_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09553__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07966_ _07966_/A _07979_/Y vssd1 vssd1 vccd1 vccd1 _13846_/Z sky130_fd_sc_hd__ebufn_2
X_09705_ _09725_/CLK line[14] vssd1 vssd1 vccd1 vccd1 _09706_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[16\].CGAND_B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06917_ _06925_/CLK line[5] vssd1 vssd1 vccd1 vccd1 _06918_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_67_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07897_ _07905_/CLK line[69] vssd1 vssd1 vccd1 vccd1 _07898_/A sky130_fd_sc_hd__dfxtp_1
X_09636_ _09636_/A _09659_/Y vssd1 vssd1 vccd1 vccd1 _13836_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12410__D line[84] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06848_ _06848_/A _06859_/Y vssd1 vssd1 vccd1 vccd1 _13848_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[26\].CLKBUF\[5\] clk vssd1 vssd1 vccd1 vccd1 _10182_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__07504__D line[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09567_ _09585_/CLK line[79] vssd1 vssd1 vccd1 vccd1 _09568_/A sky130_fd_sc_hd__dfxtp_1
X_06779_ _06785_/CLK line[70] vssd1 vssd1 vccd1 vccd1 _06780_/A sky130_fd_sc_hd__dfxtp_1
XPHY_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[20\].VALID\[7\].FF OVHB\[20\].V/CLK A[14] vssd1 vssd1 vccd1 vccd1 OVHB\[20\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08518_ _08518_/A _08539_/Y vssd1 vssd1 vccd1 vccd1 _13838_/Z sky130_fd_sc_hd__ebufn_2
XPHY_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09498_ _09498_/A _09519_/Y vssd1 vssd1 vccd1 vccd1 _13698_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08449_ _08465_/CLK line[65] vssd1 vssd1 vccd1 vccd1 _08450_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[10\].VALID\[14\].FF OVHB\[10\].V/CLK A[21] vssd1 vssd1 vccd1 vccd1 OVHB\[10\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_156_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11460_ _11460_/A _11479_/Y vssd1 vssd1 vccd1 vccd1 _13700_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[29\].VALID\[10\].TOBUF OVHB\[29\].VALID\[10\].FF/Q OVHB\[29\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04932_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_128_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_DATA\[10\].CLKBUF\[6\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10411_ _10425_/CLK line[66] vssd1 vssd1 vccd1 vccd1 _10412_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_139_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[2\].VALID\[13\].TOBUF OVHB\[2\].VALID\[13\].FF/Q OVHB\[2\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04916_/B2 sky130_fd_sc_hd__ebufn_2
X_11391_ _11405_/CLK line[2] vssd1 vssd1 vccd1 vccd1 _11392_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09728__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13130_ _13130_/A _13159_/Y vssd1 vssd1 vccd1 vccd1 _13690_/Z sky130_fd_sc_hd__ebufn_2
X_10342_ _10342_/A _10359_/Y vssd1 vssd1 vccd1 vccd1 _13702_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_164_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11696__D line[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[20\].VALID\[9\].TOBUF OVHB\[20\].VALID\[9\].FF/Q OVHB\[20\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04914_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_2_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13061_ _13085_/CLK line[12] vssd1 vssd1 vccd1 vccd1 _13062_/A sky130_fd_sc_hd__dfxtp_1
X_10273_ _10285_/CLK line[3] vssd1 vssd1 vccd1 vccd1 _10274_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_3_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05694__D line[86] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12012_ _12012_/A _12039_/Y vssd1 vssd1 vccd1 vccd1 _13692_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08070__D line[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13963_ A_h[2] vssd1 vssd1 vccd1 vccd1 _13971_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA_DATA\[3\].CLKBUF\[6\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12320__D line[48] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12914_ _13937_/X vssd1 vssd1 vccd1 vccd1 _12914_/Y sky130_fd_sc_hd__inv_2
X_13894_ _13899_/X vssd1 vssd1 vccd1 vccd1 _13894_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[19\].VALID\[8\].FF OVHB\[19\].V/CLK A[15] vssd1 vssd1 vccd1 vccd1 OVHB\[19\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_12845_ _12875_/CLK line[32] vssd1 vssd1 vccd1 vccd1 _12846_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11514__A _13926_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12776_ _12776_/A _12809_/Y vssd1 vssd1 vccd1 vccd1 _13616_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XDATA\[25\].CLKBUF\[2\] clk vssd1 vssd1 vccd1 vccd1 _09797_/CLK sky130_fd_sc_hd__clkbuf_4
XPHY_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10775__D line[105] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11233__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11727_ _11755_/CLK line[42] vssd1 vssd1 vccd1 vccd1 _11728_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13151__D line[39] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05869__D line[38] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08245__D line[100] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11658_ _11658_/A _11689_/Y vssd1 vssd1 vccd1 vccd1 _13618_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10609_ _10635_/CLK line[43] vssd1 vssd1 vccd1 vccd1 _10610_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11589_ _11615_/CLK line[107] vssd1 vssd1 vccd1 vccd1 _11590_/A sky130_fd_sc_hd__dfxtp_1
X_13328_ _13330_/CLK line[120] vssd1 vssd1 vccd1 vccd1 _13329_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_115_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[11\].VALID\[6\].FF_D A[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13259_ _13259_/A _13264_/Y vssd1 vssd1 vccd1 vccd1 _13819_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09061__TE_B _09064_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MUX.M\[2\].MUX\[3\]_A2 _13809_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07820_ _07820_/A _07839_/Y vssd1 vssd1 vccd1 vccd1 _13700_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09804__D line[59] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07174__A _13909_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07751_ _07765_/CLK line[2] vssd1 vssd1 vccd1 vccd1 _07752_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_111_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11408__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_04963_ _04965_/CLK line[8] vssd1 vssd1 vccd1 vccd1 _04964_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_49_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13326__D line[119] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06702_ _06702_/A _06719_/Y vssd1 vssd1 vccd1 vccd1 _13702_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_37_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07682_ _07682_/A _07699_/Y vssd1 vssd1 vccd1 vccd1 _13842_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_80_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09421_ _09445_/CLK line[12] vssd1 vssd1 vccd1 vccd1 _09422_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_64_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06633_ _06645_/CLK line[3] vssd1 vssd1 vccd1 vccd1 _06634_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[4\].VALID\[1\].TOBUF OVHB\[4\].VALID\[1\].FF/Q OVHB\[4\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04926_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_37_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09352_ _09352_/A _09379_/Y vssd1 vssd1 vccd1 vccd1 _13832_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[29\].VALID\[4\].TOBUF OVHB\[29\].VALID\[4\].FF/Q OVHB\[29\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04925_/B2 sky130_fd_sc_hd__ebufn_2
X_06564_ _06564_/A _06579_/Y vssd1 vssd1 vccd1 vccd1 _13844_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_100_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08303_ _08325_/CLK line[13] vssd1 vssd1 vccd1 vccd1 _08304_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_33_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05515_ _05525_/CLK line[4] vssd1 vssd1 vccd1 vccd1 _05516_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10685__D line[78] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09283_ _09305_/CLK line[77] vssd1 vssd1 vccd1 vccd1 _09284_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13061__D line[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06495_ _06505_/CLK line[68] vssd1 vssd1 vccd1 vccd1 _06496_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05779__D line[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08234_ _08234_/A _08259_/Y vssd1 vssd1 vccd1 vccd1 _13834_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08155__D line[64] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05446_ _05446_/A _05459_/Y vssd1 vssd1 vccd1 vccd1 _13846_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_178_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08165_ _08185_/CLK line[78] vssd1 vssd1 vccd1 vccd1 _08166_/A sky130_fd_sc_hd__dfxtp_1
X_05377_ _05385_/CLK line[69] vssd1 vssd1 vccd1 vccd1 _05378_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07994__D line[113] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_OVHB\[10\].VALID\[14\].FF_D A[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07116_ _07116_/A _07139_/Y vssd1 vssd1 vccd1 vccd1 _13836_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07349__A _13910_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08096_ _08096_/A _08119_/Y vssd1 vssd1 vccd1 vccd1 _13696_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_146_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XDATA\[14\].CLKBUF\[5\] clk vssd1 vssd1 vccd1 vccd1 _06542_/CLK sky130_fd_sc_hd__clkbuf_4
X_07047_ _07065_/CLK line[79] vssd1 vssd1 vccd1 vccd1 _07048_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07068__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08998_ _08998_/A _09029_/Y vssd1 vssd1 vccd1 vccd1 _13758_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_85_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05019__D line[33] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07949_ _07975_/CLK line[107] vssd1 vssd1 vccd1 vccd1 _07950_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_141_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13236__D line[92] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[31\].CGAND_A _13927_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12140__D line[89] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[20\].VALID\[13\].FF_D A[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10960_ _10960_/A _10989_/Y vssd1 vssd1 vccd1 vccd1 _13760_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07234__D line[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09619_ _09619_/A _09624_/Y vssd1 vssd1 vccd1 vccd1 _13819_/Z sky130_fd_sc_hd__ebufn_2
X_10891_ _10915_/CLK line[44] vssd1 vssd1 vccd1 vccd1 _10892_/A sky130_fd_sc_hd__dfxtp_1
XPHY_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12630_ _12630_/CLK line[57] vssd1 vssd1 vccd1 vccd1 _12631_/A sky130_fd_sc_hd__dfxtp_1
XPHY_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[31\].VALID\[2\].FF_D A[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12561_ _12561_/A _12564_/Y vssd1 vssd1 vccd1 vccd1 _13681_/Z sky130_fd_sc_hd__ebufn_2
XPHY_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_DATA\[24\].CLKBUF\[0\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11512_ _11512_/CLK _11513_/X vssd1 vssd1 vccd1 vccd1 _11510_/CLK sky130_fd_sc_hd__dlclkp_1
XPHY_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12492_ _12492_/CLK _12493_/X vssd1 vssd1 vccd1 vccd1 _12490_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__08643__A _13914_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11443_ _13926_/X wr vssd1 vssd1 vccd1 vccd1 _11443_/X sky130_fd_sc_hd__and2_1
XPHY_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[30\].VALID\[12\].FF_D A[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_OVHB\[24\].VALID\[6\].FF_D A[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11374_ _13933_/X vssd1 vssd1 vccd1 vccd1 _11374_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13113_ _13113_/A _13124_/Y vssd1 vssd1 vccd1 vccd1 _13673_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_166_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12315__D line[41] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10325_ _10355_/CLK line[32] vssd1 vssd1 vccd1 vccd1 _10326_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_125_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07409__D line[102] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[29\].VALID\[14\].FF OVHB\[29\].V/CLK A[21] vssd1 vssd1 vccd1 vccd1 OVHB\[29\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_13044_ _13050_/CLK line[118] vssd1 vssd1 vccd1 vccd1 _13045_/A sky130_fd_sc_hd__dfxtp_1
X_10256_ _10256_/A _10289_/Y vssd1 vssd1 vccd1 vccd1 _13616_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_94_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XDATA\[13\].CLKBUF\[2\] clk vssd1 vssd1 vccd1 vccd1 _06157_/CLK sky130_fd_sc_hd__clkbuf_4
X_10187_ _10215_/CLK line[106] vssd1 vssd1 vccd1 vccd1 _10188_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_207_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12050__D line[62] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13946_ _13949_/A _13949_/B _13949_/C _13949_/D vssd1 vssd1 vccd1 vccd1 _13946_/X
+ sky130_fd_sc_hd__and4bb_4
XANTENNA__07144__D line[123] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08818__A _13914_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12985__D line[96] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[12\].VALID\[10\].FF_D A[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13877_ _13877_/A _13894_/Y vssd1 vssd1 vccd1 vccd1 _13877_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06983__D line[35] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12828_ _12840_/CLK line[19] vssd1 vssd1 vccd1 vccd1 _12829_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_188_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[4\].CG clk OVHB\[4\].CGAND/X vssd1 vssd1 vccd1 vccd1 OVHB\[4\].V/CLK sky130_fd_sc_hd__dlclkp_1
X_12759_ _12759_/A _12774_/Y vssd1 vssd1 vccd1 vccd1 _13879_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_148_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05300_ _05300_/A _05319_/Y vssd1 vssd1 vccd1 vccd1 _13700_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11898__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06280_ _06280_/A _06299_/Y vssd1 vssd1 vccd1 vccd1 _13840_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_30_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05231_ _05245_/CLK line[2] vssd1 vssd1 vccd1 vccd1 _05232_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_155_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05162_ _05162_/A _05179_/Y vssd1 vssd1 vccd1 vccd1 _13842_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_116_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09970_ _09970_/CLK line[121] vssd1 vssd1 vccd1 vccd1 _09971_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12225__D line[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05093_ _05105_/CLK line[67] vssd1 vssd1 vccd1 vccd1 _05094_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[2\].VALID\[6\].TOBUF OVHB\[2\].VALID\[6\].FF/Q OVHB\[2\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04923_/A2 sky130_fd_sc_hd__ebufn_2
XANTENNA__07319__D line[75] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08921_ _08921_/A _08924_/Y vssd1 vssd1 vccd1 vccd1 _13681_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06223__D line[72] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[27\].VALID\[9\].TOBUF OVHB\[27\].VALID\[9\].FF/Q OVHB\[27\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04914_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[7\].CG_CLK clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08852_ _08852_/CLK _08853_/X vssd1 vssd1 vccd1 vccd1 _08850_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__10323__A _13923_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09534__D line[49] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07803_ _13912_/X wr vssd1 vssd1 vccd1 vccd1 _07803_/X sky130_fd_sc_hd__and2_1
XANTENNA_MUX.M\[1\].MUX\[4\]_A0 _13622_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08783_ _13914_/X wr vssd1 vssd1 vccd1 vccd1 _08783_/X sky130_fd_sc_hd__and2_1
X_05995_ _06015_/CLK line[110] vssd1 vssd1 vccd1 vccd1 _05996_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[5\].VALID\[1\].FF_D A[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07734_ _13911_/X vssd1 vssd1 vccd1 vccd1 _07734_/Y sky130_fd_sc_hd__inv_2
X_04946_ _04946_/A _04969_/Y vssd1 vssd1 vccd1 vccd1 _13626_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_37_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07665_ _07695_/CLK line[96] vssd1 vssd1 vccd1 vccd1 _07666_/A sky130_fd_sc_hd__dfxtp_1
X_09404_ _09410_/CLK line[118] vssd1 vssd1 vccd1 vccd1 _09405_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[13\].CGAND _13903_/X wr vssd1 vssd1 vccd1 vccd1 OVHB\[13\].CGAND/X sky130_fd_sc_hd__and2_4
X_06616_ _06616_/A _06649_/Y vssd1 vssd1 vccd1 vccd1 _13616_/Z sky130_fd_sc_hd__ebufn_2
X_07596_ _07596_/A _07629_/Y vssd1 vssd1 vccd1 vccd1 _13756_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_111_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09335_ _09335_/A _09344_/Y vssd1 vssd1 vccd1 vccd1 _13815_/Z sky130_fd_sc_hd__ebufn_2
X_06547_ _06575_/CLK line[106] vssd1 vssd1 vccd1 vccd1 _06548_/A sky130_fd_sc_hd__dfxtp_1
X_09266_ _09270_/CLK line[55] vssd1 vssd1 vccd1 vccd1 _09267_/A sky130_fd_sc_hd__dfxtp_1
X_06478_ _06478_/A _06509_/Y vssd1 vssd1 vccd1 vccd1 _13758_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_138_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08217_ _08217_/A _08224_/Y vssd1 vssd1 vccd1 vccd1 _13817_/Z sky130_fd_sc_hd__ebufn_2
X_05429_ _05455_/CLK line[107] vssd1 vssd1 vccd1 vccd1 _05430_/A sky130_fd_sc_hd__dfxtp_1
X_09197_ _09197_/A _09204_/Y vssd1 vssd1 vccd1 vccd1 _13677_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_153_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09709__D line[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08148_ _08150_/CLK line[56] vssd1 vssd1 vccd1 vccd1 _08149_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_119_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08079_ _08079_/A _08084_/Y vssd1 vssd1 vccd1 vccd1 _13679_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_20_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10110_ _10110_/CLK line[57] vssd1 vssd1 vccd1 vccd1 _10111_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_20_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06133__D line[45] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11090_ _11090_/CLK line[121] vssd1 vssd1 vccd1 vccd1 _11091_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11974__D line[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10041_ _10041_/A _10044_/Y vssd1 vssd1 vccd1 vccd1 _13681_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05972__D line[85] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13800_ _13820_/CLK line[94] vssd1 vssd1 vccd1 vccd1 _13801_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13544__A _13898_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11992_ _12000_/CLK line[21] vssd1 vssd1 vccd1 vccd1 _11993_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_29_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13731_ _13731_/A _13754_/Y vssd1 vssd1 vccd1 vccd1 _13731_/Z sky130_fd_sc_hd__ebufn_2
X_10943_ _10943_/A _10954_/Y vssd1 vssd1 vccd1 vccd1 _13743_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13263__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07899__D line[70] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10874_ _10880_/CLK line[22] vssd1 vssd1 vccd1 vccd1 _10875_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_32_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13662_ _13680_/CLK line[31] vssd1 vssd1 vccd1 vccd1 _13663_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06158__A _13903_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[1\].VALID\[14\].FF OVHB\[1\].V/CLK A[21] vssd1 vssd1 vccd1 vccd1 OVHB\[1\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12613_ _12613_/A _12634_/Y vssd1 vssd1 vccd1 vccd1 _13733_/Z sky130_fd_sc_hd__ebufn_2
XPHY_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13593_ _13593_/A _13614_/Y vssd1 vssd1 vccd1 vccd1 _13873_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11214__D line[49] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12544_ _12560_/CLK line[17] vssd1 vssd1 vccd1 vccd1 _12545_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06308__D line[125] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12475_ _12475_/A _12494_/Y vssd1 vssd1 vccd1 vccd1 _13875_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_177_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[4\].V_D TIE/HI vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11426_ _11440_/CLK line[18] vssd1 vssd1 vccd1 vccd1 _11427_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08523__D line[99] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_DATA\[22\].CLKBUF\[2\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13719__A _13899_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11357_ _11357_/A _11374_/Y vssd1 vssd1 vccd1 vccd1 _13877_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[17\].VALID\[14\].FF_D A[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10308_ _10320_/CLK line[19] vssd1 vssd1 vccd1 vccd1 _10309_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_193_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13438__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11288_ _11300_/CLK line[83] vssd1 vssd1 vccd1 vccd1 _11289_/A sky130_fd_sc_hd__dfxtp_1
X_13027_ _13027_/A _13054_/Y vssd1 vssd1 vccd1 vccd1 _13867_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[8\].VALID\[5\].FF OVHB\[8\].V/CLK A[12] vssd1 vssd1 vccd1 vccd1 OVHB\[8\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_10239_ _10239_/A _10254_/Y vssd1 vssd1 vccd1 vccd1 _13879_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05882__D line[58] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05780_ _05780_/A _05809_/Y vssd1 vssd1 vccd1 vccd1 _13620_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_82_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13929_ A[3] vssd1 vssd1 vccd1 vccd1 _13938_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__13604__D line[118] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[27\].VALID\[13\].FF_D A[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07450_ _07450_/CLK line[121] vssd1 vssd1 vccd1 vccd1 _07451_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_62_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06401_ _06401_/A _06404_/Y vssd1 vssd1 vccd1 vccd1 _13681_/Z sky130_fd_sc_hd__ebufn_2
X_07381_ _07381_/A _07384_/Y vssd1 vssd1 vccd1 vccd1 _13821_/Z sky130_fd_sc_hd__ebufn_2
X_09120_ _09130_/CLK line[116] vssd1 vssd1 vccd1 vccd1 _09121_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09379__A _13916_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06332_ _06332_/CLK _06333_/X vssd1 vssd1 vccd1 vccd1 _06330_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__05122__D line[95] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[25\].VALID\[12\].FF OVHB\[25\].V/CLK A[19] vssd1 vssd1 vccd1 vccd1 OVHB\[25\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10963__D line[77] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09051_ _09051_/A _09064_/Y vssd1 vssd1 vccd1 vccd1 _13811_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_175_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09098__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06263_ _13903_/X wr vssd1 vssd1 vccd1 vccd1 _06263_/X sky130_fd_sc_hd__and2_1
XFILLER_129_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08002_ _08010_/CLK line[117] vssd1 vssd1 vccd1 vccd1 _08003_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__04961__D line[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05214_ _13931_/Y vssd1 vssd1 vccd1 vccd1 _05214_/Y sky130_fd_sc_hd__inv_2
X_06194_ _13903_/X vssd1 vssd1 vccd1 vccd1 _06194_/Y sky130_fd_sc_hd__inv_2
X_05145_ _05175_/CLK line[96] vssd1 vssd1 vccd1 vccd1 _05146_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07049__D line[65] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09953_ _09953_/A _09974_/Y vssd1 vssd1 vccd1 vccd1 _13873_/Z sky130_fd_sc_hd__ebufn_2
X_05076_ _05076_/A _05109_/Y vssd1 vssd1 vccd1 vccd1 _13756_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_131_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06888__D line[120] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08904_ _08920_/CLK line[17] vssd1 vssd1 vccd1 vccd1 _08905_/A sky130_fd_sc_hd__dfxtp_1
X_09884_ _09900_/CLK line[81] vssd1 vssd1 vccd1 vccd1 _09885_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_58_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09264__D line[54] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08835_ _08835_/A _08854_/Y vssd1 vssd1 vccd1 vccd1 _13875_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10988__A _13925_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[7\].VOBUF OVHB\[7\].V/Q OVHB\[7\].INV/Y vssd1 vssd1 vccd1 vccd1 _04912_/B1
+ sky130_fd_sc_hd__ebufn_2
XOVHB\[23\].INV _13960_/X vssd1 vssd1 vccd1 vccd1 OVHB\[23\].INV/Y sky130_fd_sc_hd__inv_2
XANTENNA__10203__D line[99] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08766_ _08780_/CLK line[82] vssd1 vssd1 vccd1 vccd1 _08767_/A sky130_fd_sc_hd__dfxtp_1
X_05978_ _05980_/CLK line[88] vssd1 vssd1 vccd1 vccd1 _05979_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_26_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07717_ _07717_/A _07734_/Y vssd1 vssd1 vccd1 vccd1 _13877_/Z sky130_fd_sc_hd__ebufn_2
X_04929_ A_h[17] _04929_/B2 A_h[17] _04929_/B2 vssd1 vssd1 vccd1 vccd1 _04933_/A sky130_fd_sc_hd__a2bb2oi_2
X_08697_ _08697_/A _08714_/Y vssd1 vssd1 vccd1 vccd1 _13737_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[15\].VALID\[14\].FF OVHB\[15\].V/CLK A[21] vssd1 vssd1 vccd1 vccd1 OVHB\[15\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XOVHB\[6\].VALID\[7\].FF OVHB\[6\].V/CLK A[14] vssd1 vssd1 vccd1 vccd1 OVHB\[6\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_26_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13514__D line[91] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07648_ _07660_/CLK line[83] vssd1 vssd1 vccd1 vccd1 _07649_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_14_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07512__D line[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07579_ _07579_/A _07594_/Y vssd1 vssd1 vccd1 vccd1 _13739_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[19\].VALID\[10\].FF_D A[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09318_ _09340_/CLK line[93] vssd1 vssd1 vccd1 vccd1 _09319_/A sky130_fd_sc_hd__dfxtp_1
X_10590_ _10600_/CLK line[20] vssd1 vssd1 vccd1 vccd1 _10591_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[20\].VALID\[9\].FF_D A[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09249_ _09249_/A _09274_/Y vssd1 vssd1 vccd1 vccd1 _13729_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09439__D line[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12260_ _12280_/CLK line[30] vssd1 vssd1 vccd1 vccd1 _12261_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_110_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XOVHB\[15\].VALID\[13\].TOBUF OVHB\[15\].VALID\[13\].FF/Q OVHB\[15\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04916_/B2 sky130_fd_sc_hd__ebufn_2
X_11211_ _11211_/A _11234_/Y vssd1 vssd1 vccd1 vccd1 _13731_/Z sky130_fd_sc_hd__ebufn_2
X_12191_ _12191_/A _12214_/Y vssd1 vssd1 vccd1 vccd1 _13871_/Z sky130_fd_sc_hd__ebufn_2
X_11142_ _11160_/CLK line[31] vssd1 vssd1 vccd1 vccd1 _11143_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_150_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11059__A _13925_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11073_ _11073_/A _11094_/Y vssd1 vssd1 vccd1 vccd1 _13873_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_49_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06798__D line[93] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[9\].VALID\[6\].TOBUF OVHB\[9\].VALID\[6\].FF/Q OVHB\[9\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04923_/A2 sky130_fd_sc_hd__ebufn_2
XANTENNA__09174__D line[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10024_ _10040_/CLK line[17] vssd1 vssd1 vccd1 vccd1 _10025_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_76_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11975_ _11975_/A _12004_/Y vssd1 vssd1 vccd1 vccd1 _13655_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_91_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13714_ _13714_/A _13719_/Y vssd1 vssd1 vccd1 vccd1 _13714_/Z sky130_fd_sc_hd__ebufn_2
X_10926_ _10950_/CLK line[60] vssd1 vssd1 vccd1 vccd1 _10927_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07422__D line[122] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10857_ _10857_/A _10884_/Y vssd1 vssd1 vccd1 vccd1 _13657_/Z sky130_fd_sc_hd__ebufn_2
X_13645_ _13645_/CLK line[9] vssd1 vssd1 vccd1 vccd1 _13646_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_72_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06038__D line[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10788_ _10810_/CLK line[125] vssd1 vssd1 vccd1 vccd1 _10789_/A sky130_fd_sc_hd__dfxtp_1
X_13576_ _13576_/A _13579_/Y vssd1 vssd1 vccd1 vccd1 _13856_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_188_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11879__D line[97] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XOVHB\[4\].VALID\[9\].FF OVHB\[4\].V/CLK A[16] vssd1 vssd1 vccd1 vccd1 OVHB\[4\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_12527_ _12527_/CLK _12528_/X vssd1 vssd1 vccd1 vccd1 _12525_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_8_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MUX.M\[3\].MUX\[5\]_A2 _13799_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09349__D line[107] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08253__D line[104] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12458_ _13935_/X wr vssd1 vssd1 vccd1 vccd1 _12458_/X sky130_fd_sc_hd__and2_1
XFILLER_172_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11409_ _13926_/X vssd1 vssd1 vccd1 vccd1 _11409_/Y sky130_fd_sc_hd__inv_2
X_12389_ _13935_/X vssd1 vssd1 vccd1 vccd1 _12389_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12353__A _13935_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XDATA\[4\].CLKBUF\[6\] clk vssd1 vssd1 vccd1 vccd1 _12457_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_98_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12503__D line[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06950_ _06960_/CLK line[20] vssd1 vssd1 vccd1 vccd1 _06951_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[1\].VALID\[4\].FF_D A[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05901_ _05901_/A _05914_/Y vssd1 vssd1 vccd1 vccd1 _13741_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_79_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06501__D line[71] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06881_ _06881_/A _06894_/Y vssd1 vssd1 vccd1 vccd1 _13881_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[20\].CLKBUF\[4\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11119__D line[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08620_ _08640_/CLK line[30] vssd1 vssd1 vccd1 vccd1 _08621_/A sky130_fd_sc_hd__dfxtp_1
X_05832_ _05840_/CLK line[21] vssd1 vssd1 vccd1 vccd1 _05833_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_67_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09812__D line[63] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MUX.M\[1\].MUX\[1\]_A3 _13856_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08551_ _08551_/A _08574_/Y vssd1 vssd1 vccd1 vccd1 _13871_/Z sky130_fd_sc_hd__ebufn_2
X_05763_ _05763_/A _05774_/Y vssd1 vssd1 vccd1 vccd1 _13883_/Z sky130_fd_sc_hd__ebufn_2
X_07502_ _07520_/CLK line[31] vssd1 vssd1 vccd1 vccd1 _07503_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08428__D line[56] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08482_ _08500_/CLK line[95] vssd1 vssd1 vccd1 vccd1 _08483_/A sky130_fd_sc_hd__dfxtp_1
X_05694_ _05700_/CLK line[86] vssd1 vssd1 vccd1 vccd1 _05695_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[16\].VALID\[1\].TOBUF OVHB\[16\].VALID\[1\].FF/Q OVHB\[16\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04926_/B2 sky130_fd_sc_hd__ebufn_2
X_07433_ _07433_/A _07454_/Y vssd1 vssd1 vccd1 vccd1 _13873_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_211_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12528__A _13936_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07364_ _07380_/CLK line[81] vssd1 vssd1 vccd1 vccd1 _07365_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_210_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09103_ _09103_/A _09134_/Y vssd1 vssd1 vccd1 vccd1 _13863_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10693__D line[67] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06315_ _06315_/A _06334_/Y vssd1 vssd1 vccd1 vccd1 _13875_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_176_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07295_ _07295_/A _07314_/Y vssd1 vssd1 vccd1 vccd1 _13735_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05787__D line[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09034_ _09060_/CLK line[91] vssd1 vssd1 vccd1 vccd1 _09035_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08163__D line[77] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06246_ _06260_/CLK line[82] vssd1 vssd1 vccd1 vccd1 _06247_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_117_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06177_ _06177_/A _06194_/Y vssd1 vssd1 vccd1 vccd1 _13737_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_132_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05128_ _05140_/CLK line[83] vssd1 vssd1 vccd1 vccd1 _05129_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_104_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05059_ _05059_/A _05074_/Y vssd1 vssd1 vccd1 vccd1 _13739_/Z sky130_fd_sc_hd__ebufn_2
X_09936_ _09936_/A _09939_/Y vssd1 vssd1 vccd1 vccd1 _13856_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06411__D line[44] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09867_ _09867_/CLK _09868_/X vssd1 vssd1 vccd1 vccd1 _09865_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__11029__D line[107] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XDATA\[3\].CLKBUF\[3\] clk vssd1 vssd1 vccd1 vccd1 _12072_/CLK sky130_fd_sc_hd__clkbuf_4
X_08818_ _13914_/X wr vssd1 vssd1 vccd1 vccd1 _08818_/X sky130_fd_sc_hd__and2_1
XFILLER_93_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05027__D line[37] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08188__A _13932_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09798_ _13921_/X wr vssd1 vssd1 vccd1 vccd1 _09798_/X sky130_fd_sc_hd__and2_1
XFILLER_45_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10868__D line[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08749_ _13914_/X vssd1 vssd1 vccd1 vccd1 _08749_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13244__D line[81] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[21\].VALID\[10\].FF OVHB\[21\].V/CLK A[17] vssd1 vssd1 vccd1 vccd1 OVHB\[21\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_26_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08338__D line[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11760_ _11790_/CLK line[48] vssd1 vssd1 vccd1 vccd1 _11761_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[16\].VALID\[1\].FF_D A[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10711_ _10711_/A _10744_/Y vssd1 vssd1 vccd1 vccd1 _13791_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11691_ _11691_/A _11724_/Y vssd1 vssd1 vccd1 vccd1 _13651_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10642_ _10670_/CLK line[58] vssd1 vssd1 vccd1 vccd1 _10643_/A sky130_fd_sc_hd__dfxtp_1
X_13430_ _13430_/A _13439_/Y vssd1 vssd1 vccd1 vccd1 _13710_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13361_ _13365_/CLK line[7] vssd1 vssd1 vccd1 vccd1 _13362_/A sky130_fd_sc_hd__dfxtp_1
X_10573_ _10573_/A _10604_/Y vssd1 vssd1 vccd1 vccd1 _13653_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_158_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12312_ _12312_/A _12319_/Y vssd1 vssd1 vccd1 vccd1 _13712_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[13\].VALID\[1\].FF OVHB\[13\].V/CLK A[8] vssd1 vssd1 vccd1 vccd1 OVHB\[13\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_13292_ _13292_/A _13299_/Y vssd1 vssd1 vccd1 vccd1 _13852_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_182_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[22\].VALID\[0\].TOBUF OVHB\[22\].VALID\[0\].FF/Q OVHB\[22\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04924_/B2 sky130_fd_sc_hd__ebufn_2
X_12243_ _12245_/CLK line[8] vssd1 vssd1 vccd1 vccd1 _12244_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10108__D line[56] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XOVHB\[30\].VALID\[5\].FF OVHB\[30\].V/CLK A[12] vssd1 vssd1 vccd1 vccd1 OVHB\[30\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_135_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12174_ _12174_/A _12179_/Y vssd1 vssd1 vccd1 vccd1 _13854_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08801__D line[98] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDATA\[23\].CLKBUF\[7\] clk vssd1 vssd1 vccd1 vccd1 _09412_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__13419__D line[33] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11125_ _11125_/CLK line[9] vssd1 vssd1 vccd1 vccd1 _11126_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_96_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XOVHB\[11\].VALID\[12\].FF OVHB\[11\].V/CLK A[19] vssd1 vssd1 vccd1 vccd1 OVHB\[11\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[19\].CLKBUF\[5\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11056_ _11056_/A _11059_/Y vssd1 vssd1 vccd1 vccd1 _13856_/Z sky130_fd_sc_hd__ebufn_2
X_10007_ _10007_/CLK _10008_/X vssd1 vssd1 vccd1 vccd1 _10005_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_36_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_OVHB\[7\].VALID\[8\].FF_D A[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07152__D line[127] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDATA\[2\].CLKBUF\[0\] clk vssd1 vssd1 vccd1 vccd1 _11127_/CLK sky130_fd_sc_hd__clkbuf_4
X_11958_ _11958_/A _11969_/Y vssd1 vssd1 vccd1 vccd1 _13638_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_83_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12993__D line[109] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10909_ _10915_/CLK line[38] vssd1 vssd1 vccd1 vccd1 _10910_/A sky130_fd_sc_hd__dfxtp_1
X_11889_ _11895_/CLK line[102] vssd1 vssd1 vccd1 vccd1 _11890_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06991__D line[39] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13628_ _13628_/A _13649_/Y vssd1 vssd1 vccd1 vccd1 _13628_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_158_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13559_ _13575_/CLK line[97] vssd1 vssd1 vccd1 vccd1 _13560_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06100_ _06120_/CLK line[30] vssd1 vssd1 vccd1 vccd1 _06101_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09079__D line[97] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07080_ _07100_/CLK line[94] vssd1 vssd1 vccd1 vccd1 _07081_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[29\].VALID\[6\].FF OVHB\[29\].V/CLK A[13] vssd1 vssd1 vccd1 vccd1 OVHB\[29\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__05400__D line[94] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06031_ _06031_/A _06054_/Y vssd1 vssd1 vccd1 vccd1 _13871_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10018__D line[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_MUX.M\[2\].MUX\[6\]_A0 _13675_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XOVHB\[14\].VALID\[6\].TOBUF OVHB\[14\].VALID\[6\].FF/Q OVHB\[14\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04923_/A2 sky130_fd_sc_hd__ebufn_2
XANTENNA__12233__D line[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13907__A A[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07982_ _08010_/CLK line[122] vssd1 vssd1 vccd1 vccd1 _07983_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[11\].VALID\[3\].FF OVHB\[11\].V/CLK A[10] vssd1 vssd1 vccd1 vccd1 OVHB\[11\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07327__D line[79] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09721_ _09725_/CLK line[7] vssd1 vssd1 vccd1 vccd1 _09722_/A sky130_fd_sc_hd__dfxtp_1
X_06933_ _06933_/A _06964_/Y vssd1 vssd1 vccd1 vccd1 _13653_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[8\].INV _13942_/Y vssd1 vssd1 vccd1 vccd1 OVHB\[8\].INV/Y sky130_fd_sc_hd__inv_2
XFILLER_67_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XDATA\[22\].CLKBUF\[4\] clk vssd1 vssd1 vccd1 vccd1 _09027_/CLK sky130_fd_sc_hd__clkbuf_4
X_06864_ _06890_/CLK line[123] vssd1 vssd1 vccd1 vccd1 _06865_/A sky130_fd_sc_hd__dfxtp_1
X_09652_ _09652_/A _09659_/Y vssd1 vssd1 vccd1 vccd1 _13852_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_95_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09542__D line[53] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08603_ _08605_/CLK line[8] vssd1 vssd1 vccd1 vccd1 _08604_/A sky130_fd_sc_hd__dfxtp_1
X_05815_ _05815_/A _05844_/Y vssd1 vssd1 vccd1 vccd1 _13655_/Z sky130_fd_sc_hd__ebufn_2
X_09583_ _09585_/CLK line[72] vssd1 vssd1 vccd1 vccd1 _09584_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[29\].VALID\[1\].FF_D A[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06795_ _06795_/A _06824_/Y vssd1 vssd1 vccd1 vccd1 _13795_/Z sky130_fd_sc_hd__ebufn_2
X_08534_ _08534_/A _08539_/Y vssd1 vssd1 vccd1 vccd1 _13854_/Z sky130_fd_sc_hd__ebufn_2
X_05746_ _05770_/CLK line[124] vssd1 vssd1 vccd1 vccd1 _05747_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_23_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MUX.M\[0\].MUX\[2\]_A1 _13702_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08465_ _08465_/CLK line[73] vssd1 vssd1 vccd1 vccd1 _08466_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05677_ _05677_/A _05704_/Y vssd1 vssd1 vccd1 vccd1 _13797_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_211_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[9\].VALID\[10\].TOBUF OVHB\[9\].VALID\[10\].FF/Q OVHB\[9\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04932_/B2 sky130_fd_sc_hd__ebufn_2
XPHY_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07416_ _07416_/A _07419_/Y vssd1 vssd1 vccd1 vccd1 _13856_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_168_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08396_ _08396_/A _08399_/Y vssd1 vssd1 vccd1 vccd1 _13716_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_196_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07347_ _07347_/CLK _07348_/X vssd1 vssd1 vccd1 vccd1 _07345_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_195_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12408__D line[83] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07278_ _13910_/X wr vssd1 vssd1 vccd1 vccd1 _07278_/X sky130_fd_sc_hd__and2_1
XFILLER_12_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09017_ _09025_/CLK line[69] vssd1 vssd1 vccd1 vccd1 _09018_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13089__A _13938_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06229_ _13903_/X vssd1 vssd1 vccd1 vccd1 _06229_/Y sky130_fd_sc_hd__inv_2
XFILLER_128_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09717__D line[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[27\].VALID\[8\].FF OVHB\[27\].V/CLK A[15] vssd1 vssd1 vccd1 vccd1 OVHB\[27\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06141__D line[34] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09919_ _09935_/CLK line[97] vssd1 vssd1 vccd1 vccd1 _09920_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_120_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11982__D line[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12930_ _12930_/A _12949_/Y vssd1 vssd1 vccd1 vccd1 _13770_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_92_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[6\].VALID\[14\].FF OVHB\[6\].V/CLK A[21] vssd1 vssd1 vccd1 vccd1 OVHB\[6\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__09452__D line[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05980__D line[89] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_206_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10598__D line[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12861_ _12875_/CLK line[34] vssd1 vssd1 vccd1 vccd1 _12862_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_206_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08068__D line[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11812_ _11812_/A _11829_/Y vssd1 vssd1 vccd1 vccd1 _13772_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[20\].VALID\[5\].TOBUF OVHB\[20\].VALID\[5\].FF/Q OVHB\[20\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04927_/B2 sky130_fd_sc_hd__ebufn_2
XDATA\[21\].CLKBUF\[1\] clk vssd1 vssd1 vccd1 vccd1 _08642_/CLK sky130_fd_sc_hd__clkbuf_4
XPHY_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12792_ _12792_/A _12809_/Y vssd1 vssd1 vccd1 vccd1 _13632_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11743_ _11755_/CLK line[35] vssd1 vssd1 vccd1 vccd1 _11744_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XDATA\[11\].CLKBUF\[7\] clk vssd1 vssd1 vccd1 vccd1 _05772_/CLK sky130_fd_sc_hd__clkbuf_4
XPHY_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11674_ _11674_/A _11689_/Y vssd1 vssd1 vccd1 vccd1 _13634_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07700__D line[112] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13413_ _13435_/CLK line[45] vssd1 vssd1 vccd1 vccd1 _13414_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10625_ _10635_/CLK line[36] vssd1 vssd1 vccd1 vccd1 _10626_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11222__D line[53] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13344_ _13344_/A _13369_/Y vssd1 vssd1 vccd1 vccd1 _13624_/Z sky130_fd_sc_hd__ebufn_2
X_10556_ _10556_/A _10569_/Y vssd1 vssd1 vccd1 vccd1 _13636_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06316__D line[114] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10487_ _10495_/CLK line[101] vssd1 vssd1 vccd1 vccd1 _10488_/A sky130_fd_sc_hd__dfxtp_1
X_13275_ _13295_/CLK line[110] vssd1 vssd1 vccd1 vccd1 _13276_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09627__D line[106] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06613__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12226_ _12226_/A _12249_/Y vssd1 vssd1 vccd1 vccd1 _13626_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08531__D line[103] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13149__D line[38] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12157_ _12175_/CLK line[111] vssd1 vssd1 vccd1 vccd1 _12158_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_69_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11108_ _11108_/A _11129_/Y vssd1 vssd1 vccd1 vccd1 _13628_/Z sky130_fd_sc_hd__ebufn_2
X_12088_ _12088_/A _12109_/Y vssd1 vssd1 vccd1 vccd1 _13768_/Z sky130_fd_sc_hd__ebufn_2
X_11039_ _11055_/CLK line[97] vssd1 vssd1 vccd1 vccd1 _11040_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_37_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05890__D line[62] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[17\].CLKBUF\[7\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05600_ _05630_/CLK line[48] vssd1 vssd1 vccd1 vccd1 _05601_/A sky130_fd_sc_hd__dfxtp_1
X_06580_ _06610_/CLK line[112] vssd1 vssd1 vccd1 vccd1 _06581_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_33_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05531_ _05531_/A _05564_/Y vssd1 vssd1 vccd1 vccd1 _13651_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_178_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08250_ _08250_/A _08259_/Y vssd1 vssd1 vccd1 vccd1 _13850_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_33_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08706__D line[55] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05462_ _05490_/CLK line[122] vssd1 vssd1 vccd1 vccd1 _05463_/A sky130_fd_sc_hd__dfxtp_1
X_07201_ _07205_/CLK line[7] vssd1 vssd1 vccd1 vccd1 _07202_/A sky130_fd_sc_hd__dfxtp_1
X_08181_ _08185_/CLK line[71] vssd1 vssd1 vccd1 vccd1 _08182_/A sky130_fd_sc_hd__dfxtp_1
X_05393_ _05393_/A _05424_/Y vssd1 vssd1 vccd1 vccd1 _13793_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11132__D line[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07132_ _07132_/A _07139_/Y vssd1 vssd1 vccd1 vccd1 _13852_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[10\].CLKBUF\[4\] clk vssd1 vssd1 vccd1 vccd1 _05387_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_118_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05130__D line[84] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10971__D line[66] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07063_ _07065_/CLK line[72] vssd1 vssd1 vccd1 vccd1 _07064_/A sky130_fd_sc_hd__dfxtp_1
X_06014_ _06014_/A _06019_/Y vssd1 vssd1 vccd1 vccd1 _13854_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08441__D line[76] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13059__D line[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XOVHB\[29\].VALID\[0\].TOBUF OVHB\[29\].VALID\[0\].FF/Q OVHB\[29\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04924_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_102_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07057__D line[69] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12898__D line[51] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07965_ _07975_/CLK line[100] vssd1 vssd1 vccd1 vccd1 _07966_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_68_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09704_ _09704_/A _09729_/Y vssd1 vssd1 vccd1 vccd1 _13624_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_56_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06916_ _06916_/A _06929_/Y vssd1 vssd1 vccd1 vccd1 _13636_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_68_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07896_ _07896_/A _07909_/Y vssd1 vssd1 vccd1 vccd1 _13776_/Z sky130_fd_sc_hd__ebufn_2
X_09635_ _09655_/CLK line[110] vssd1 vssd1 vccd1 vccd1 _09636_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[12\].VALID\[4\].FF_D A[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06847_ _06855_/CLK line[101] vssd1 vssd1 vccd1 vccd1 _06848_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11307__D line[106] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10211__D line[103] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06778_ _06778_/A _06789_/Y vssd1 vssd1 vccd1 vccd1 _13778_/Z sky130_fd_sc_hd__ebufn_2
X_09566_ _09566_/A _09589_/Y vssd1 vssd1 vccd1 vccd1 _13766_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[25\].VALID\[11\].TOBUF OVHB\[25\].VALID\[11\].FF/Q OVHB\[25\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04915_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__05305__D line[36] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08517_ _08535_/CLK line[111] vssd1 vssd1 vccd1 vccd1 _08518_/A sky130_fd_sc_hd__dfxtp_1
X_05729_ _05735_/CLK line[102] vssd1 vssd1 vccd1 vccd1 _05730_/A sky130_fd_sc_hd__dfxtp_1
XPHY_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09497_ _09515_/CLK line[47] vssd1 vssd1 vccd1 vccd1 _09498_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13522__D line[95] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08616__D line[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08448_ _08448_/A _08469_/Y vssd1 vssd1 vccd1 vccd1 _13768_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07520__D line[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12138__D line[88] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08379_ _08395_/CLK line[33] vssd1 vssd1 vccd1 vccd1 _08380_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10410_ _10410_/A _10429_/Y vssd1 vssd1 vccd1 vccd1 _13770_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_99_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11390_ _11390_/A _11409_/Y vssd1 vssd1 vccd1 vccd1 _13630_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05040__D line[48] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10341_ _10355_/CLK line[34] vssd1 vssd1 vccd1 vccd1 _10342_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_109_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13060_ _13060_/A _13089_/Y vssd1 vssd1 vccd1 vccd1 _13620_/Z sky130_fd_sc_hd__ebufn_2
X_10272_ _10272_/A _10289_/Y vssd1 vssd1 vccd1 vccd1 _13632_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_2_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12011_ _12035_/CLK line[44] vssd1 vssd1 vccd1 vccd1 _12012_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_2_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13962_ A_h[1] vssd1 vssd1 vccd1 vccd1 _13971_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_59_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09182__D line[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12913_ _13937_/X wr vssd1 vssd1 vccd1 vccd1 _12913_/X sky130_fd_sc_hd__and2_1
X_13893_ _13899_/X wr vssd1 vssd1 vccd1 vccd1 _13893_/X sky130_fd_sc_hd__and2_1
XFILLER_73_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10121__D line[76] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12844_ _13937_/X vssd1 vssd1 vccd1 vccd1 _12844_/Y sky130_fd_sc_hd__inv_2
XANTENNA__05215__D line[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12775_ _12805_/CLK line[0] vssd1 vssd1 vccd1 vccd1 _12776_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11726_ _11726_/A _11759_/Y vssd1 vssd1 vccd1 vccd1 _13686_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07430__D line[126] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[4\].VALID\[13\].FF_D A[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12048__D line[61] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11657_ _11685_/CLK line[10] vssd1 vssd1 vccd1 vccd1 _11658_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10608_ _10608_/A _10639_/Y vssd1 vssd1 vccd1 vccd1 _13688_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06046__D line[119] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11588_ _11588_/A _11619_/Y vssd1 vssd1 vccd1 vccd1 _13828_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11887__D line[101] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13327_ _13327_/A _13334_/Y vssd1 vssd1 vccd1 vccd1 _13887_/Z sky130_fd_sc_hd__ebufn_2
X_10539_ _10565_/CLK line[11] vssd1 vssd1 vccd1 vccd1 _10540_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09357__D line[111] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XOVHB\[2\].VALID\[12\].FF OVHB\[2\].V/CLK A[19] vssd1 vssd1 vccd1 vccd1 OVHB\[2\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_13258_ _13260_/CLK line[88] vssd1 vssd1 vccd1 vccd1 _13259_/A sky130_fd_sc_hd__dfxtp_1
X_12209_ _12209_/A _12214_/Y vssd1 vssd1 vccd1 vccd1 _13889_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.M\[2\].MUX\[3\]_A3 _13879_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13189_ _13189_/A _13194_/Y vssd1 vssd1 vccd1 vccd1 _13749_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_123_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__04929__B1 A_h[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[25\].VALID\[4\].FF_D A[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12511__D line[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_04962_ _04962_/A _04969_/Y vssd1 vssd1 vccd1 vccd1 _13642_/Z sky130_fd_sc_hd__ebufn_2
X_07750_ _07750_/A _07769_/Y vssd1 vssd1 vccd1 vccd1 _13630_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07605__D line[78] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06701_ _06715_/CLK line[34] vssd1 vssd1 vccd1 vccd1 _06702_/A sky130_fd_sc_hd__dfxtp_1
X_07681_ _07695_/CLK line[98] vssd1 vssd1 vccd1 vccd1 _07682_/A sky130_fd_sc_hd__dfxtp_1
X_09420_ _09420_/A _09449_/Y vssd1 vssd1 vccd1 vccd1 _13620_/Z sky130_fd_sc_hd__ebufn_2
X_06632_ _06632_/A _06649_/Y vssd1 vssd1 vccd1 vccd1 _13632_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09820__D line[52] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[2\].VALID\[2\].TOBUF OVHB\[2\].VALID\[2\].FF/Q OVHB\[2\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04930_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__05703__A _13901_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09351_ _09375_/CLK line[108] vssd1 vssd1 vccd1 vccd1 _09352_/A sky130_fd_sc_hd__dfxtp_1
X_06563_ _06575_/CLK line[99] vssd1 vssd1 vccd1 vccd1 _06564_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[18\].VALID\[8\].FF_D A[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[27\].VALID\[5\].TOBUF OVHB\[27\].VALID\[5\].FF/Q OVHB\[27\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04927_/B2 sky130_fd_sc_hd__ebufn_2
X_05514_ _05514_/A _05529_/Y vssd1 vssd1 vccd1 vccd1 _13634_/Z sky130_fd_sc_hd__ebufn_2
X_08302_ _08302_/A _08329_/Y vssd1 vssd1 vccd1 vccd1 _13622_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09282_ _09282_/A _09309_/Y vssd1 vssd1 vccd1 vccd1 _13762_/Z sky130_fd_sc_hd__ebufn_2
X_06494_ _06494_/A _06509_/Y vssd1 vssd1 vccd1 vccd1 _13774_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_20_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08233_ _08255_/CLK line[109] vssd1 vssd1 vccd1 vccd1 _08234_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_193_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05445_ _05455_/CLK line[100] vssd1 vssd1 vccd1 vccd1 _05446_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_20_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08164_ _08164_/A _08189_/Y vssd1 vssd1 vccd1 vccd1 _13764_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_118_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05376_ _05376_/A _05389_/Y vssd1 vssd1 vccd1 vccd1 _13776_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[0\].VALID\[0\].FF OVHB\[0\].V/CLK A[7] vssd1 vssd1 vccd1 vccd1 OVHB\[0\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11797__D line[74] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MUX.SEL1BUF\[3\]_A A[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07115_ _07135_/CLK line[110] vssd1 vssd1 vccd1 vccd1 _07116_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[11\].CLKBUF\[0\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08095_ _08115_/CLK line[46] vssd1 vssd1 vccd1 vccd1 _08096_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_161_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05795__D line[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08171__D line[66] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07046_ _07046_/A _07069_/Y vssd1 vssd1 vccd1 vccd1 _13766_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_161_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[26\].VALID\[10\].FF OVHB\[26\].V/CLK A[17] vssd1 vssd1 vccd1 vccd1 OVHB\[26\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_08997_ _09025_/CLK line[74] vssd1 vssd1 vccd1 vccd1 _08998_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_85_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07948_ _07948_/A _07979_/Y vssd1 vssd1 vccd1 vccd1 _13828_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[31\].CGAND_B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07879_ _07905_/CLK line[75] vssd1 vssd1 vccd1 vccd1 _07880_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11037__D line[111] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09618_ _09620_/CLK line[88] vssd1 vssd1 vccd1 vccd1 _09619_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_18_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_DATA\[4\].CLKBUF\[0\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05035__D line[41] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10890_ _10890_/A _10919_/Y vssd1 vssd1 vccd1 vccd1 _13690_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09730__D line[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10876__D line[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09549_ _09549_/A _09554_/Y vssd1 vssd1 vccd1 vccd1 _13749_/Z sky130_fd_sc_hd__ebufn_2
XPHY_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13252__D line[85] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12560_ _12560_/CLK line[25] vssd1 vssd1 vccd1 vccd1 _12561_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08346__D line[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08924__A _13915_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_DATA\[30\].CLKBUF\[2\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11511_ _11511_/A _11514_/Y vssd1 vssd1 vccd1 vccd1 _13751_/Z sky130_fd_sc_hd__ebufn_2
XPHY_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12491_ _12491_/A _12494_/Y vssd1 vssd1 vccd1 vccd1 _13891_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08643__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11442_ _11442_/CLK _11443_/X vssd1 vssd1 vccd1 vccd1 _11440_/CLK sky130_fd_sc_hd__dlclkp_1
XPHY_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[16\].VALID\[12\].FF OVHB\[16\].V/CLK A[19] vssd1 vssd1 vccd1 vccd1 OVHB\[16\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_11373_ _13933_/X wr vssd1 vssd1 vccd1 vccd1 _11373_/X sky130_fd_sc_hd__and2_1
XANTENNA__11500__D line[52] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13112_ _13120_/CLK line[21] vssd1 vssd1 vccd1 vccd1 _13113_/A sky130_fd_sc_hd__dfxtp_1
X_10324_ _13923_/X vssd1 vssd1 vccd1 vccd1 _10324_/Y sky130_fd_sc_hd__inv_2
X_10255_ _10285_/CLK line[0] vssd1 vssd1 vccd1 vccd1 _10256_/A sky130_fd_sc_hd__dfxtp_1
X_13043_ _13043_/A _13054_/Y vssd1 vssd1 vccd1 vccd1 _13883_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_59_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09905__D line[96] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10186_ _10186_/A _10219_/Y vssd1 vssd1 vccd1 vccd1 _13826_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13427__D line[37] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__04927__A1_N A_h[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13945_ _13949_/C _13949_/B _13949_/A _13949_/D vssd1 vssd1 vccd1 vccd1 _13945_/X
+ sky130_fd_sc_hd__and4b_4
XANTENNA__08818__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13876_ _13890_/CLK line[114] vssd1 vssd1 vccd1 vccd1 _13877_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_201_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10786__D line[124] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12827_ _12827_/A _12844_/Y vssd1 vssd1 vccd1 vccd1 _13667_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_22_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13162__D line[58] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12758_ _12770_/CLK line[115] vssd1 vssd1 vccd1 vccd1 _12759_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07160__D line[116] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11709_ _11709_/A _11724_/Y vssd1 vssd1 vccd1 vccd1 _13669_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_175_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12689_ _12689_/A _12704_/Y vssd1 vssd1 vccd1 vccd1 _13809_/Z sky130_fd_sc_hd__ebufn_2
X_05230_ _05230_/A _05249_/Y vssd1 vssd1 vccd1 vccd1 _13630_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_190_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05161_ _05175_/CLK line[98] vssd1 vssd1 vccd1 vccd1 _05162_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11410__D line[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09087__D line[101] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05092_ _05092_/A _05109_/Y vssd1 vssd1 vccd1 vccd1 _13772_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[0\].VALID\[7\].TOBUF OVHB\[0\].VALID\[7\].FF/Q OVHB\[0\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/A2 sky130_fd_sc_hd__ebufn_2
XANTENNA__10026__D line[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08920_ _08920_/CLK line[25] vssd1 vssd1 vccd1 vccd1 _08921_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10604__A _13924_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08851_ _08851_/A _08854_/Y vssd1 vssd1 vccd1 vccd1 _13891_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_111_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13337__D line[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10323__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07802_ _07802_/CLK _07803_/X vssd1 vssd1 vccd1 vccd1 _07800_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__12241__D line[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__04959__D line[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08782_ _08782_/CLK _08783_/X vssd1 vssd1 vccd1 vccd1 _08780_/CLK sky130_fd_sc_hd__dlclkp_1
X_05994_ _05994_/A _06019_/Y vssd1 vssd1 vccd1 vccd1 _13834_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.M\[1\].MUX\[4\]_A1 _13692_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07335__D line[68] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_04945_ _04965_/CLK line[14] vssd1 vssd1 vccd1 vccd1 _04946_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_84_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07733_ _13911_/X wr vssd1 vssd1 vccd1 vccd1 _07733_/X sky130_fd_sc_hd__and2_1
XFILLER_37_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07664_ _13911_/X vssd1 vssd1 vccd1 vccd1 _07664_/Y sky130_fd_sc_hd__inv_2
XANTENNA__09550__D line[57] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09403_ _09403_/A _09414_/Y vssd1 vssd1 vccd1 vccd1 _13883_/Z sky130_fd_sc_hd__ebufn_2
X_06615_ _06645_/CLK line[0] vssd1 vssd1 vccd1 vccd1 _06616_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_13_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07595_ _07625_/CLK line[64] vssd1 vssd1 vccd1 vccd1 _07596_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[29\].CLKBUF\[3\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09334_ _09340_/CLK line[86] vssd1 vssd1 vccd1 vccd1 _09335_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_40_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06546_ _06546_/A _06579_/Y vssd1 vssd1 vccd1 vccd1 _13826_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07070__D line[80] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06477_ _06505_/CLK line[74] vssd1 vssd1 vccd1 vccd1 _06478_/A sky130_fd_sc_hd__dfxtp_1
X_09265_ _09265_/A _09274_/Y vssd1 vssd1 vccd1 vccd1 _13745_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_178_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13800__D line[94] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05428_ _05428_/A _05459_/Y vssd1 vssd1 vccd1 vccd1 _13828_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_138_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08216_ _08220_/CLK line[87] vssd1 vssd1 vccd1 vccd1 _08217_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[3\].VOBUF OVHB\[3\].V/Q OVHB\[3\].INV/Y vssd1 vssd1 vccd1 vccd1 _04912_/B1
+ sky130_fd_sc_hd__ebufn_2
X_09196_ _09200_/CLK line[23] vssd1 vssd1 vccd1 vccd1 _09197_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06264__A _13903_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05359_ _05385_/CLK line[75] vssd1 vssd1 vccd1 vccd1 _05360_/A sky130_fd_sc_hd__dfxtp_1
X_08147_ _08147_/A _08154_/Y vssd1 vssd1 vccd1 vccd1 _13747_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12416__D line[87] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08078_ _08080_/CLK line[24] vssd1 vssd1 vccd1 vccd1 _08079_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_20_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07029_ _07029_/A _07034_/Y vssd1 vssd1 vccd1 vccd1 _13749_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09725__D line[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10040_ _10040_/CLK line[25] vssd1 vssd1 vccd1 vccd1 _10041_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12151__D line[108] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07245__D line[32] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XDATA\[31\].CLKBUF\[6\] clk vssd1 vssd1 vccd1 vccd1 _11897_/CLK sky130_fd_sc_hd__clkbuf_4
X_11991_ _11991_/A _12004_/Y vssd1 vssd1 vccd1 vccd1 _13671_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11990__D line[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13730_ _13750_/CLK line[62] vssd1 vssd1 vccd1 vccd1 _13731_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_28_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10942_ _10950_/CLK line[53] vssd1 vssd1 vccd1 vccd1 _10943_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06439__A _13904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09460__D line[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13661_ _13661_/A _13684_/Y vssd1 vssd1 vccd1 vccd1 _13661_/Z sky130_fd_sc_hd__ebufn_2
X_10873_ _10873_/A _10884_/Y vssd1 vssd1 vccd1 vccd1 _13673_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06158__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[31\].VALID\[9\].TOBUF OVHB\[31\].VALID\[9\].FF/Q OVHB\[31\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04914_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__08076__D line[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12612_ _12630_/CLK line[63] vssd1 vssd1 vccd1 vccd1 _12613_/A sky130_fd_sc_hd__dfxtp_1
XPHY_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13592_ _13610_/CLK line[127] vssd1 vssd1 vccd1 vccd1 _13593_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_101_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[9\].VALID\[2\].TOBUF OVHB\[9\].VALID\[2\].FF/Q OVHB\[9\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04930_/B2 sky130_fd_sc_hd__ebufn_2
XPHY_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12543_ _12543_/A _12564_/Y vssd1 vssd1 vccd1 vccd1 _13663_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_157_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_DATA\[2\].CLKBUF\[2\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12474_ _12490_/CLK line[113] vssd1 vssd1 vccd1 vccd1 _12475_/A sky130_fd_sc_hd__dfxtp_1
X_11425_ _11425_/A _11444_/Y vssd1 vssd1 vccd1 vccd1 _13665_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12326__D line[60] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11230__D line[57] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDATA\[0\].CLKBUF\[5\] clk vssd1 vssd1 vccd1 vccd1 _05142_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_153_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06324__D line[118] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11356_ _11370_/CLK line[114] vssd1 vssd1 vccd1 vccd1 _11357_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_140_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10307_ _10307_/A _10324_/Y vssd1 vssd1 vccd1 vccd1 _13667_/Z sky130_fd_sc_hd__ebufn_2
X_11287_ _11287_/A _11304_/Y vssd1 vssd1 vccd1 vccd1 _13807_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09635__D line[110] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[21\].VALID\[7\].FF_D A[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13026_ _13050_/CLK line[124] vssd1 vssd1 vccd1 vccd1 _13027_/A sky130_fd_sc_hd__dfxtp_1
X_10238_ _10250_/CLK line[115] vssd1 vssd1 vccd1 vccd1 _10239_/A sky130_fd_sc_hd__dfxtp_1
X_10169_ _10169_/A _10184_/Y vssd1 vssd1 vccd1 vccd1 _13809_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_120_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07733__A _13911_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[27\].CG_CLK clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13928_ A[2] vssd1 vssd1 vccd1 vccd1 _13938_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_34_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13859_ _13899_/X vssd1 vssd1 vccd1 vccd1 _13859_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11405__D line[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06400_ _06400_/CLK line[25] vssd1 vssd1 vccd1 vccd1 _06401_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[30\].CLKBUF\[3\] clk vssd1 vssd1 vccd1 vccd1 _11512_/CLK sky130_fd_sc_hd__clkbuf_4
XOVHB\[12\].VALID\[10\].FF OVHB\[12\].V/CLK A[17] vssd1 vssd1 vccd1 vccd1 OVHB\[12\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_34_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07380_ _07380_/CLK line[89] vssd1 vssd1 vccd1 vccd1 _07381_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_210_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06331_ _06331_/A _06334_/Y vssd1 vssd1 vccd1 vccd1 _13891_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_148_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_187_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09050_ _09060_/CLK line[84] vssd1 vssd1 vccd1 vccd1 _09051_/A sky130_fd_sc_hd__dfxtp_1
X_06262_ _06262_/CLK _06263_/X vssd1 vssd1 vccd1 vccd1 _06260_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_191_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08001_ _08001_/A _08014_/Y vssd1 vssd1 vccd1 vccd1 _13881_/Z sky130_fd_sc_hd__ebufn_2
X_05213_ _13931_/Y wr vssd1 vssd1 vccd1 vccd1 _05213_/X sky130_fd_sc_hd__and2_1
X_06193_ _13903_/X wr vssd1 vssd1 vccd1 vccd1 _06193_/X sky130_fd_sc_hd__and2_1
XFILLER_128_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11140__D line[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05144_ _13931_/Y vssd1 vssd1 vccd1 vccd1 _05144_/Y sky130_fd_sc_hd__inv_2
XANTENNA__07908__A _13912_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06234__D line[91] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMUX.SEL1BUF\[2\] A[1] vssd1 vssd1 vccd1 vccd1 MUX.SEL1BUF\[2\]/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09952_ _09970_/CLK line[127] vssd1 vssd1 vccd1 vccd1 _09953_/A sky130_fd_sc_hd__dfxtp_1
X_05075_ _05105_/CLK line[64] vssd1 vssd1 vccd1 vccd1 _05076_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_98_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08903_ _08903_/A _08924_/Y vssd1 vssd1 vccd1 vccd1 _13663_/Z sky130_fd_sc_hd__ebufn_2
X_09883_ _09883_/A _09904_/Y vssd1 vssd1 vccd1 vccd1 _13803_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13067__D line[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08834_ _08850_/CLK line[113] vssd1 vssd1 vccd1 vccd1 _08835_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_112_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07065__D line[73] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10988__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08765_ _08765_/A _08784_/Y vssd1 vssd1 vccd1 vccd1 _13805_/Z sky130_fd_sc_hd__ebufn_2
X_05977_ _05977_/A _05984_/Y vssd1 vssd1 vccd1 vccd1 _13817_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_38_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07716_ _07730_/CLK line[114] vssd1 vssd1 vccd1 vccd1 _07717_/A sky130_fd_sc_hd__dfxtp_1
X_04928_ _04928_/A _04928_/B _04928_/C _04928_/D vssd1 vssd1 vccd1 vccd1 _04934_/C
+ sky130_fd_sc_hd__or4_2
X_08696_ _08710_/CLK line[50] vssd1 vssd1 vccd1 vccd1 _08697_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_81_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[21\].VALID\[14\].FF_D A[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07647_ _07647_/A _07664_/Y vssd1 vssd1 vccd1 vccd1 _13807_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_202_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11315__D line[110] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[2\].VALID\[2\].FF_D A[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[21\].VALID\[1\].FF OVHB\[21\].V/CLK A[8] vssd1 vssd1 vccd1 vccd1 OVHB\[21\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06409__D line[43] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05313__D line[40] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07578_ _07590_/CLK line[51] vssd1 vssd1 vccd1 vccd1 _07579_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_22_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XOVHB\[11\].VALID\[14\].TOBUF OVHB\[11\].VALID\[14\].FF/Q OVHB\[11\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/B2 sky130_fd_sc_hd__ebufn_2
X_09317_ _09317_/A _09344_/Y vssd1 vssd1 vccd1 vccd1 _13797_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_40_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06529_ _06529_/A _06544_/Y vssd1 vssd1 vccd1 vccd1 _13809_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13530__D line[84] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08624__D line[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09248_ _09270_/CLK line[61] vssd1 vssd1 vccd1 vccd1 _09249_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[27\].CLKBUF\[5\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09179_ _09179_/A _09204_/Y vssd1 vssd1 vccd1 vccd1 _13659_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_166_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XOVHB\[22\].CG clk OVHB\[22\].CGAND/X vssd1 vssd1 vccd1 vccd1 OVHB\[22\].V/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_147_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11210_ _11230_/CLK line[62] vssd1 vssd1 vccd1 vccd1 _11211_/A sky130_fd_sc_hd__dfxtp_1
X_12190_ _12210_/CLK line[126] vssd1 vssd1 vccd1 vccd1 _12191_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[31\].VALID\[13\].FF_D A[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11141_ _11141_/A _11164_/Y vssd1 vssd1 vccd1 vccd1 _13661_/Z sky130_fd_sc_hd__ebufn_2
X_11072_ _11090_/CLK line[127] vssd1 vssd1 vccd1 vccd1 _11073_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_1_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10023_ _10023_/A _10044_/Y vssd1 vssd1 vccd1 vccd1 _13663_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[7\].VALID\[7\].TOBUF OVHB\[7\].VALID\[7\].FF/Q OVHB\[7\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/A2 sky130_fd_sc_hd__ebufn_2
XFILLER_1_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13705__D line[36] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11974_ _12000_/CLK line[27] vssd1 vssd1 vccd1 vccd1 _11975_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_16_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09190__D line[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05073__A _13931_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13713_ _13715_/CLK line[40] vssd1 vssd1 vccd1 vccd1 _13714_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_16_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10925_ _10925_/A _10954_/Y vssd1 vssd1 vccd1 vccd1 _13725_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_204_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[13\].VALID\[11\].FF_D A[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13644_ _13644_/A _13649_/Y vssd1 vssd1 vccd1 vccd1 _13644_/Z sky130_fd_sc_hd__ebufn_2
X_10856_ _10880_/CLK line[28] vssd1 vssd1 vccd1 vccd1 _10857_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_72_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05223__D line[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13575_ _13575_/CLK line[105] vssd1 vssd1 vccd1 vccd1 _13576_/A sky130_fd_sc_hd__dfxtp_1
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10787_ _10787_/A _10814_/Y vssd1 vssd1 vccd1 vccd1 _13867_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13440__D line[48] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XOVHB\[7\].VALID\[12\].FF OVHB\[7\].V/CLK A[19] vssd1 vssd1 vccd1 vccd1 OVHB\[7\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12526_ _12526_/A _12529_/Y vssd1 vssd1 vccd1 vccd1 _13646_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_118_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MUX.M\[3\].MUX\[5\]_A3 _13869_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12056__D line[50] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12457_ _12457_/CLK _12458_/X vssd1 vssd1 vccd1 vccd1 _12455_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__12634__A _13936_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11408_ _13926_/X wr vssd1 vssd1 vccd1 vccd1 _11408_/X sky130_fd_sc_hd__and2_1
XFILLER_126_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12388_ _13935_/X wr vssd1 vssd1 vccd1 vccd1 _12388_/X sky130_fd_sc_hd__and2_1
XANTENNA__11895__D line[105] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12353__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[0\].V OVHB\[0\].V/CLK TIE/HI rst_n vssd1 vssd1 vccd1 vccd1 OVHB\[0\].V/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_DATA\[0\].CLKBUF\[4\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06989__D line[38] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11339_ _13933_/X vssd1 vssd1 vccd1 vccd1 _11339_/Y sky130_fd_sc_hd__inv_2
XANTENNA_OVHB\[23\].VALID\[10\].FF_D A[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09365__D line[100] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05248__A _13900_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10304__D line[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05900_ _05910_/CLK line[52] vssd1 vssd1 vccd1 vccd1 _05901_/A sky130_fd_sc_hd__dfxtp_1
X_13009_ _13015_/CLK line[102] vssd1 vssd1 vccd1 vccd1 _13010_/A sky130_fd_sc_hd__dfxtp_1
X_06880_ _06890_/CLK line[116] vssd1 vssd1 vccd1 vccd1 _06881_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05831_ _05831_/A _05844_/Y vssd1 vssd1 vccd1 vccd1 _13671_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[31\].VALID\[14\].TOBUF OVHB\[31\].VALID\[14\].FF/Q OVHB\[31\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_55_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13615__D line[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08550_ _08570_/CLK line[126] vssd1 vssd1 vccd1 vccd1 _08551_/A sky130_fd_sc_hd__dfxtp_1
X_05762_ _05770_/CLK line[117] vssd1 vssd1 vccd1 vccd1 _05763_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07613__D line[67] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07501_ _07501_/A _07524_/Y vssd1 vssd1 vccd1 vccd1 _13661_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_63_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05693_ _05693_/A _05704_/Y vssd1 vssd1 vccd1 vccd1 _13813_/Z sky130_fd_sc_hd__ebufn_2
X_08481_ _08481_/A _08504_/Y vssd1 vssd1 vccd1 vccd1 _13801_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12809__A _13937_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07432_ _07450_/CLK line[127] vssd1 vssd1 vccd1 vccd1 _07433_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[14\].VALID\[2\].TOBUF OVHB\[14\].VALID\[2\].FF/Q OVHB\[14\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04930_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__08294__A _13932_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12528__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07363_ _07363_/A _07384_/Y vssd1 vssd1 vccd1 vccd1 _13803_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[8\].VALID\[6\].FF_D A[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09102_ _09130_/CLK line[122] vssd1 vssd1 vccd1 vccd1 _09103_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__04972__D line[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06314_ _06330_/CLK line[113] vssd1 vssd1 vccd1 vccd1 _06315_/A sky130_fd_sc_hd__dfxtp_1
X_07294_ _07310_/CLK line[49] vssd1 vssd1 vccd1 vccd1 _07295_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_136_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XOVHB\[18\].VALID\[4\].FF OVHB\[18\].V/CLK A[11] vssd1 vssd1 vccd1 vccd1 OVHB\[18\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_09033_ _09033_/A _09064_/Y vssd1 vssd1 vccd1 vccd1 _13793_/Z sky130_fd_sc_hd__ebufn_2
X_06245_ _06245_/A _06264_/Y vssd1 vssd1 vccd1 vccd1 _13805_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_129_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06176_ _06190_/CLK line[50] vssd1 vssd1 vccd1 vccd1 _06177_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_132_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05127_ _05127_/A _05144_/Y vssd1 vssd1 vccd1 vccd1 _13807_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06899__D line[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09275__D line[64] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05058_ _05070_/CLK line[51] vssd1 vssd1 vccd1 vccd1 _05059_/A sky130_fd_sc_hd__dfxtp_1
X_09935_ _09935_/CLK line[105] vssd1 vssd1 vccd1 vccd1 _09936_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_131_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09866_ _09866_/A _09869_/Y vssd1 vssd1 vccd1 vccd1 _13786_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08469__A _13913_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08817_ _08817_/CLK _08818_/X vssd1 vssd1 vccd1 vccd1 _08815_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_85_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09797_ _09797_/CLK _09798_/X vssd1 vssd1 vccd1 vccd1 _09795_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__08188__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[3\].V_D TIE/HI vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08748_ _13914_/X wr vssd1 vssd1 vccd1 vccd1 _08748_/X sky130_fd_sc_hd__and2_1
XFILLER_26_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08679_ _13914_/X vssd1 vssd1 vccd1 vccd1 _08679_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11045__D line[100] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10710_ _10740_/CLK line[80] vssd1 vssd1 vccd1 vccd1 _10711_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_26_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06139__D line[33] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11690_ _11720_/CLK line[16] vssd1 vssd1 vccd1 vccd1 _11691_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10641_ _10641_/A _10674_/Y vssd1 vssd1 vccd1 vccd1 _13721_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05978__D line[88] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13260__D line[89] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13360_ _13360_/A _13369_/Y vssd1 vssd1 vccd1 vccd1 _13640_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08354__D line[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10572_ _10600_/CLK line[26] vssd1 vssd1 vccd1 vccd1 _10573_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_158_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12311_ _12315_/CLK line[39] vssd1 vssd1 vccd1 vccd1 _12312_/A sky130_fd_sc_hd__dfxtp_1
X_13291_ _13295_/CLK line[103] vssd1 vssd1 vccd1 vccd1 _13292_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_158_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12242_ _12242_/A _12249_/Y vssd1 vssd1 vccd1 vccd1 _13642_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[20\].VALID\[1\].TOBUF OVHB\[20\].VALID\[1\].FF/Q OVHB\[20\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04926_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__12604__D line[59] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12173_ _12175_/CLK line[104] vssd1 vssd1 vccd1 vccd1 _12174_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_3_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XOVHB\[16\].VALID\[6\].FF OVHB\[16\].V/CLK A[13] vssd1 vssd1 vccd1 vccd1 OVHB\[16\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_11124_ _11124_/A _11129_/Y vssd1 vssd1 vccd1 vccd1 _13644_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09763__A _13921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06602__D line[117] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[25\].CLKBUF\[7\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11055_ _11055_/CLK line[105] vssd1 vssd1 vccd1 vccd1 _11056_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09913__D line[109] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10006_ _10006_/A _10009_/Y vssd1 vssd1 vccd1 vccd1 _13646_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13435__D line[41] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08529__D line[102] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11957_ _11965_/CLK line[5] vssd1 vssd1 vccd1 vccd1 _11958_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_205_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10908_ _10908_/A _10919_/Y vssd1 vssd1 vccd1 vccd1 _13708_/Z sky130_fd_sc_hd__ebufn_2
X_11888_ _11888_/A _11899_/Y vssd1 vssd1 vccd1 vccd1 _13848_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[28\].VALID\[14\].FF_D A[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10794__D line[113] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13627_ _13645_/CLK line[15] vssd1 vssd1 vccd1 vccd1 _13628_/A sky130_fd_sc_hd__dfxtp_1
X_10839_ _10845_/CLK line[6] vssd1 vssd1 vccd1 vccd1 _10840_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10149__A _13922_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13170__D line[62] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05888__D line[61] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08264__D line[123] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09938__A _13921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13558_ _13558_/A _13579_/Y vssd1 vssd1 vccd1 vccd1 _13838_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_192_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12509_ _12525_/CLK line[1] vssd1 vssd1 vccd1 vccd1 _12510_/A sky130_fd_sc_hd__dfxtp_1
X_13489_ _13505_/CLK line[65] vssd1 vssd1 vccd1 vccd1 _13490_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[22\].INV _13959_/X vssd1 vssd1 vccd1 vccd1 OVHB\[22\].INV/Y sky130_fd_sc_hd__inv_2
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06030_ _06050_/CLK line[126] vssd1 vssd1 vccd1 vccd1 _06031_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.M\[2\].MUX\[6\]_A1 _13745_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09095__D line[105] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06512__D line[90] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[12\].VALID\[7\].TOBUF OVHB\[12\].VALID\[7\].FF/Q OVHB\[12\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/A2 sky130_fd_sc_hd__ebufn_2
X_07981_ _07981_/A _08014_/Y vssd1 vssd1 vccd1 vccd1 _13861_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10034__D line[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09720_ _09720_/A _09729_/Y vssd1 vssd1 vccd1 vccd1 _13640_/Z sky130_fd_sc_hd__ebufn_2
X_06932_ _06960_/CLK line[26] vssd1 vssd1 vccd1 vccd1 _06933_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05128__D line[83] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09651_ _09655_/CLK line[103] vssd1 vssd1 vccd1 vccd1 _09652_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10969__D line[65] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[31\].V_RESET_B rst_n vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06863_ _06863_/A _06894_/Y vssd1 vssd1 vccd1 vccd1 _13863_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_94_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[5\].VALID\[11\].TOBUF OVHB\[5\].VALID\[11\].FF/Q OVHB\[5\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04915_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__13345__D line[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08602_ _08602_/A _08609_/Y vssd1 vssd1 vccd1 vccd1 _13642_/Z sky130_fd_sc_hd__ebufn_2
X_05814_ _05840_/CLK line[27] vssd1 vssd1 vccd1 vccd1 _05815_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_103_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08439__D line[75] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09582_ _09582_/A _09589_/Y vssd1 vssd1 vccd1 vccd1 _13782_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07343__D line[72] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XOVHB\[14\].VALID\[8\].FF OVHB\[14\].V/CLK A[15] vssd1 vssd1 vccd1 vccd1 OVHB\[14\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_06794_ _06820_/CLK line[91] vssd1 vssd1 vccd1 vccd1 _06795_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_208_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[3\].VALID\[10\].FF OVHB\[3\].V/CLK A[17] vssd1 vssd1 vccd1 vccd1 OVHB\[3\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_08533_ _08535_/CLK line[104] vssd1 vssd1 vccd1 vccd1 _08534_/A sky130_fd_sc_hd__dfxtp_1
X_05745_ _05745_/A _05774_/Y vssd1 vssd1 vccd1 vccd1 _13865_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11443__A _13926_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08464_ _08464_/A _08469_/Y vssd1 vssd1 vccd1 vccd1 _13784_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.M\[0\].MUX\[2\]_A2 _13772_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05676_ _05700_/CLK line[92] vssd1 vssd1 vccd1 vccd1 _05677_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07415_ _07415_/CLK line[105] vssd1 vssd1 vccd1 vccd1 _07416_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_211_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08395_ _08395_/CLK line[41] vssd1 vssd1 vccd1 vccd1 _08396_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07346_ _07346_/A _07349_/Y vssd1 vssd1 vccd1 vccd1 _13786_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10209__D line[102] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07277_ _07277_/CLK _07278_/X vssd1 vssd1 vccd1 vccd1 _07275_/CLK sky130_fd_sc_hd__dlclkp_1
X_09016_ _09016_/A _09029_/Y vssd1 vssd1 vccd1 vccd1 _13776_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_128_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08902__D line[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06228_ _13903_/X wr vssd1 vssd1 vccd1 vccd1 _06228_/X sky130_fd_sc_hd__and2_1
XFILLER_151_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06159_ _13903_/X vssd1 vssd1 vccd1 vccd1 _06159_/Y sky130_fd_sc_hd__inv_2
XANTENNA__07518__D line[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11618__A _13926_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09918_ _09918_/A _09939_/Y vssd1 vssd1 vccd1 vccd1 _13838_/Z sky130_fd_sc_hd__ebufn_2
X_09849_ _09865_/CLK line[65] vssd1 vssd1 vccd1 vccd1 _09850_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_58_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12860_ _12860_/A _12879_/Y vssd1 vssd1 vccd1 vccd1 _13700_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_170_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07253__D line[45] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11811_ _11825_/CLK line[66] vssd1 vssd1 vccd1 vccd1 _11812_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12791_ _12805_/CLK line[2] vssd1 vssd1 vccd1 vccd1 _12792_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_14_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11742_ _11742_/A _11759_/Y vssd1 vssd1 vccd1 vccd1 _13702_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11673_ _11685_/CLK line[3] vssd1 vssd1 vccd1 vccd1 _11674_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13412_ _13412_/A _13439_/Y vssd1 vssd1 vccd1 vccd1 _13692_/Z sky130_fd_sc_hd__ebufn_2
X_10624_ _10624_/A _10639_/Y vssd1 vssd1 vccd1 vccd1 _13704_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_OVHB\[13\].VALID\[2\].FF_D A[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05501__D line[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13343_ _13365_/CLK line[13] vssd1 vssd1 vccd1 vccd1 _13344_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10119__D line[75] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10555_ _10565_/CLK line[4] vssd1 vssd1 vccd1 vccd1 _10556_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_185_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07278__A _13910_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13274_ _13274_/A _13299_/Y vssd1 vssd1 vccd1 vccd1 _13834_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_154_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10486_ _10486_/A _10499_/Y vssd1 vssd1 vccd1 vccd1 _13846_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_142_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12225_ _12245_/CLK line[14] vssd1 vssd1 vccd1 vccd1 _12226_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12334__D line[49] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07428__D line[125] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12156_ _12156_/A _12179_/Y vssd1 vssd1 vccd1 vccd1 _13836_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_96_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11107_ _11125_/CLK line[15] vssd1 vssd1 vccd1 vccd1 _11108_/A sky130_fd_sc_hd__dfxtp_1
X_12087_ _12105_/CLK line[79] vssd1 vssd1 vccd1 vccd1 _12088_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09643__D line[99] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11038_ _11038_/A _11059_/Y vssd1 vssd1 vccd1 vccd1 _13838_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[17\].VALID\[10\].FF OVHB\[17\].V/CLK A[17] vssd1 vssd1 vccd1 vccd1 OVHB\[17\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_37_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12989_ _13015_/CLK line[107] vssd1 vssd1 vccd1 vccd1 _12990_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[28\].VALID\[13\].TOBUF OVHB\[28\].VALID\[13\].FF/Q OVHB\[28\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04916_/B2 sky130_fd_sc_hd__ebufn_2
X_05530_ _05560_/CLK line[16] vssd1 vssd1 vccd1 vccd1 _05531_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_32_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_OVHB\[4\].VALID\[9\].FF_D A[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05461_ _05461_/A _05494_/Y vssd1 vssd1 vccd1 vccd1 _13861_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12509__D line[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07200_ _07200_/A _07209_/Y vssd1 vssd1 vccd1 vccd1 _13640_/Z sky130_fd_sc_hd__ebufn_2
X_08180_ _08180_/A _08189_/Y vssd1 vssd1 vccd1 vccd1 _13780_/Z sky130_fd_sc_hd__ebufn_2
X_05392_ _05420_/CLK line[90] vssd1 vssd1 vccd1 vccd1 _05393_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_192_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07131_ _07135_/CLK line[103] vssd1 vssd1 vccd1 vccd1 _07132_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_158_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09818__D line[51] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07062_ _07062_/A _07069_/Y vssd1 vssd1 vccd1 vccd1 _13782_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_161_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06013_ _06015_/CLK line[104] vssd1 vssd1 vccd1 vccd1 _06014_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_145_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13918__A A[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06242__D line[95] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[27\].VALID\[1\].TOBUF OVHB\[27\].VALID\[1\].FF/Q OVHB\[27\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04926_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_99_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07964_ _07964_/A _07979_/Y vssd1 vssd1 vccd1 vccd1 _13844_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[21\].VALID\[12\].TOBUF OVHB\[21\].VALID\[12\].FF/Q OVHB\[21\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04929_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_114_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09703_ _09725_/CLK line[13] vssd1 vssd1 vccd1 vccd1 _09704_/A sky130_fd_sc_hd__dfxtp_1
X_06915_ _06925_/CLK line[4] vssd1 vssd1 vccd1 vccd1 _06916_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10699__D line[70] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07895_ _07905_/CLK line[68] vssd1 vssd1 vccd1 vccd1 _07896_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13075__D line[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09634_ _09634_/A _09659_/Y vssd1 vssd1 vccd1 vccd1 _13834_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08169__D line[65] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06846_ _06846_/A _06859_/Y vssd1 vssd1 vccd1 vccd1 _13846_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_55_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09565_ _09585_/CLK line[78] vssd1 vssd1 vccd1 vccd1 _09566_/A sky130_fd_sc_hd__dfxtp_1
X_06777_ _06785_/CLK line[69] vssd1 vssd1 vccd1 vccd1 _06778_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[7\].VALID\[1\].FF OVHB\[7\].V/CLK A[8] vssd1 vssd1 vccd1 vccd1 OVHB\[7\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_82_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08516_ _08516_/A _08539_/Y vssd1 vssd1 vccd1 vccd1 _13836_/Z sky130_fd_sc_hd__ebufn_2
XPHY_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05728_ _05728_/A _05739_/Y vssd1 vssd1 vccd1 vccd1 _13848_/Z sky130_fd_sc_hd__ebufn_2
XPHY_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09496_ _09496_/A _09519_/Y vssd1 vssd1 vccd1 vccd1 _13696_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[26\].VALID\[2\].FF_D A[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08447_ _08465_/CLK line[79] vssd1 vssd1 vccd1 vccd1 _08448_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05659_ _05665_/CLK line[70] vssd1 vssd1 vccd1 vccd1 _05660_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_169_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11323__D line[99] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06417__D line[47] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08378_ _08378_/A _08399_/Y vssd1 vssd1 vccd1 vccd1 _13698_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_139_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07329_ _07345_/CLK line[65] vssd1 vssd1 vccd1 vccd1 _07330_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_99_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08632__D line[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10340_ _10340_/A _10359_/Y vssd1 vssd1 vccd1 vccd1 _13700_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_191_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[19\].VALID\[6\].FF_D A[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10271_ _10285_/CLK line[2] vssd1 vssd1 vccd1 vccd1 _10272_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_2_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12010_ _12010_/A _12039_/Y vssd1 vssd1 vccd1 vccd1 _13690_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_2_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05991__D line[108] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13961_ A_h[0] vssd1 vssd1 vccd1 vccd1 _13971_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_93_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[19\].VALID\[7\].TOBUF OVHB\[19\].VALID\[7\].FF/Q OVHB\[19\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/A2 sky130_fd_sc_hd__ebufn_2
XFILLER_101_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12912_ _12912_/CLK _12913_/X vssd1 vssd1 vccd1 vccd1 _12910_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_19_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13892_ _13892_/CLK _13893_/X vssd1 vssd1 vccd1 vccd1 _13890_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_74_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12843_ _13937_/X wr vssd1 vssd1 vccd1 vccd1 _12843_/X sky130_fd_sc_hd__and2_1
XANTENNA__12179__A _13934_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13713__D line[40] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[18\].CLKBUF\[1\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08807__D line[101] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12774_ _13936_/X vssd1 vssd1 vccd1 vccd1 _12774_/Y sky130_fd_sc_hd__inv_2
XPHY_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11725_ _11755_/CLK line[32] vssd1 vssd1 vccd1 vccd1 _11726_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11656_ _11656_/A _11689_/Y vssd1 vssd1 vccd1 vccd1 _13616_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05231__D line[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[7\].INV _13982_/X vssd1 vssd1 vccd1 vccd1 OVHB\[7\].INV/Y sky130_fd_sc_hd__inv_2
XOVHB\[5\].VALID\[3\].FF OVHB\[5\].V/CLK A[10] vssd1 vssd1 vccd1 vccd1 OVHB\[5\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_10607_ _10635_/CLK line[42] vssd1 vssd1 vccd1 vccd1 _10608_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11587_ _11615_/CLK line[106] vssd1 vssd1 vccd1 vccd1 _11588_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_10_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13326_ _13330_/CLK line[119] vssd1 vssd1 vccd1 vccd1 _13327_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08542__D line[122] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10538_ _10538_/A _10569_/Y vssd1 vssd1 vccd1 vccd1 _13618_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_155_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12064__D line[54] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13257_ _13257_/A _13264_/Y vssd1 vssd1 vccd1 vccd1 _13817_/Z sky130_fd_sc_hd__ebufn_2
X_10469_ _10495_/CLK line[107] vssd1 vssd1 vccd1 vccd1 _10470_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[27\].V OVHB\[27\].V/CLK TIE/HI rst_n vssd1 vssd1 vccd1 vccd1 OVHB\[27\].V/Q
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07158__D line[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12208_ _12210_/CLK line[120] vssd1 vssd1 vccd1 vccd1 _12209_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_97_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12999__D line[97] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13188_ _13190_/CLK line[56] vssd1 vssd1 vccd1 vccd1 _13189_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_96_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12139_ _12139_/A _12144_/Y vssd1 vssd1 vccd1 vccd1 _13819_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__04929__B2 _04929_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09373__D line[104] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_04961_ _04965_/CLK line[7] vssd1 vssd1 vccd1 vccd1 _04962_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_38_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10312__D line[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06700_ _06700_/A _06719_/Y vssd1 vssd1 vccd1 vccd1 _13700_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13473__A _13898_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07680_ _07680_/A _07699_/Y vssd1 vssd1 vccd1 vccd1 _13840_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05406__D line[82] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06631_ _06645_/CLK line[2] vssd1 vssd1 vccd1 vccd1 _06632_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13623__D line[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09350_ _09350_/A _09379_/Y vssd1 vssd1 vccd1 vccd1 _13830_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08717__D line[74] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05703__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06562_ _06562_/A _06579_/Y vssd1 vssd1 vccd1 vccd1 _13842_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[0\].VALID\[3\].TOBUF OVHB\[0\].VALID\[3\].FF/Q OVHB\[0\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04919_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_205_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07621__D line[71] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08301_ _08325_/CLK line[12] vssd1 vssd1 vccd1 vccd1 _08302_/A sky130_fd_sc_hd__dfxtp_1
X_05513_ _05525_/CLK line[3] vssd1 vssd1 vccd1 vccd1 _05514_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12239__D line[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09281_ _09305_/CLK line[76] vssd1 vssd1 vccd1 vccd1 _09282_/A sky130_fd_sc_hd__dfxtp_1
X_06493_ _06505_/CLK line[67] vssd1 vssd1 vccd1 vccd1 _06494_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[25\].VALID\[6\].TOBUF OVHB\[25\].VALID\[6\].FF/Q OVHB\[25\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04923_/A2 sky130_fd_sc_hd__ebufn_2
X_08232_ _08232_/A _08259_/Y vssd1 vssd1 vccd1 vccd1 _13832_/Z sky130_fd_sc_hd__ebufn_2
X_05444_ _05444_/A _05459_/Y vssd1 vssd1 vccd1 vccd1 _13844_/Z sky130_fd_sc_hd__ebufn_2
X_08163_ _08185_/CLK line[77] vssd1 vssd1 vccd1 vccd1 _08164_/A sky130_fd_sc_hd__dfxtp_1
X_05375_ _05385_/CLK line[68] vssd1 vssd1 vccd1 vccd1 _05376_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_109_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09548__D line[56] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07114_ _07114_/A _07139_/Y vssd1 vssd1 vccd1 vccd1 _13834_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__04980__D line[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08094_ _08094_/A _08119_/Y vssd1 vssd1 vccd1 vccd1 _13694_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13648__A _13899_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07045_ _07065_/CLK line[78] vssd1 vssd1 vccd1 vccd1 _07046_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[18\].V OVHB\[18\].V/CLK TIE/HI rst_n vssd1 vssd1 vccd1 vccd1 OVHB\[18\].V/Q
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XOVHB\[3\].VALID\[5\].FF OVHB\[3\].V/CLK A[12] vssd1 vssd1 vccd1 vccd1 OVHB\[3\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_08996_ _08996_/A _09029_/Y vssd1 vssd1 vccd1 vccd1 _13756_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_125_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09283__D line[77] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07947_ _07975_/CLK line[106] vssd1 vssd1 vccd1 vccd1 _07948_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10222__D line[122] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07878_ _07878_/A _07909_/Y vssd1 vssd1 vccd1 vccd1 _13758_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_28_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09617_ _09617_/A _09624_/Y vssd1 vssd1 vccd1 vccd1 _13817_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_18_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06829_ _06855_/CLK line[107] vssd1 vssd1 vccd1 vccd1 _06830_/A sky130_fd_sc_hd__dfxtp_1
X_09548_ _09550_/CLK line[56] vssd1 vssd1 vccd1 vccd1 _09549_/A sky130_fd_sc_hd__dfxtp_1
XPHY_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07531__D line[44] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12149__D line[107] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09479_ _09479_/A _09484_/Y vssd1 vssd1 vccd1 vccd1 _13679_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_34_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11053__D line[104] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11510_ _11510_/CLK line[57] vssd1 vssd1 vccd1 vccd1 _11511_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_184_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06147__D line[37] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12490_ _12490_/CLK line[121] vssd1 vssd1 vccd1 vccd1 _12491_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11988__D line[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11441_ _11441_/A _11444_/Y vssd1 vssd1 vccd1 vccd1 _13681_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_156_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09458__D line[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11372_ _11372_/CLK _11373_/X vssd1 vssd1 vccd1 vccd1 _11370_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_50_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13111_ _13111_/A _13124_/Y vssd1 vssd1 vccd1 vccd1 _13671_/Z sky130_fd_sc_hd__ebufn_2
X_10323_ _13923_/X wr vssd1 vssd1 vccd1 vccd1 _10323_/X sky130_fd_sc_hd__and2_1
XFILLER_166_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13042_ _13050_/CLK line[117] vssd1 vssd1 vccd1 vccd1 _13043_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[31\].VALID\[5\].TOBUF OVHB\[31\].VALID\[5\].FF/Q OVHB\[31\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04927_/B2 sky130_fd_sc_hd__ebufn_2
X_10254_ _13922_/X vssd1 vssd1 vccd1 vccd1 _10254_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12612__D line[63] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10185_ _10215_/CLK line[96] vssd1 vssd1 vccd1 vccd1 _10186_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_78_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07706__D line[124] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[0\].VALID\[10\].FF_D A[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06610__D line[121] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11228__D line[56] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13944_ _13949_/C _13949_/A _13949_/B _13949_/D vssd1 vssd1 vccd1 vccd1 _13944_/X
+ sky130_fd_sc_hd__and4bb_4
XANTENNA__09921__D line[98] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[1\].VALID\[7\].FF OVHB\[1\].V/CLK A[14] vssd1 vssd1 vccd1 vccd1 OVHB\[1\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_13875_ _13875_/A _13894_/Y vssd1 vssd1 vccd1 vccd1 _13875_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_201_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12826_ _12840_/CLK line[18] vssd1 vssd1 vccd1 vccd1 _12827_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_62_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12757_ _12757_/A _12774_/Y vssd1 vssd1 vccd1 vccd1 _13877_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_91_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11708_ _11720_/CLK line[19] vssd1 vssd1 vccd1 vccd1 _11709_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06057__D line[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12688_ _12700_/CLK line[83] vssd1 vssd1 vccd1 vccd1 _12689_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11639_ _11639_/A _11654_/Y vssd1 vssd1 vccd1 vccd1 _13879_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_30_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_DATA\[16\].CLKBUF\[3\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05896__D line[50] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05160_ _05160_/A _05179_/Y vssd1 vssd1 vccd1 vccd1 _13840_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08272__D line[127] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13309_ _13309_/A _13334_/Y vssd1 vssd1 vccd1 vccd1 _13869_/Z sky130_fd_sc_hd__ebufn_2
X_05091_ _05105_/CLK line[66] vssd1 vssd1 vccd1 vccd1 _05092_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_170_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08850_ _08850_/CLK line[121] vssd1 vssd1 vccd1 vccd1 _08851_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[8\].VALID\[10\].FF OVHB\[8\].V/CLK A[17] vssd1 vssd1 vccd1 vccd1 OVHB\[8\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_07801_ _07801_/A _07804_/Y vssd1 vssd1 vccd1 vccd1 _13681_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06520__D line[94] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08781_ _08781_/A _08784_/Y vssd1 vssd1 vccd1 vccd1 _13821_/Z sky130_fd_sc_hd__ebufn_2
X_05993_ _06015_/CLK line[109] vssd1 vssd1 vccd1 vccd1 _05994_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11138__D line[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MUX.M\[1\].MUX\[4\]_A2 _13762_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07732_ _07732_/CLK _07733_/X vssd1 vssd1 vccd1 vccd1 _07730_/CLK sky130_fd_sc_hd__dlclkp_1
X_04944_ _04944_/A _04969_/Y vssd1 vssd1 vccd1 vccd1 _13624_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05136__D line[87] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[9\].CLKBUF\[3\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10977__D line[69] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07663_ _13911_/X wr vssd1 vssd1 vccd1 vccd1 _07663_/X sky130_fd_sc_hd__and2_1
XOVHB\[18\].VALID\[11\].TOBUF OVHB\[18\].VALID\[11\].FF/Q OVHB\[18\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04915_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__13353__D line[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09402_ _09410_/CLK line[117] vssd1 vssd1 vccd1 vccd1 _09403_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_92_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06614_ _13904_/X vssd1 vssd1 vccd1 vccd1 _06614_/Y sky130_fd_sc_hd__inv_2
XANTENNA_OVHB\[22\].VALID\[5\].FF_D A[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08447__D line[79] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07594_ _13911_/X vssd1 vssd1 vccd1 vccd1 _07594_/Y sky130_fd_sc_hd__inv_2
XFILLER_197_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09333_ _09333_/A _09344_/Y vssd1 vssd1 vccd1 vccd1 _13813_/Z sky130_fd_sc_hd__ebufn_2
X_06545_ _06575_/CLK line[96] vssd1 vssd1 vccd1 vccd1 _06546_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_178_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09264_ _09270_/CLK line[54] vssd1 vssd1 vccd1 vccd1 _09265_/A sky130_fd_sc_hd__dfxtp_1
X_06476_ _06476_/A _06509_/Y vssd1 vssd1 vccd1 vccd1 _13756_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_139_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08215_ _08215_/A _08224_/Y vssd1 vssd1 vccd1 vccd1 _13815_/Z sky130_fd_sc_hd__ebufn_2
X_05427_ _05455_/CLK line[106] vssd1 vssd1 vccd1 vccd1 _05428_/A sky130_fd_sc_hd__dfxtp_1
X_09195_ _09195_/A _09204_/Y vssd1 vssd1 vccd1 vccd1 _13675_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[15\].VALID\[9\].FF_D A[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11601__D line[98] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08146_ _08150_/CLK line[55] vssd1 vssd1 vccd1 vccd1 _08147_/A sky130_fd_sc_hd__dfxtp_1
X_05358_ _05358_/A _05389_/Y vssd1 vssd1 vccd1 vccd1 _13758_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_4_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08077_ _08077_/A _08084_/Y vssd1 vssd1 vccd1 vccd1 _13677_/Z sky130_fd_sc_hd__ebufn_2
X_05289_ _05315_/CLK line[43] vssd1 vssd1 vccd1 vccd1 _05290_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08910__D line[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07028_ _07030_/CLK line[56] vssd1 vssd1 vccd1 vccd1 _07029_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_161_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13528__D line[83] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XOVHB\[11\].VALID\[10\].TOBUF OVHB\[11\].VALID\[10\].FF/Q OVHB\[11\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04932_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_0_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[28\].VALID\[2\].FF OVHB\[28\].V/CLK A[9] vssd1 vssd1 vccd1 vccd1 OVHB\[28\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_48_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08979_ _08979_/A _08994_/Y vssd1 vssd1 vccd1 vccd1 _13739_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_88_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XOVHB\[6\].CGAND _13937_/X wr vssd1 vssd1 vccd1 vccd1 OVHB\[6\].CGAND/X sky130_fd_sc_hd__and2_4
X_11990_ _12000_/CLK line[20] vssd1 vssd1 vccd1 vccd1 _11991_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05046__D line[60] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10887__D line[42] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10941_ _10941_/A _10954_/Y vssd1 vssd1 vccd1 vccd1 _13741_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_204_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13660_ _13680_/CLK line[30] vssd1 vssd1 vccd1 vccd1 _13661_/A sky130_fd_sc_hd__dfxtp_1
X_10872_ _10880_/CLK line[21] vssd1 vssd1 vccd1 vccd1 _10873_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07261__D line[34] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12611_ _12611_/A _12634_/Y vssd1 vssd1 vccd1 vccd1 _13731_/Z sky130_fd_sc_hd__ebufn_2
XPHY_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13591_ _13591_/A _13614_/Y vssd1 vssd1 vccd1 vccd1 _13871_/Z sky130_fd_sc_hd__ebufn_2
XPHY_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12542_ _12560_/CLK line[31] vssd1 vssd1 vccd1 vccd1 _12543_/A sky130_fd_sc_hd__dfxtp_1
XPHY_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XOVHB\[7\].VALID\[3\].TOBUF OVHB\[7\].VALID\[3\].FF/Q OVHB\[7\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04919_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_157_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12473_ _12473_/A _12494_/Y vssd1 vssd1 vccd1 vccd1 _13873_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[5\].VALID\[14\].FF_D A[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09188__D line[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11424_ _11440_/CLK line[17] vssd1 vssd1 vccd1 vccd1 _11425_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_172_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_OVHB\[3\].VALID\[0\].FF_D A[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10127__D line[79] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11355_ _11355_/A _11374_/Y vssd1 vssd1 vccd1 vccd1 _13875_/Z sky130_fd_sc_hd__ebufn_2
X_10306_ _10320_/CLK line[18] vssd1 vssd1 vccd1 vccd1 _10307_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08820__D line[112] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11286_ _11300_/CLK line[82] vssd1 vssd1 vccd1 vccd1 _11287_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12342__D line[53] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13025_ _13025_/A _13054_/Y vssd1 vssd1 vccd1 vccd1 _13865_/Z sky130_fd_sc_hd__ebufn_2
X_10237_ _10237_/A _10254_/Y vssd1 vssd1 vccd1 vccd1 _13877_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07436__D line[114] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10168_ _10180_/CLK line[83] vssd1 vssd1 vccd1 vccd1 _10169_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07733__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10099_ _10099_/A _10114_/Y vssd1 vssd1 vccd1 vccd1 _13739_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09651__D line[103] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13927_ _13927_/A _13927_/B _13927_/C _13927_/D vssd1 vssd1 vccd1 vccd1 _13927_/X
+ sky130_fd_sc_hd__and4_4
XFILLER_35_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13858_ _13899_/X wr vssd1 vssd1 vccd1 vccd1 _13858_/X sky130_fd_sc_hd__and2_1
XOVHB\[26\].VALID\[4\].FF OVHB\[26\].V/CLK A[11] vssd1 vssd1 vccd1 vccd1 OVHB\[26\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_34_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12809_ _13937_/X vssd1 vssd1 vccd1 vccd1 _12809_/Y sky130_fd_sc_hd__inv_2
X_13789_ _13899_/X vssd1 vssd1 vccd1 vccd1 _13789_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[28\].VALID\[9\].FF_D A[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06330_ _06330_/CLK line[121] vssd1 vssd1 vccd1 vccd1 _06331_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_187_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12517__D line[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06261_ _06261_/A _06264_/Y vssd1 vssd1 vccd1 vccd1 _13821_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[29\].CLKBUF\[1\] clk vssd1 vssd1 vccd1 vccd1 _10882_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_30_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XOVHB\[31\].VALID\[10\].TOBUF OVHB\[31\].VALID\[10\].FF/Q OVHB\[31\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04932_/B2 sky130_fd_sc_hd__ebufn_2
X_08000_ _08010_/CLK line[116] vssd1 vssd1 vccd1 vccd1 _08001_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[2\].CGAND_A _13933_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05212_ _05212_/CLK _05213_/X vssd1 vssd1 vccd1 vccd1 _05210_/CLK sky130_fd_sc_hd__dlclkp_1
X_06192_ _06192_/CLK _06193_/X vssd1 vssd1 vccd1 vccd1 _06190_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_144_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XDATA\[19\].CLKBUF\[7\] clk vssd1 vssd1 vccd1 vccd1 _08012_/CLK sky130_fd_sc_hd__clkbuf_4
X_05143_ _13931_/Y wr vssd1 vssd1 vccd1 vccd1 _05143_/X sky130_fd_sc_hd__and2_1
XFILLER_7_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07908__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09826__D line[55] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09951_ _09951_/A _09974_/Y vssd1 vssd1 vccd1 vccd1 _13871_/Z sky130_fd_sc_hd__ebufn_2
X_05074_ _13931_/Y vssd1 vssd1 vccd1 vccd1 _05074_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08902_ _08920_/CLK line[31] vssd1 vssd1 vccd1 vccd1 _08903_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[14\].CLKBUF\[5\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12252__D line[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09882_ _09900_/CLK line[95] vssd1 vssd1 vccd1 vccd1 _09883_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_85_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08833_ _08833_/A _08854_/Y vssd1 vssd1 vccd1 vccd1 _13873_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06250__D line[84] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08764_ _08780_/CLK line[81] vssd1 vssd1 vccd1 vccd1 _08765_/A sky130_fd_sc_hd__dfxtp_1
X_05976_ _05980_/CLK line[87] vssd1 vssd1 vccd1 vccd1 _05977_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_73_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09561__D line[76] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[7\].VALID\[10\].FF_D A[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07715_ _07715_/A _07734_/Y vssd1 vssd1 vccd1 vccd1 _13875_/Z sky130_fd_sc_hd__ebufn_2
X_04927_ A_h[10] _04927_/B2 A_h[10] _04927_/B2 vssd1 vssd1 vccd1 vccd1 _04928_/D sky130_fd_sc_hd__a2bb2oi_2
X_08695_ _08695_/A _08714_/Y vssd1 vssd1 vccd1 vccd1 _13735_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13083__D line[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MUX.M\[0\].MUX\[5\]_A0 _13638_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10500__D line[112] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08177__D line[69] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07646_ _07660_/CLK line[82] vssd1 vssd1 vccd1 vccd1 _07647_/A sky130_fd_sc_hd__dfxtp_1
X_07577_ _07577_/A _07594_/Y vssd1 vssd1 vccd1 vccd1 _13737_/Z sky130_fd_sc_hd__ebufn_2
X_09316_ _09340_/CLK line[92] vssd1 vssd1 vccd1 vccd1 _09317_/A sky130_fd_sc_hd__dfxtp_1
X_06528_ _06540_/CLK line[83] vssd1 vssd1 vccd1 vccd1 _06529_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[7\].CLKBUF\[5\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09247_ _09247_/A _09274_/Y vssd1 vssd1 vccd1 vccd1 _13727_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12427__D line[106] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06459_ _06459_/A _06474_/Y vssd1 vssd1 vccd1 vccd1 _13739_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__04926__A1_N A_h[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11331__D line[103] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[24\].VALID\[6\].FF OVHB\[24\].V/CLK A[13] vssd1 vssd1 vccd1 vccd1 OVHB\[24\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06425__D line[36] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09178_ _09200_/CLK line[29] vssd1 vssd1 vccd1 vccd1 _09179_/A sky130_fd_sc_hd__dfxtp_1
X_08129_ _08129_/A _08154_/Y vssd1 vssd1 vccd1 vccd1 _13729_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_181_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09736__D line[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08640__D line[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11140_ _11160_/CLK line[30] vssd1 vssd1 vccd1 vccd1 _11141_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13258__D line[88] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[9\].VALID\[4\].FF_D A[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11071_ _11071_/A _11094_/Y vssd1 vssd1 vccd1 vccd1 _13871_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_0_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XDATA\[18\].CLKBUF\[4\] clk vssd1 vssd1 vccd1 vccd1 _07627_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_103_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10022_ _10040_/CLK line[31] vssd1 vssd1 vccd1 vccd1 _10023_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_49_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06160__D line[48] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[5\].VALID\[8\].TOBUF OVHB\[5\].VALID\[8\].FF/Q OVHB\[5\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04931_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_56_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05354__A _13900_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11973_ _11973_/A _12004_/Y vssd1 vssd1 vccd1 vccd1 _13653_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11506__D line[55] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13712_ _13712_/A _13719_/Y vssd1 vssd1 vccd1 vccd1 _13712_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08087__D line[42] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10924_ _10950_/CLK line[59] vssd1 vssd1 vccd1 vccd1 _10925_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05073__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10855_ _10855_/A _10884_/Y vssd1 vssd1 vccd1 vccd1 _13655_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_31_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13643_ _13645_/CLK line[8] vssd1 vssd1 vccd1 vccd1 _13644_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_71_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13574_ _13574_/A _13579_/Y vssd1 vssd1 vccd1 vccd1 _13854_/Z sky130_fd_sc_hd__ebufn_2
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08815__D line[105] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10786_ _10810_/CLK line[124] vssd1 vssd1 vccd1 vccd1 _10787_/A sky130_fd_sc_hd__dfxtp_1
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12525_ _12525_/CLK line[9] vssd1 vssd1 vccd1 vccd1 _12526_/A sky130_fd_sc_hd__dfxtp_1
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11241__D line[76] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06335__D line[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12456_ _12456_/A _12459_/Y vssd1 vssd1 vccd1 vccd1 _13856_/Z sky130_fd_sc_hd__ebufn_2
X_11407_ _11407_/CLK _11408_/X vssd1 vssd1 vccd1 vccd1 _11405_/CLK sky130_fd_sc_hd__dlclkp_1
X_12387_ _12387_/CLK _12388_/X vssd1 vssd1 vccd1 vccd1 _12385_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_207_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05529__A _13901_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08550__D line[126] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11338_ _13933_/X wr vssd1 vssd1 vccd1 vccd1 _11338_/X sky130_fd_sc_hd__and2_1
XFILLER_140_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13168__D line[61] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05248__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11269_ _13933_/X vssd1 vssd1 vccd1 vccd1 _11269_/Y sky130_fd_sc_hd__inv_2
XANTENNA__07166__D line[119] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[22\].VALID\[8\].FF OVHB\[22\].V/CLK A[15] vssd1 vssd1 vccd1 vccd1 OVHB\[22\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_13008_ _13008_/A _13019_/Y vssd1 vssd1 vccd1 vccd1 _13848_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[30\].V_RESET_B rst_n vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[30\].VALID\[13\].FF OVHB\[30\].V/CLK A[20] vssd1 vssd1 vccd1 vccd1 OVHB\[30\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_05830_ _05840_/CLK line[20] vssd1 vssd1 vccd1 vccd1 _05831_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XDATA\[17\].CLKBUF\[1\] clk vssd1 vssd1 vccd1 vccd1 _07242_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_82_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05761_ _05761_/A _05774_/Y vssd1 vssd1 vccd1 vccd1 _13881_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_48_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11416__D line[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07500_ _07520_/CLK line[30] vssd1 vssd1 vccd1 vccd1 _07501_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10320__D line[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08480_ _08500_/CLK line[94] vssd1 vssd1 vccd1 vccd1 _08481_/A sky130_fd_sc_hd__dfxtp_1
X_05692_ _05700_/CLK line[85] vssd1 vssd1 vccd1 vccd1 _05693_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05414__D line[86] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07431_ _07431_/A _07454_/Y vssd1 vssd1 vccd1 vccd1 _13871_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13631__D line[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XOVHB\[12\].VALID\[3\].TOBUF OVHB\[12\].VALID\[3\].FF/Q OVHB\[12\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04919_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__08725__D line[78] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07362_ _07380_/CLK line[95] vssd1 vssd1 vccd1 vccd1 _07363_/A sky130_fd_sc_hd__dfxtp_1
X_09101_ _09101_/A _09134_/Y vssd1 vssd1 vccd1 vccd1 _13861_/Z sky130_fd_sc_hd__ebufn_2
X_06313_ _06313_/A _06334_/Y vssd1 vssd1 vccd1 vccd1 _13873_/Z sky130_fd_sc_hd__ebufn_2
X_07293_ _07293_/A _07314_/Y vssd1 vssd1 vccd1 vccd1 _13733_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_30_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09032_ _09060_/CLK line[90] vssd1 vssd1 vccd1 vccd1 _09033_/A sky130_fd_sc_hd__dfxtp_1
X_06244_ _06260_/CLK line[81] vssd1 vssd1 vccd1 vccd1 _06245_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_190_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06823__A _13905_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10990__D line[80] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06175_ _06175_/A _06194_/Y vssd1 vssd1 vccd1 vccd1 _13735_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_117_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05126_ _05140_/CLK line[82] vssd1 vssd1 vccd1 vccd1 _05127_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_171_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05057_ _05057_/A _05074_/Y vssd1 vssd1 vccd1 vccd1 _13737_/Z sky130_fd_sc_hd__ebufn_2
X_09934_ _09934_/A _09939_/Y vssd1 vssd1 vccd1 vccd1 _13854_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07076__D line[92] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09865_ _09865_/CLK line[73] vssd1 vssd1 vccd1 vccd1 _09866_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_58_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13806__D line[82] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08816_ _08816_/A _08819_/Y vssd1 vssd1 vccd1 vccd1 _13856_/Z sky130_fd_sc_hd__ebufn_2
X_09796_ _09796_/A _09799_/Y vssd1 vssd1 vccd1 vccd1 _13716_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_133_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09291__D line[66] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08747_ _08747_/CLK _08748_/X vssd1 vssd1 vccd1 vccd1 _08745_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA_DATA\[12\].CLKBUF\[7\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05959_ _05959_/A _05984_/Y vssd1 vssd1 vccd1 vccd1 _13799_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10230__D line[126] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08678_ _13914_/X wr vssd1 vssd1 vccd1 vccd1 _08678_/X sky130_fd_sc_hd__and2_1
XANTENNA__05324__D line[59] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_DECH.DEC0.AND2_A_N A_h[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07629_ _13911_/X vssd1 vssd1 vccd1 vccd1 _07629_/Y sky130_fd_sc_hd__inv_2
XPHY_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10640_ _10670_/CLK line[48] vssd1 vssd1 vccd1 vccd1 _10641_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12157__D line[111] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10571_ _10571_/A _10604_/Y vssd1 vssd1 vccd1 vccd1 _13651_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_42_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12310_ _12310_/A _12319_/Y vssd1 vssd1 vccd1 vccd1 _13710_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_166_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06155__D line[41] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13290_ _13290_/A _13299_/Y vssd1 vssd1 vccd1 vccd1 _13850_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11996__D line[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12241_ _12245_/CLK line[7] vssd1 vssd1 vccd1 vccd1 _12242_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09466__D line[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[5\].CLKBUF\[7\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12172_ _12172_/A _12179_/Y vssd1 vssd1 vccd1 vccd1 _13852_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_107_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11123_ _11125_/CLK line[8] vssd1 vssd1 vccd1 vccd1 _11124_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09763__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10405__D line[78] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11054_ _11054_/A _11059_/Y vssd1 vssd1 vccd1 vccd1 _13854_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[31\].VALID\[8\].FF_D A[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10005_ _10005_/CLK line[9] vssd1 vssd1 vccd1 vccd1 _10006_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12620__D line[52] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07714__D line[113] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[8\].VALID\[13\].TOBUF OVHB\[8\].VALID\[13\].FF/Q OVHB\[8\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04916_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_36_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11956_ _11956_/A _11969_/Y vssd1 vssd1 vccd1 vccd1 _13636_/Z sky130_fd_sc_hd__ebufn_2
X_10907_ _10915_/CLK line[37] vssd1 vssd1 vccd1 vccd1 _10908_/A sky130_fd_sc_hd__dfxtp_1
X_11887_ _11895_/CLK line[101] vssd1 vssd1 vccd1 vccd1 _11888_/A sky130_fd_sc_hd__dfxtp_1
X_10838_ _10838_/A _10849_/Y vssd1 vssd1 vccd1 vccd1 _13638_/Z sky130_fd_sc_hd__ebufn_2
X_13626_ _13626_/A _13649_/Y vssd1 vssd1 vccd1 vccd1 _13626_/Z sky130_fd_sc_hd__ebufn_2
X_13557_ _13575_/CLK line[111] vssd1 vssd1 vccd1 vccd1 _13558_/A sky130_fd_sc_hd__dfxtp_1
X_10769_ _10775_/CLK line[102] vssd1 vssd1 vccd1 vccd1 _10770_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09938__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06065__D line[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12508_ _12508_/A _12529_/Y vssd1 vssd1 vccd1 vccd1 _13628_/Z sky130_fd_sc_hd__ebufn_2
X_13488_ _13488_/A _13509_/Y vssd1 vssd1 vccd1 vccd1 _13768_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_145_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12439_ _12455_/CLK line[97] vssd1 vssd1 vccd1 vccd1 _12440_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08280__D line[116] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MUX.M\[2\].MUX\[6\]_A2 _13815_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[1\].VALID\[12\].TOBUF OVHB\[1\].VALID\[12\].FF/Q OVHB\[1\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04929_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_99_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07980_ _08010_/CLK line[112] vssd1 vssd1 vccd1 vccd1 _07981_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[14\].VALID\[0\].FF_D A[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06931_ _06931_/A _06964_/Y vssd1 vssd1 vccd1 vccd1 _13651_/Z sky130_fd_sc_hd__ebufn_2
XMUX.M\[1\].MUX\[0\] _13644_/Z _13714_/Z _13784_/Z _13854_/Z MUX.SEL0BUF\[1\]/X MUX.SEL1BUF\[1\]/X
+ vssd1 vssd1 vccd1 vccd1 Do[8] sky130_fd_sc_hd__mux4_1
XOVHB\[10\].VALID\[8\].TOBUF OVHB\[10\].VALID\[8\].FF/Q OVHB\[10\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04931_/B2 sky130_fd_sc_hd__ebufn_2
X_09650_ _09650_/A _09659_/Y vssd1 vssd1 vccd1 vccd1 _13850_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12530__D line[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06862_ _06890_/CLK line[122] vssd1 vssd1 vccd1 vccd1 _06863_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_83_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08601_ _08605_/CLK line[7] vssd1 vssd1 vccd1 vccd1 _08602_/A sky130_fd_sc_hd__dfxtp_1
X_05813_ _05813_/A _05844_/Y vssd1 vssd1 vccd1 vccd1 _13653_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_82_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09581_ _09585_/CLK line[71] vssd1 vssd1 vccd1 vccd1 _09582_/A sky130_fd_sc_hd__dfxtp_1
X_06793_ _06793_/A _06824_/Y vssd1 vssd1 vccd1 vccd1 _13793_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11146__D line[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[11\].CG_CLK clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11724__A _13927_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08532_ _08532_/A _08539_/Y vssd1 vssd1 vccd1 vccd1 _13852_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[12\].CG clk OVHB\[12\].CGAND/X vssd1 vssd1 vccd1 vccd1 OVHB\[12\].V/CLK sky130_fd_sc_hd__dlclkp_1
X_05744_ _05770_/CLK line[123] vssd1 vssd1 vccd1 vccd1 _05745_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_63_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11443__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10985__D line[73] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08463_ _08465_/CLK line[72] vssd1 vssd1 vccd1 vccd1 _08464_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_35_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05675_ _05675_/A _05704_/Y vssd1 vssd1 vccd1 vccd1 _13795_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13361__D line[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MUX.M\[0\].MUX\[2\]_A3 _13842_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07414_ _07414_/A _07419_/Y vssd1 vssd1 vccd1 vccd1 _13854_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_196_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08455__D line[68] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08394_ _08394_/A _08399_/Y vssd1 vssd1 vccd1 vccd1 _13714_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07345_ _07345_/CLK line[73] vssd1 vssd1 vccd1 vccd1 _07346_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_149_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07276_ _07276_/A _07279_/Y vssd1 vssd1 vccd1 vccd1 _13716_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_176_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09015_ _09025_/CLK line[68] vssd1 vssd1 vccd1 vccd1 _09016_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_164_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06227_ _06227_/CLK _06228_/X vssd1 vssd1 vccd1 vccd1 _06225_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_191_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12705__D line[96] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_OVHB\[5\].VALID\[7\].FF_D A[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06703__D line[35] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08190__D line[80] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06158_ _13903_/X wr vssd1 vssd1 vccd1 vccd1 _06158_/X sky130_fd_sc_hd__and2_1
XFILLER_144_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05109_ _13931_/Y vssd1 vssd1 vccd1 vccd1 _05109_/Y sky130_fd_sc_hd__inv_2
X_06089_ _13903_/X vssd1 vssd1 vccd1 vccd1 _06089_/Y sky130_fd_sc_hd__inv_2
XANTENNA__07384__A _13910_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11618__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09917_ _09935_/CLK line[111] vssd1 vssd1 vccd1 vccd1 _09918_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13536__D line[87] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[26\].CLKBUF\[1\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09848_ _09848_/A _09869_/Y vssd1 vssd1 vccd1 vccd1 _13768_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_100_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09779_ _09795_/CLK line[33] vssd1 vssd1 vccd1 vccd1 _09780_/A sky130_fd_sc_hd__dfxtp_1
X_11810_ _11810_/A _11829_/Y vssd1 vssd1 vccd1 vccd1 _13770_/Z sky130_fd_sc_hd__ebufn_2
X_12790_ _12790_/A _12809_/Y vssd1 vssd1 vccd1 vccd1 _13630_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05054__D line[49] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10895__D line[46] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11741_ _11755_/CLK line[34] vssd1 vssd1 vccd1 vccd1 _11742_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13271__D line[108] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05989__D line[107] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08365__D line[32] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11672_ _11672_/A _11689_/Y vssd1 vssd1 vccd1 vccd1 _13632_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMUX.M\[0\].MUX\[2\] _13632_/Z _13702_/Z _13772_/Z _13842_/Z MUX.SEL0BUF\[0\]/X MUX.SEL1BUF\[0\]/X
+ vssd1 vssd1 vccd1 vccd1 Do[2] sky130_fd_sc_hd__mux4_1
XPHY_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[14\].VALID\[12\].FF_D A[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10623_ _10635_/CLK line[35] vssd1 vssd1 vccd1 vccd1 _10624_/A sky130_fd_sc_hd__dfxtp_1
X_13411_ _13435_/CLK line[44] vssd1 vssd1 vccd1 vccd1 _13412_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13342_ _13342_/A _13369_/Y vssd1 vssd1 vccd1 vccd1 _13622_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07559__A _13911_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[19\].VALID\[3\].TOBUF OVHB\[19\].VALID\[3\].FF/Q OVHB\[19\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04919_/B2 sky130_fd_sc_hd__ebufn_2
X_10554_ _10554_/A _10569_/Y vssd1 vssd1 vccd1 vccd1 _13634_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_185_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07278__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13273_ _13295_/CLK line[109] vssd1 vssd1 vccd1 vccd1 _13274_/A sky130_fd_sc_hd__dfxtp_1
X_10485_ _10495_/CLK line[100] vssd1 vssd1 vccd1 vccd1 _10486_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09196__D line[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12224_ _12224_/A _12249_/Y vssd1 vssd1 vccd1 vccd1 _13624_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[27\].VALID\[0\].FF_D A[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12155_ _12175_/CLK line[110] vssd1 vssd1 vccd1 vccd1 _12156_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10135__D line[68] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05229__D line[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11106_ _11106_/A _11129_/Y vssd1 vssd1 vccd1 vccd1 _13626_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[24\].VALID\[11\].FF_D A[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12086_ _12086_/A _12109_/Y vssd1 vssd1 vccd1 vccd1 _13766_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13446__D line[60] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[24\].VALID\[14\].TOBUF OVHB\[24\].VALID\[14\].FF/Q OVHB\[24\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_49_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12350__D line[57] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11037_ _11055_/CLK line[111] vssd1 vssd1 vccd1 vccd1 _11038_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_92_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07444__D line[118] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12988_ _12988_/A _13019_/Y vssd1 vssd1 vccd1 vccd1 _13828_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_17_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11939_ _11965_/CLK line[11] vssd1 vssd1 vccd1 vccd1 _11940_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[7\].CG clk OVHB\[7\].CGAND/X vssd1 vssd1 vccd1 vccd1 OVHB\[7\].V/CLK sky130_fd_sc_hd__dlclkp_1
X_05460_ _05490_/CLK line[112] vssd1 vssd1 vccd1 vccd1 _05461_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08853__A _13914_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13609_ _13609_/A _13614_/Y vssd1 vssd1 vccd1 vccd1 _13889_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_20_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05391_ _05391_/A _05424_/Y vssd1 vssd1 vccd1 vccd1 _13791_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_186_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07130_ _07130_/A _07139_/Y vssd1 vssd1 vccd1 vccd1 _13850_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_158_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12525__D line[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07061_ _07065_/CLK line[71] vssd1 vssd1 vccd1 vccd1 _07062_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07619__D line[70] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06012_ _06012_/A _06019_/Y vssd1 vssd1 vccd1 vccd1 _13852_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[2\].V_D TIE/HI vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10045__D line[32] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[25\].VALID\[2\].TOBUF OVHB\[25\].VALID\[2\].FF/Q OVHB\[25\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04930_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.M\[1\].MUX\[7\]_A0 _13628_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07963_ _07975_/CLK line[99] vssd1 vssd1 vccd1 vccd1 _07964_/A sky130_fd_sc_hd__dfxtp_1
X_09702_ _09702_/A _09729_/Y vssd1 vssd1 vccd1 vccd1 _13622_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12260__D line[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06914_ _06914_/A _06929_/Y vssd1 vssd1 vccd1 vccd1 _13634_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[8\].CLKBUF\[5\] clk vssd1 vssd1 vccd1 vccd1 _13542_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__04978__D line[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07894_ _07894_/A _07909_/Y vssd1 vssd1 vccd1 vccd1 _13774_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07354__D line[91] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09633_ _09655_/CLK line[109] vssd1 vssd1 vccd1 vccd1 _09634_/A sky130_fd_sc_hd__dfxtp_1
X_06845_ _06855_/CLK line[100] vssd1 vssd1 vccd1 vccd1 _06846_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_83_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09564_ _09564_/A _09589_/Y vssd1 vssd1 vccd1 vccd1 _13764_/Z sky130_fd_sc_hd__ebufn_2
X_06776_ _06776_/A _06789_/Y vssd1 vssd1 vccd1 vccd1 _13776_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_130_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08515_ _08535_/CLK line[110] vssd1 vssd1 vccd1 vccd1 _08516_/A sky130_fd_sc_hd__dfxtp_1
X_05727_ _05735_/CLK line[101] vssd1 vssd1 vccd1 vccd1 _05728_/A sky130_fd_sc_hd__dfxtp_1
X_09495_ _09515_/CLK line[46] vssd1 vssd1 vccd1 vccd1 _09496_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_130_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08446_ _08446_/A _08469_/Y vssd1 vssd1 vccd1 vccd1 _13766_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08185__D line[73] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05658_ _05658_/A _05669_/Y vssd1 vssd1 vccd1 vccd1 _13778_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05602__D line[58] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08377_ _08395_/CLK line[47] vssd1 vssd1 vccd1 vccd1 _08378_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05589_ _05595_/CLK line[38] vssd1 vssd1 vccd1 vccd1 _05590_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_7_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07328_ _07328_/A _07349_/Y vssd1 vssd1 vccd1 vccd1 _13768_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_177_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07259_ _07275_/CLK line[33] vssd1 vssd1 vccd1 vccd1 _07260_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12435__D line[110] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07529__D line[43] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06433__D line[40] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10270_ _10270_/A _10289_/Y vssd1 vssd1 vccd1 vccd1 _13630_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_191_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10533__A _13923_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09744__D line[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13960_ _13960_/A _13960_/B _13960_/C _13960_/D vssd1 vssd1 vccd1 vccd1 _13960_/X
+ sky130_fd_sc_hd__and4_4
XFILLER_48_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12911_ _12911_/A _12914_/Y vssd1 vssd1 vccd1 vccd1 _13751_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[17\].VALID\[8\].TOBUF OVHB\[17\].VALID\[8\].FF/Q OVHB\[17\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04931_/B2 sky130_fd_sc_hd__ebufn_2
X_13891_ _13891_/A _13894_/Y vssd1 vssd1 vccd1 vccd1 _13891_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[21\].INV _13958_/X vssd1 vssd1 vccd1 vccd1 OVHB\[21\].INV/Y sky130_fd_sc_hd__inv_2
X_12842_ _12842_/CLK _12843_/X vssd1 vssd1 vccd1 vccd1 _12840_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_64_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XDATA\[7\].CLKBUF\[2\] clk vssd1 vssd1 vccd1 vccd1 _13157_/CLK sky130_fd_sc_hd__clkbuf_4
XPHY_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_DATA\[24\].CLKBUF\[3\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12773_ _13936_/X wr vssd1 vssd1 vccd1 vccd1 _12773_/X sky130_fd_sc_hd__and2_1
XPHY_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XOVHB\[31\].VALID\[1\].TOBUF OVHB\[31\].VALID\[1\].FF/Q OVHB\[31\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04926_/B2 sky130_fd_sc_hd__ebufn_2
XPHY_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08095__D line[46] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11724_ _13927_/X vssd1 vssd1 vccd1 vccd1 _11724_/Y sky130_fd_sc_hd__inv_2
XANTENNA__06608__D line[120] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11655_ _11685_/CLK line[0] vssd1 vssd1 vccd1 vccd1 _11656_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10708__A _13924_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09919__D line[97] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10606_ _10606_/A _10639_/Y vssd1 vssd1 vccd1 vccd1 _13686_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06193__A _13903_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11586_ _11586_/A _11619_/Y vssd1 vssd1 vccd1 vccd1 _13826_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_167_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10537_ _10565_/CLK line[10] vssd1 vssd1 vccd1 vccd1 _10538_/A sky130_fd_sc_hd__dfxtp_1
X_13325_ _13325_/A _13334_/Y vssd1 vssd1 vccd1 vccd1 _13885_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_182_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06343__D line[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10468_ _10468_/A _10499_/Y vssd1 vssd1 vccd1 vccd1 _13828_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[10\].VALID\[3\].FF_D A[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13256_ _13260_/CLK line[87] vssd1 vssd1 vccd1 vccd1 _13257_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[8\].VALID\[8\].FF OVHB\[8\].V/CLK A[15] vssd1 vssd1 vccd1 vccd1 OVHB\[8\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_12207_ _12207_/A _12214_/Y vssd1 vssd1 vccd1 vccd1 _13887_/Z sky130_fd_sc_hd__ebufn_2
X_13187_ _13187_/A _13194_/Y vssd1 vssd1 vccd1 vccd1 _13747_/Z sky130_fd_sc_hd__ebufn_2
X_10399_ _10425_/CLK line[75] vssd1 vssd1 vccd1 vccd1 _10400_/A sky130_fd_sc_hd__dfxtp_1
X_12138_ _12140_/CLK line[88] vssd1 vssd1 vccd1 vccd1 _12139_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_150_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13176__D line[50] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDATA\[27\].CLKBUF\[6\] clk vssd1 vssd1 vccd1 vccd1 _10497_/CLK sky130_fd_sc_hd__clkbuf_4
XMUX.M\[3\].MUX\[7\] _13663_/Z _13733_/Z _13803_/Z _13873_/Z MUX.SEL0BUF\[3\]/X MUX.SEL1BUF\[3\]/X
+ vssd1 vssd1 vccd1 vccd1 Do[31] sky130_fd_sc_hd__mux4_1
XANTENNA__13754__A _13899_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_04960_ _04960_/A _04969_/Y vssd1 vssd1 vccd1 vccd1 _13640_/Z sky130_fd_sc_hd__ebufn_2
X_12069_ _12069_/A _12074_/Y vssd1 vssd1 vccd1 vccd1 _13749_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_65_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13473__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06630_ _06630_/A _06649_/Y vssd1 vssd1 vccd1 vccd1 _13630_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_53_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06368__A _13904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06561_ _06575_/CLK line[98] vssd1 vssd1 vccd1 vccd1 _06562_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11424__D line[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08300_ _08300_/A _08329_/Y vssd1 vssd1 vccd1 vccd1 _13620_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_33_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05512_ _05512_/A _05529_/Y vssd1 vssd1 vccd1 vccd1 _13632_/Z sky130_fd_sc_hd__ebufn_2
X_09280_ _09280_/A _09309_/Y vssd1 vssd1 vccd1 vccd1 _13760_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06518__D line[93] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06492_ _06492_/A _06509_/Y vssd1 vssd1 vccd1 vccd1 _13772_/Z sky130_fd_sc_hd__ebufn_2
X_08231_ _08255_/CLK line[108] vssd1 vssd1 vccd1 vccd1 _08232_/A sky130_fd_sc_hd__dfxtp_1
X_05443_ _05455_/CLK line[99] vssd1 vssd1 vccd1 vccd1 _05444_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[23\].VALID\[7\].TOBUF OVHB\[23\].VALID\[7\].FF/Q OVHB\[23\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/A2 sky130_fd_sc_hd__ebufn_2
XANTENNA__08733__D line[67] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08162_ _08162_/A _08189_/Y vssd1 vssd1 vccd1 vccd1 _13762_/Z sky130_fd_sc_hd__ebufn_2
X_05374_ _05374_/A _05389_/Y vssd1 vssd1 vccd1 vccd1 _13774_/Z sky130_fd_sc_hd__ebufn_2
X_07113_ _07135_/CLK line[109] vssd1 vssd1 vccd1 vccd1 _07114_/A sky130_fd_sc_hd__dfxtp_1
X_08093_ _08115_/CLK line[45] vssd1 vssd1 vccd1 vccd1 _08094_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_109_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13929__A A[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07044_ _07044_/A _07069_/Y vssd1 vssd1 vccd1 vccd1 _13764_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13648__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08995_ _09025_/CLK line[64] vssd1 vssd1 vccd1 vccd1 _08996_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_197_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07946_ _07946_/A _07979_/Y vssd1 vssd1 vccd1 vccd1 _13826_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07084__D line[81] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07877_ _07905_/CLK line[74] vssd1 vssd1 vccd1 vccd1 _07878_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_95_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13814__D line[86] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09616_ _09620_/CLK line[87] vssd1 vssd1 vccd1 vccd1 _09617_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_44_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08908__D line[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDATA\[26\].CLKBUF\[3\] clk vssd1 vssd1 vccd1 vccd1 _10112_/CLK sky130_fd_sc_hd__clkbuf_4
X_06828_ _06828_/A _06859_/Y vssd1 vssd1 vccd1 vccd1 _13828_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_83_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06759_ _06785_/CLK line[75] vssd1 vssd1 vccd1 vccd1 _06760_/A sky130_fd_sc_hd__dfxtp_1
X_09547_ _09547_/A _09554_/Y vssd1 vssd1 vccd1 vccd1 _13747_/Z sky130_fd_sc_hd__ebufn_2
XPHY_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09589__A _13920_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09478_ _09480_/CLK line[24] vssd1 vssd1 vccd1 vccd1 _09479_/A sky130_fd_sc_hd__dfxtp_1
XPHY_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05332__D line[63] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08429_ _08429_/A _08434_/Y vssd1 vssd1 vccd1 vccd1 _13749_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11440_ _11440_/CLK line[25] vssd1 vssd1 vccd1 vccd1 _11441_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XOVHB\[2\].CGAND _13933_/X wr vssd1 vssd1 vccd1 vccd1 OVHB\[2\].CGAND/X sky130_fd_sc_hd__and2_4
XANTENNA__12165__D line[100] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11371_ _11371_/A _11374_/Y vssd1 vssd1 vccd1 vccd1 _13891_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[23\].VALID\[3\].FF_D A[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07259__D line[33] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13110_ _13120_/CLK line[20] vssd1 vssd1 vccd1 vccd1 _13111_/A sky130_fd_sc_hd__dfxtp_1
X_10322_ _10322_/CLK _10323_/X vssd1 vssd1 vccd1 vccd1 _10320_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_50_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13041_ _13041_/A _13054_/Y vssd1 vssd1 vccd1 vccd1 _13881_/Z sky130_fd_sc_hd__ebufn_2
X_10253_ _13922_/X wr vssd1 vssd1 vccd1 vccd1 _10253_/X sky130_fd_sc_hd__and2_1
XANTENNA__09474__D line[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[17\].VALID\[0\].FF OVHB\[17\].V/CLK A[7] vssd1 vssd1 vccd1 vccd1 OVHB\[17\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_10184_ _13922_/X vssd1 vssd1 vccd1 vccd1 _10184_/Y sky130_fd_sc_hd__inv_2
XANTENNA_OVHB\[16\].VALID\[7\].FF_D A[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10413__D line[67] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05507__D line[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13943_ _13949_/C _13949_/B _13949_/A _13949_/D vssd1 vssd1 vccd1 vccd1 _13943_/X
+ sky130_fd_sc_hd__and4bb_4
XANTENNA__13724__D line[59] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11094__A _13925_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13874_ _13890_/CLK line[113] vssd1 vssd1 vccd1 vccd1 _13875_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07722__D line[117] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12825_ _12825_/A _12844_/Y vssd1 vssd1 vccd1 vccd1 _13665_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_91_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12756_ _12770_/CLK line[114] vssd1 vssd1 vccd1 vccd1 _12757_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XDATA\[25\].CLKBUF\[0\] clk vssd1 vssd1 vccd1 vccd1 _09727_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_187_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11707_ _11707_/A _11724_/Y vssd1 vssd1 vccd1 vccd1 _13667_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12687_ _12687_/A _12704_/Y vssd1 vssd1 vccd1 vccd1 _13807_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09649__D line[102] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11638_ _11650_/CLK line[115] vssd1 vssd1 vccd1 vccd1 _11639_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[15\].CLKBUF\[6\] clk vssd1 vssd1 vccd1 vccd1 _06857_/CLK sky130_fd_sc_hd__clkbuf_4
XPHY_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_DATA\[22\].CLKBUF\[5\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12075__D line[64] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11569_ _11569_/A _11584_/Y vssd1 vssd1 vccd1 vccd1 _13809_/Z sky130_fd_sc_hd__ebufn_2
X_13308_ _13330_/CLK line[125] vssd1 vssd1 vccd1 vccd1 _13309_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06073__D line[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05090_ _05090_/A _05109_/Y vssd1 vssd1 vccd1 vccd1 _13770_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11269__A _13933_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12803__D line[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13239_ _13239_/A _13264_/Y vssd1 vssd1 vccd1 vccd1 _13799_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_171_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09384__D line[123] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[14\].VALID\[12\].TOBUF OVHB\[14\].VALID\[12\].FF/Q OVHB\[14\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04929_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_97_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07800_ _07800_/CLK line[25] vssd1 vssd1 vccd1 vccd1 _07801_/A sky130_fd_sc_hd__dfxtp_1
X_08780_ _08780_/CLK line[89] vssd1 vssd1 vccd1 vccd1 _08781_/A sky130_fd_sc_hd__dfxtp_1
X_05992_ _05992_/A _06019_/Y vssd1 vssd1 vccd1 vccd1 _13832_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_111_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MUX.M\[1\].MUX\[4\]_A3 _13832_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07731_ _07731_/A _07734_/Y vssd1 vssd1 vccd1 vccd1 _13891_/Z sky130_fd_sc_hd__ebufn_2
X_04943_ _04965_/CLK line[13] vssd1 vssd1 vccd1 vccd1 _04944_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_38_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07662_ _07662_/CLK _07663_/X vssd1 vssd1 vccd1 vccd1 _07660_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_1_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07632__D line[90] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[15\].VALID\[2\].FF OVHB\[15\].V/CLK A[9] vssd1 vssd1 vccd1 vccd1 OVHB\[15\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_09401_ _09401_/A _09414_/Y vssd1 vssd1 vccd1 vccd1 _13881_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_80_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06613_ _13904_/X wr vssd1 vssd1 vccd1 vccd1 _06613_/X sky130_fd_sc_hd__and2_1
X_07593_ _13911_/X wr vssd1 vssd1 vccd1 vccd1 _07593_/X sky130_fd_sc_hd__and2_1
XANTENNA__11154__D line[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09332_ _09340_/CLK line[85] vssd1 vssd1 vccd1 vccd1 _09333_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_197_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06544_ _13904_/X vssd1 vssd1 vccd1 vccd1 _06544_/Y sky130_fd_sc_hd__inv_2
XANTENNA__06248__D line[83] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09263_ _09263_/A _09274_/Y vssd1 vssd1 vccd1 vccd1 _13743_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[31\].VALID\[11\].FF OVHB\[31\].V/CLK A[18] vssd1 vssd1 vccd1 vccd1 OVHB\[31\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_06475_ _06505_/CLK line[64] vssd1 vssd1 vccd1 vccd1 _06476_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_194_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09559__D line[75] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08214_ _08220_/CLK line[86] vssd1 vssd1 vccd1 vccd1 _08215_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08463__D line[72] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05426_ _05426_/A _05459_/Y vssd1 vssd1 vccd1 vccd1 _13826_/Z sky130_fd_sc_hd__ebufn_2
X_09194_ _09200_/CLK line[22] vssd1 vssd1 vccd1 vccd1 _09195_/A sky130_fd_sc_hd__dfxtp_1
X_08145_ _08145_/A _08154_/Y vssd1 vssd1 vccd1 vccd1 _13745_/Z sky130_fd_sc_hd__ebufn_2
X_05357_ _05385_/CLK line[74] vssd1 vssd1 vccd1 vccd1 _05358_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12563__A _13936_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08076_ _08080_/CLK line[23] vssd1 vssd1 vccd1 vccd1 _08077_/A sky130_fd_sc_hd__dfxtp_1
X_05288_ _05288_/A _05319_/Y vssd1 vssd1 vccd1 vccd1 _13688_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[14\].CLKBUF\[3\] clk vssd1 vssd1 vccd1 vccd1 _06472_/CLK sky130_fd_sc_hd__clkbuf_4
X_07027_ _07027_/A _07034_/Y vssd1 vssd1 vccd1 vccd1 _13747_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_122_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[29\].VALID\[7\].FF_D A[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12713__D line[109] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07807__D line[42] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06711__D line[39] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11329__D line[102] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08978_ _08990_/CLK line[51] vssd1 vssd1 vccd1 vccd1 _08979_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_130_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[6\].INV _13981_/X vssd1 vssd1 vccd1 vccd1 OVHB\[6\].INV/Y sky130_fd_sc_hd__inv_2
X_07929_ _07929_/A _07944_/Y vssd1 vssd1 vccd1 vccd1 _13809_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_152_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XOVHB\[21\].VALID\[13\].FF OVHB\[21\].V/CLK A[20] vssd1 vssd1 vccd1 vccd1 OVHB\[21\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08638__D line[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10940_ _10950_/CLK line[52] vssd1 vssd1 vccd1 vccd1 _10941_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11064__D line[123] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10871_ _10871_/A _10884_/Y vssd1 vssd1 vccd1 vccd1 _13671_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12738__A _13936_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12610_ _12630_/CLK line[62] vssd1 vssd1 vccd1 vccd1 _12611_/A sky130_fd_sc_hd__dfxtp_1
XPHY_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13590_ _13610_/CLK line[126] vssd1 vssd1 vccd1 vccd1 _13591_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05062__D line[53] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12541_ _12541_/A _12564_/Y vssd1 vssd1 vccd1 vccd1 _13661_/Z sky130_fd_sc_hd__ebufn_2
XPHY_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05997__D line[111] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XOVHB\[5\].VALID\[4\].TOBUF OVHB\[5\].VALID\[4\].FF/Q OVHB\[5\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04925_/B2 sky130_fd_sc_hd__ebufn_2
XPHY_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08373__D line[45] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[13\].VALID\[4\].FF OVHB\[13\].V/CLK A[11] vssd1 vssd1 vccd1 vccd1 OVHB\[13\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_12472_ _12490_/CLK line[127] vssd1 vssd1 vccd1 vccd1 _12473_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_200_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11423_ _11423_/A _11444_/Y vssd1 vssd1 vccd1 vccd1 _13663_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_137_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XOVHB\[30\].VALID\[8\].FF OVHB\[30\].V/CLK A[15] vssd1 vssd1 vccd1 vccd1 OVHB\[30\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_165_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11354_ _11370_/CLK line[113] vssd1 vssd1 vccd1 vccd1 _11355_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_4_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10305_ _10305_/A _10324_/Y vssd1 vssd1 vccd1 vccd1 _13665_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_98_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11285_ _11285_/A _11304_/Y vssd1 vssd1 vccd1 vccd1 _13805_/Z sky130_fd_sc_hd__ebufn_2
X_10236_ _10250_/CLK line[114] vssd1 vssd1 vccd1 vccd1 _10237_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06621__D line[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13024_ _13050_/CLK line[123] vssd1 vssd1 vccd1 vccd1 _13025_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11239__D line[75] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10143__D line[72] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDATA\[13\].CLKBUF\[0\] clk vssd1 vssd1 vccd1 vccd1 _06087_/CLK sky130_fd_sc_hd__clkbuf_4
X_10167_ _10167_/A _10184_/Y vssd1 vssd1 vccd1 vccd1 _13807_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05237__D line[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08398__A _13913_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10098_ _10110_/CLK line[51] vssd1 vssd1 vccd1 vccd1 _10099_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_82_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13454__D line[49] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13926_ _13927_/A _13927_/B _13927_/C _13927_/D vssd1 vssd1 vccd1 vccd1 _13926_/X
+ sky130_fd_sc_hd__and4b_4
XANTENNA__08548__D line[125] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13857_ _13857_/CLK _13858_/X vssd1 vssd1 vccd1 vccd1 _13855_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_207_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12808_ _13937_/X wr vssd1 vssd1 vccd1 vccd1 _12808_/X sky130_fd_sc_hd__and2_1
XFILLER_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13788_ _13899_/X wr vssd1 vssd1 vccd1 vccd1 _13788_/X sky130_fd_sc_hd__and2_1
X_12739_ _13936_/X vssd1 vssd1 vccd1 vccd1 _12739_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11702__D line[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06260_ _06260_/CLK line[89] vssd1 vssd1 vccd1 vccd1 _06261_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[29\].VALID\[9\].FF OVHB\[29\].V/CLK A[16] vssd1 vssd1 vccd1 vccd1 OVHB\[29\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__05700__D line[89] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05211_ _05211_/A _05214_/Y vssd1 vssd1 vccd1 vccd1 _13891_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10318__D line[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[21\].CGAND_A _13914_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[2\].CGAND_B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06191_ _06191_/A _06194_/Y vssd1 vssd1 vccd1 vccd1 _13751_/Z sky130_fd_sc_hd__ebufn_2
X_05142_ _05142_/CLK _05143_/X vssd1 vssd1 vccd1 vccd1 _05140_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__13629__D line[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[6\].CGAND_A _13937_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09950_ _09970_/CLK line[126] vssd1 vssd1 vccd1 vccd1 _09951_/A sky130_fd_sc_hd__dfxtp_1
X_05073_ _13931_/Y wr vssd1 vssd1 vccd1 vccd1 _05073_/X sky130_fd_sc_hd__and2_1
XOVHB\[11\].VALID\[6\].FF OVHB\[11\].V/CLK A[13] vssd1 vssd1 vccd1 vccd1 OVHB\[11\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_171_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08901_ _08901_/A _08924_/Y vssd1 vssd1 vccd1 vccd1 _13661_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[20\].CLKBUF\[7\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09881_ _09881_/A _09904_/Y vssd1 vssd1 vccd1 vccd1 _13801_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10053__D line[45] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08832_ _08850_/CLK line[127] vssd1 vssd1 vccd1 vccd1 _08833_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05147__D line[106] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08763_ _08763_/A _08784_/Y vssd1 vssd1 vccd1 vccd1 _13803_/Z sky130_fd_sc_hd__ebufn_2
X_05975_ _05975_/A _05984_/Y vssd1 vssd1 vccd1 vccd1 _13815_/Z sky130_fd_sc_hd__ebufn_2
X_04926_ A_h[6] _04926_/B2 A_h[6] _04926_/B2 vssd1 vssd1 vccd1 vccd1 _04928_/C sky130_fd_sc_hd__a2bb2oi_2
XANTENNA__04986__D line[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07714_ _07730_/CLK line[113] vssd1 vssd1 vccd1 vccd1 _07715_/A sky130_fd_sc_hd__dfxtp_1
X_08694_ _08710_/CLK line[49] vssd1 vssd1 vccd1 vccd1 _08695_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07362__D line[95] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MUX.M\[0\].MUX\[5\]_A1 _13708_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07645_ _07645_/A _07664_/Y vssd1 vssd1 vccd1 vccd1 _13805_/Z sky130_fd_sc_hd__ebufn_2
X_07576_ _07590_/CLK line[50] vssd1 vssd1 vccd1 vccd1 _07577_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_41_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09315_ _09315_/A _09344_/Y vssd1 vssd1 vccd1 vccd1 _13795_/Z sky130_fd_sc_hd__ebufn_2
X_06527_ _06527_/A _06544_/Y vssd1 vssd1 vccd1 vccd1 _13807_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10078__A _13922_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09289__D line[65] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06458_ _06470_/CLK line[51] vssd1 vssd1 vccd1 vccd1 _06459_/A sky130_fd_sc_hd__dfxtp_1
X_09246_ _09270_/CLK line[60] vssd1 vssd1 vccd1 vccd1 _09247_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05610__D line[62] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05409_ _05409_/A _05424_/Y vssd1 vssd1 vccd1 vccd1 _13809_/Z sky130_fd_sc_hd__ebufn_2
X_09177_ _09177_/A _09204_/Y vssd1 vssd1 vccd1 vccd1 _13657_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10228__D line[125] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06389_ _06389_/A _06404_/Y vssd1 vssd1 vccd1 vccd1 _13669_/Z sky130_fd_sc_hd__ebufn_2
X_08128_ _08150_/CLK line[61] vssd1 vssd1 vccd1 vccd1 _08129_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_162_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08059_ _08059_/A _08084_/Y vssd1 vssd1 vccd1 vccd1 _13659_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_134_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12443__D line[99] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07537__D line[47] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11070_ _11090_/CLK line[126] vssd1 vssd1 vccd1 vccd1 _11071_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10021_ _10021_/A _10044_/Y vssd1 vssd1 vccd1 vccd1 _13661_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_49_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09752__D line[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[3\].VALID\[9\].TOBUF OVHB\[3\].VALID\[9\].FF/Q OVHB\[3\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04914_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[1\].VALID\[11\].FF_D A[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11972_ _12000_/CLK line[26] vssd1 vssd1 vccd1 vccd1 _11973_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_56_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13711_ _13715_/CLK line[39] vssd1 vssd1 vccd1 vccd1 _13712_/A sky130_fd_sc_hd__dfxtp_1
X_10923_ _10923_/A _10954_/Y vssd1 vssd1 vccd1 vccd1 _13723_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_16_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13642_ _13642_/A _13649_/Y vssd1 vssd1 vccd1 vccd1 _13642_/Z sky130_fd_sc_hd__ebufn_2
X_10854_ _10880_/CLK line[27] vssd1 vssd1 vccd1 vccd1 _10855_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_72_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12618__D line[51] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13573_ _13575_/CLK line[104] vssd1 vssd1 vccd1 vccd1 _13574_/A sky130_fd_sc_hd__dfxtp_1
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10785_ _10785_/A _10814_/Y vssd1 vssd1 vccd1 vccd1 _13865_/Z sky130_fd_sc_hd__ebufn_2
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12524_ _12524_/A _12529_/Y vssd1 vssd1 vccd1 vccd1 _13644_/Z sky130_fd_sc_hd__ebufn_2
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13299__A _13938_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12455_ _12455_/CLK line[105] vssd1 vssd1 vccd1 vccd1 _12456_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09927__D line[101] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11406_ _11406_/A _11409_/Y vssd1 vssd1 vccd1 vccd1 _13646_/Z sky130_fd_sc_hd__ebufn_2
X_12386_ _12386_/A _12389_/Y vssd1 vssd1 vccd1 vccd1 _13786_/Z sky130_fd_sc_hd__ebufn_2
X_11337_ _11337_/CLK _11338_/X vssd1 vssd1 vccd1 vccd1 _11335_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__06351__D line[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11268_ _13933_/X wr vssd1 vssd1 vccd1 vccd1 _11268_/X sky130_fd_sc_hd__and2_1
XANTENNA_OVHB\[0\].VALID\[1\].FF_D A[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13007_ _13015_/CLK line[101] vssd1 vssd1 vccd1 vccd1 _13008_/A sky130_fd_sc_hd__dfxtp_1
X_10219_ _13922_/X vssd1 vssd1 vccd1 vccd1 _10219_/Y sky130_fd_sc_hd__inv_2
X_11199_ _13933_/X vssd1 vssd1 vccd1 vccd1 _11199_/Y sky130_fd_sc_hd__inv_2
XANTENNA__09662__D line[122] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13184__D line[54] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05760_ _05770_/CLK line[116] vssd1 vssd1 vccd1 vccd1 _05761_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08278__D line[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13909_ _13916_/A _13916_/B _13916_/C _13916_/D vssd1 vssd1 vccd1 vccd1 _13909_/Y
+ sky130_fd_sc_hd__nor4b_4
X_05691_ _05691_/A _05704_/Y vssd1 vssd1 vccd1 vccd1 _13811_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_35_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07430_ _07450_/CLK line[126] vssd1 vssd1 vccd1 vccd1 _07431_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07910__D line[80] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07361_ _07361_/A _07384_/Y vssd1 vssd1 vccd1 vccd1 _13801_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11432__D line[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XOVHB\[10\].VALID\[4\].TOBUF OVHB\[10\].VALID\[4\].FF/Q OVHB\[10\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04925_/B2 sky130_fd_sc_hd__ebufn_2
X_06312_ _06330_/CLK line[127] vssd1 vssd1 vccd1 vccd1 _06313_/A sky130_fd_sc_hd__dfxtp_1
X_09100_ _09130_/CLK line[112] vssd1 vssd1 vccd1 vccd1 _09101_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_31_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07292_ _07310_/CLK line[63] vssd1 vssd1 vccd1 vccd1 _07293_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06526__D line[82] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09031_ _09031_/A _09064_/Y vssd1 vssd1 vccd1 vccd1 _13791_/Z sky130_fd_sc_hd__ebufn_2
X_06243_ _06243_/A _06264_/Y vssd1 vssd1 vccd1 vccd1 _13803_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_175_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06823__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09837__D line[74] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08741__D line[71] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06174_ _06190_/CLK line[49] vssd1 vssd1 vccd1 vccd1 _06175_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13359__D line[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05125_ _05125_/A _05144_/Y vssd1 vssd1 vccd1 vccd1 _13805_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_117_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05056_ _05070_/CLK line[50] vssd1 vssd1 vccd1 vccd1 _05057_/A sky130_fd_sc_hd__dfxtp_1
X_09933_ _09935_/CLK line[104] vssd1 vssd1 vccd1 vccd1 _09934_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_100_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09864_ _09864_/A _09869_/Y vssd1 vssd1 vccd1 vccd1 _13784_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_133_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08815_ _08815_/CLK line[105] vssd1 vssd1 vccd1 vccd1 _08816_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13094__D line[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09795_ _09795_/CLK line[41] vssd1 vssd1 vccd1 vccd1 _09796_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11607__D line[101] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08746_ _08746_/A _08749_/Y vssd1 vssd1 vccd1 vccd1 _13786_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07092__D line[85] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05958_ _05980_/CLK line[93] vssd1 vssd1 vccd1 vccd1 _05959_/A sky130_fd_sc_hd__dfxtp_1
X_05889_ _05889_/A _05914_/Y vssd1 vssd1 vccd1 vccd1 _13729_/Z sky130_fd_sc_hd__ebufn_2
X_08677_ _08677_/CLK _08678_/X vssd1 vssd1 vccd1 vccd1 _08675_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_198_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08916__D line[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07628_ _13911_/X wr vssd1 vssd1 vccd1 vccd1 _07628_/X sky130_fd_sc_hd__and2_1
XFILLER_199_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[0\].CG_CLK clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07559_ _13911_/X vssd1 vssd1 vccd1 vccd1 _07559_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11342__D line[122] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10570_ _10600_/CLK line[16] vssd1 vssd1 vccd1 vccd1 _10571_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05340__D line[52] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09229_ _09235_/CLK line[38] vssd1 vssd1 vccd1 vccd1 _09230_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_181_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XDATA\[5\].CLKBUF\[7\] clk vssd1 vssd1 vccd1 vccd1 _12772_/CLK sky130_fd_sc_hd__clkbuf_4
X_12240_ _12240_/A _12249_/Y vssd1 vssd1 vccd1 vccd1 _13640_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08651__D line[44] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13269__D line[107] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12173__D line[104] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12171_ _12175_/CLK line[103] vssd1 vssd1 vccd1 vccd1 _12172_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07267__D line[37] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[4\].VALID\[14\].TOBUF OVHB\[4\].VALID\[14\].FF/Q OVHB\[4\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/B2 sky130_fd_sc_hd__ebufn_2
X_11122_ _11122_/A _11129_/Y vssd1 vssd1 vccd1 vccd1 _13642_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_3_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11053_ _11055_/CLK line[104] vssd1 vssd1 vccd1 vccd1 _11054_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_89_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10004_ _10004_/A _10009_/Y vssd1 vssd1 vccd1 vccd1 _13644_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_76_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11517__D line[74] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[6\].VALID\[5\].FF_D A[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10421__D line[71] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05515__D line[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_DEC.DEC0.AND2_B A[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[2\].VALID\[1\].FF OVHB\[2\].V/CLK A[8] vssd1 vssd1 vccd1 vccd1 OVHB\[2\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_11955_ _11965_/CLK line[4] vssd1 vssd1 vccd1 vccd1 _11956_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13732__D line[63] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10906_ _10906_/A _10919_/Y vssd1 vssd1 vccd1 vccd1 _13706_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08826__D line[124] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11886_ _11886_/A _11899_/Y vssd1 vssd1 vccd1 vccd1 _13846_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07730__D line[121] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13625_ _13645_/CLK line[14] vssd1 vssd1 vccd1 vccd1 _13626_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12348__D line[56] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10837_ _10845_/CLK line[5] vssd1 vssd1 vccd1 vccd1 _10838_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_9_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XOVHB\[24\].VALID\[10\].TOBUF OVHB\[24\].VALID\[10\].FF/Q OVHB\[24\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04932_/B2 sky130_fd_sc_hd__ebufn_2
X_13556_ _13556_/A _13579_/Y vssd1 vssd1 vccd1 vccd1 _13836_/Z sky130_fd_sc_hd__ebufn_2
X_10768_ _10768_/A _10779_/Y vssd1 vssd1 vccd1 vccd1 _13848_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05250__D line[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12507_ _12525_/CLK line[15] vssd1 vssd1 vccd1 vccd1 _12508_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_146_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13487_ _13505_/CLK line[79] vssd1 vssd1 vccd1 vccd1 _13488_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_8_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10699_ _10705_/CLK line[70] vssd1 vssd1 vccd1 vccd1 _10700_/A sky130_fd_sc_hd__dfxtp_1
X_12438_ _12438_/A _12459_/Y vssd1 vssd1 vccd1 vccd1 _13838_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12083__D line[77] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MUX.M\[2\].MUX\[6\]_A3 _13885_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12369_ _12385_/CLK line[65] vssd1 vssd1 vccd1 vccd1 _12370_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07177__D line[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06081__D line[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XDATA\[4\].CLKBUF\[4\] clk vssd1 vssd1 vccd1 vccd1 _12387_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_114_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06930_ _06960_/CLK line[16] vssd1 vssd1 vccd1 vccd1 _06931_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09392__D line[127] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07905__D line[73] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06861_ _06861_/A _06894_/Y vssd1 vssd1 vccd1 vccd1 _13861_/Z sky130_fd_sc_hd__ebufn_2
X_08600_ _08600_/A _08609_/Y vssd1 vssd1 vccd1 vccd1 _13640_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10331__D line[44] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__04925__A1_N A_h[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05812_ _05840_/CLK line[26] vssd1 vssd1 vccd1 vccd1 _05813_/A sky130_fd_sc_hd__dfxtp_1
X_09580_ _09580_/A _09589_/Y vssd1 vssd1 vccd1 vccd1 _13780_/Z sky130_fd_sc_hd__ebufn_2
X_06792_ _06820_/CLK line[90] vssd1 vssd1 vccd1 vccd1 _06793_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_94_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05425__D line[96] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08531_ _08535_/CLK line[103] vssd1 vssd1 vccd1 vccd1 _08532_/A sky130_fd_sc_hd__dfxtp_1
X_05743_ _05743_/A _05774_/Y vssd1 vssd1 vccd1 vccd1 _13863_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[13\].CLKBUF\[1\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[8\].VALID\[11\].FF_D A[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08462_ _08462_/A _08469_/Y vssd1 vssd1 vccd1 vccd1 _13782_/Z sky130_fd_sc_hd__ebufn_2
X_05674_ _05700_/CLK line[91] vssd1 vssd1 vccd1 vccd1 _05675_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07640__D line[94] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07413_ _07415_/CLK line[104] vssd1 vssd1 vccd1 vccd1 _07414_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12258__D line[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08393_ _08395_/CLK line[40] vssd1 vssd1 vccd1 vccd1 _08394_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_51_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07344_ _07344_/A _07349_/Y vssd1 vssd1 vccd1 vccd1 _13784_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06256__D line[87] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[0\].VALID\[3\].FF OVHB\[0\].V/CLK A[10] vssd1 vssd1 vccd1 vccd1 OVHB\[0\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_149_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07275_ _07275_/CLK line[41] vssd1 vssd1 vccd1 vccd1 _07276_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_148_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09567__D line[79] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06226_ _06226_/A _06229_/Y vssd1 vssd1 vccd1 vccd1 _13786_/Z sky130_fd_sc_hd__ebufn_2
X_09014_ _09014_/A _09029_/Y vssd1 vssd1 vccd1 vccd1 _13774_/Z sky130_fd_sc_hd__ebufn_2
X_06157_ _06157_/CLK _06158_/X vssd1 vssd1 vccd1 vccd1 _06155_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__10506__D line[124] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_DATA\[6\].CLKBUF\[1\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05108_ _13931_/Y wr vssd1 vssd1 vccd1 vccd1 _05108_/X sky130_fd_sc_hd__and2_1
XFILLER_144_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XOVHB\[26\].VALID\[13\].FF OVHB\[26\].V/CLK A[20] vssd1 vssd1 vccd1 vccd1 OVHB\[26\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_06088_ _13903_/X wr vssd1 vssd1 vccd1 vccd1 _06088_/X sky130_fd_sc_hd__and2_1
XANTENNA__12721__D line[98] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05039_ _13931_/Y vssd1 vssd1 vccd1 vccd1 _05039_/Y sky130_fd_sc_hd__inv_2
X_09916_ _09916_/A _09939_/Y vssd1 vssd1 vccd1 vccd1 _13836_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07815__D line[46] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09847_ _09865_/CLK line[79] vssd1 vssd1 vccd1 vccd1 _09848_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_85_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XDATA\[3\].CLKBUF\[1\] clk vssd1 vssd1 vccd1 vccd1 _12002_/CLK sky130_fd_sc_hd__clkbuf_4
X_09778_ _09778_/A _09799_/Y vssd1 vssd1 vccd1 vccd1 _13698_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_39_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05913__A _13902_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08729_ _08745_/CLK line[65] vssd1 vssd1 vccd1 vccd1 _08730_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11740_ _11740_/A _11759_/Y vssd1 vssd1 vccd1 vccd1 _13700_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11671_ _11685_/CLK line[2] vssd1 vssd1 vccd1 vccd1 _11672_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11072__D line[127] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13410_ _13410_/A _13439_/Y vssd1 vssd1 vccd1 vccd1 _13690_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06166__D line[60] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10622_ _10622_/A _10639_/Y vssd1 vssd1 vccd1 vccd1 _13702_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05070__D line[57] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13341_ _13365_/CLK line[12] vssd1 vssd1 vccd1 vccd1 _13342_/A sky130_fd_sc_hd__dfxtp_1
X_10553_ _10565_/CLK line[3] vssd1 vssd1 vccd1 vccd1 _10554_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_139_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[17\].VALID\[4\].TOBUF OVHB\[17\].VALID\[4\].FF/Q OVHB\[17\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04925_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__08381__D line[34] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13272_ _13272_/A _13299_/Y vssd1 vssd1 vccd1 vccd1 _13832_/Z sky130_fd_sc_hd__ebufn_2
X_10484_ _10484_/A _10499_/Y vssd1 vssd1 vccd1 vccd1 _13844_/Z sky130_fd_sc_hd__ebufn_2
X_12223_ _12245_/CLK line[13] vssd1 vssd1 vccd1 vccd1 _12224_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12154_ _12154_/A _12179_/Y vssd1 vssd1 vccd1 vccd1 _13834_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[23\].CLKBUF\[5\] clk vssd1 vssd1 vccd1 vccd1 _09342_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_2_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11105_ _11125_/CLK line[14] vssd1 vssd1 vccd1 vccd1 _11106_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_78_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12085_ _12105_/CLK line[78] vssd1 vssd1 vccd1 vccd1 _12086_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_104_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11036_ _11036_/A _11059_/Y vssd1 vssd1 vccd1 vccd1 _13836_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11247__D line[79] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05245__D line[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09940__D line[112] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13462__D line[53] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12987_ _13015_/CLK line[106] vssd1 vssd1 vccd1 vccd1 _12988_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_205_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08556__D line[114] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11938_ _11938_/A _11969_/Y vssd1 vssd1 vccd1 vccd1 _13618_/Z sky130_fd_sc_hd__ebufn_2
X_11869_ _11895_/CLK line[107] vssd1 vssd1 vccd1 vccd1 _11870_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08853__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13608_ _13610_/CLK line[120] vssd1 vssd1 vccd1 vccd1 _13609_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_60_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05390_ _05420_/CLK line[80] vssd1 vssd1 vccd1 vccd1 _05391_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_186_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13539_ _13539_/A _13544_/Y vssd1 vssd1 vccd1 vccd1 _13819_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11710__D line[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07060_ _07060_/A _07069_/Y vssd1 vssd1 vccd1 vccd1 _13780_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06804__D line[81] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06011_ _06015_/CLK line[103] vssd1 vssd1 vccd1 vccd1 _06012_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_160_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13637__D line[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07962_ _07962_/A _07979_/Y vssd1 vssd1 vccd1 vccd1 _13842_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.M\[1\].MUX\[7\]_A1 _13698_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09701_ _09725_/CLK line[12] vssd1 vssd1 vccd1 vccd1 _09702_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[23\].VALID\[3\].TOBUF OVHB\[23\].VALID\[3\].FF/Q OVHB\[23\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04919_/B2 sky130_fd_sc_hd__ebufn_2
X_06913_ _06925_/CLK line[3] vssd1 vssd1 vccd1 vccd1 _06914_/A sky130_fd_sc_hd__dfxtp_1
X_07893_ _07905_/CLK line[67] vssd1 vssd1 vccd1 vccd1 _07894_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[22\].CLKBUF\[2\] clk vssd1 vssd1 vccd1 vccd1 _08957_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__10061__D line[34] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09632_ _09632_/A _09659_/Y vssd1 vssd1 vccd1 vccd1 _13832_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_55_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06844_ _06844_/A _06859_/Y vssd1 vssd1 vccd1 vccd1 _13844_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[11\].VALID\[1\].FF_D A[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05155__D line[110] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10996__D line[92] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09563_ _09585_/CLK line[77] vssd1 vssd1 vccd1 vccd1 _09564_/A sky130_fd_sc_hd__dfxtp_1
X_06775_ _06785_/CLK line[68] vssd1 vssd1 vccd1 vccd1 _06776_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13372__D line[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__04994__D line[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08514_ _08514_/A _08539_/Y vssd1 vssd1 vccd1 vccd1 _13834_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_130_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13950__A A_h[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05726_ _05726_/A _05739_/Y vssd1 vssd1 vccd1 vccd1 _13846_/Z sky130_fd_sc_hd__ebufn_2
X_09494_ _09494_/A _09519_/Y vssd1 vssd1 vccd1 vccd1 _13694_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07370__D line[84] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08445_ _08465_/CLK line[78] vssd1 vssd1 vccd1 vccd1 _08446_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05657_ _05665_/CLK line[69] vssd1 vssd1 vccd1 vccd1 _05658_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05588_ _05588_/A _05599_/Y vssd1 vssd1 vccd1 vccd1 _13708_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08376_ _08376_/A _08399_/Y vssd1 vssd1 vccd1 vccd1 _13696_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_211_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_DATA\[11\].CLKBUF\[3\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07327_ _07345_/CLK line[79] vssd1 vssd1 vccd1 vccd1 _07328_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_149_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11620__D line[112] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09297__D line[69] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[25\].VALID\[0\].FF OVHB\[25\].V/CLK A[7] vssd1 vssd1 vccd1 vccd1 OVHB\[25\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_07258_ _07258_/A _07279_/Y vssd1 vssd1 vccd1 vccd1 _13698_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10236__D line[114] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06209_ _06225_/CLK line[65] vssd1 vssd1 vccd1 vccd1 _06210_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_136_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07189_ _07205_/CLK line[1] vssd1 vssd1 vccd1 vccd1 _07190_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10814__A _13924_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13547__D line[106] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10533__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12451__D line[103] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[2\].VALID\[8\].FF_D A[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07545__D line[36] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12910_ _12910_/CLK line[57] vssd1 vssd1 vccd1 vccd1 _12911_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_48_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_DATA\[4\].CLKBUF\[3\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13890_ _13890_/CLK line[121] vssd1 vssd1 vccd1 vccd1 _13891_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09760__D line[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XOVHB\[15\].VALID\[9\].TOBUF OVHB\[15\].VALID\[9\].FF/Q OVHB\[15\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04914_/B2 sky130_fd_sc_hd__ebufn_2
X_12841_ _12841_/A _12844_/Y vssd1 vssd1 vccd1 vccd1 _13681_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_64_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12772_ _12772_/CLK _12773_/X vssd1 vssd1 vccd1 vccd1 _12770_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_199_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07280__D line[48] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[30\].CLKBUF\[5\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ _13927_/X wr vssd1 vssd1 vccd1 vccd1 _11723_/X sky130_fd_sc_hd__and2_1
XFILLER_15_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XDATA\[11\].CLKBUF\[5\] clk vssd1 vssd1 vccd1 vccd1 _05702_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_159_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11654_ _13926_/X vssd1 vssd1 vccd1 vccd1 _11654_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06474__A _13904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10708__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10605_ _10635_/CLK line[32] vssd1 vssd1 vccd1 vccd1 _10606_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12626__D line[55] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[22\].VALID\[11\].FF OVHB\[22\].V/CLK A[18] vssd1 vssd1 vccd1 vccd1 OVHB\[22\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11585_ _11615_/CLK line[96] vssd1 vssd1 vccd1 vccd1 _11586_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06193__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13324_ _13330_/CLK line[118] vssd1 vssd1 vccd1 vccd1 _13325_/A sky130_fd_sc_hd__dfxtp_1
X_10536_ _10536_/A _10569_/Y vssd1 vssd1 vccd1 vccd1 _13616_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_183_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13255_ _13255_/A _13264_/Y vssd1 vssd1 vccd1 vccd1 _13815_/Z sky130_fd_sc_hd__ebufn_2
X_10467_ _10495_/CLK line[106] vssd1 vssd1 vccd1 vccd1 _10468_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_89_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09935__D line[105] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12206_ _12210_/CLK line[119] vssd1 vssd1 vccd1 vccd1 _12207_/A sky130_fd_sc_hd__dfxtp_1
X_13186_ _13190_/CLK line[55] vssd1 vssd1 vccd1 vccd1 _13187_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_123_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10398_ _10398_/A _10429_/Y vssd1 vssd1 vccd1 vccd1 _13758_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12361__D line[76] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12137_ _12137_/A _12144_/Y vssd1 vssd1 vccd1 vccd1 _13817_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07455__D line[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[23\].VALID\[2\].FF OVHB\[23\].V/CLK A[9] vssd1 vssd1 vccd1 vccd1 OVHB\[23\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[31\].V_D TIE/HI vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[24\].VALID\[1\].FF_D A[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12068_ _12070_/CLK line[56] vssd1 vssd1 vccd1 vccd1 _12069_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_111_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11019_ _11019_/A _11024_/Y vssd1 vssd1 vccd1 vccd1 _13819_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_37_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06649__A _13905_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09670__D line[126] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06368__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[12\].VALID\[13\].FF OVHB\[12\].V/CLK A[20] vssd1 vssd1 vccd1 vccd1 OVHB\[12\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08286__D line[119] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06560_ _06560_/A _06579_/Y vssd1 vssd1 vccd1 vccd1 _13840_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[17\].VALID\[5\].FF_D A[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05511_ _05525_/CLK line[2] vssd1 vssd1 vccd1 vccd1 _05512_/A sky130_fd_sc_hd__dfxtp_1
X_06491_ _06505_/CLK line[66] vssd1 vssd1 vccd1 vccd1 _06492_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_60_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05442_ _05442_/A _05459_/Y vssd1 vssd1 vccd1 vccd1 _13842_/Z sky130_fd_sc_hd__ebufn_2
X_08230_ _08230_/A _08259_/Y vssd1 vssd1 vccd1 vccd1 _13830_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_60_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12536__D line[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05373_ _05385_/CLK line[67] vssd1 vssd1 vccd1 vccd1 _05374_/A sky130_fd_sc_hd__dfxtp_1
X_08161_ _08185_/CLK line[76] vssd1 vssd1 vccd1 vccd1 _08162_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[21\].VALID\[8\].TOBUF OVHB\[21\].VALID\[8\].FF/Q OVHB\[21\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04931_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_119_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11440__D line[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07112_ _07112_/A _07139_/Y vssd1 vssd1 vccd1 vccd1 _13832_/Z sky130_fd_sc_hd__ebufn_2
X_08092_ _08092_/A _08119_/Y vssd1 vssd1 vccd1 vccd1 _13692_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[10\].CLKBUF\[2\] clk vssd1 vssd1 vccd1 vccd1 _05317_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__06534__D line[86] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07043_ _07065_/CLK line[77] vssd1 vssd1 vccd1 vccd1 _07044_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_161_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09845__D line[78] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08994_ _13915_/X vssd1 vssd1 vccd1 vccd1 _08994_/Y sky130_fd_sc_hd__inv_2
XANTENNA__07943__A _13912_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07945_ _07975_/CLK line[96] vssd1 vssd1 vccd1 vccd1 _07946_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_55_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07876_ _07876_/A _07909_/Y vssd1 vssd1 vccd1 vccd1 _13756_/Z sky130_fd_sc_hd__ebufn_2
X_09615_ _09615_/A _09624_/Y vssd1 vssd1 vccd1 vccd1 _13815_/Z sky130_fd_sc_hd__ebufn_2
X_06827_ _06855_/CLK line[106] vssd1 vssd1 vccd1 vccd1 _06828_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_55_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11615__D line[105] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[29\].CLKBUF\[6\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06709__D line[38] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09546_ _09550_/CLK line[55] vssd1 vssd1 vccd1 vccd1 _09547_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[21\].VALID\[4\].FF OVHB\[21\].V/CLK A[11] vssd1 vssd1 vccd1 vccd1 OVHB\[21\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08196__D line[92] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06758_ _06758_/A _06789_/Y vssd1 vssd1 vccd1 vccd1 _13758_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_36_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05709_ _05735_/CLK line[107] vssd1 vssd1 vccd1 vccd1 _05710_/A sky130_fd_sc_hd__dfxtp_1
XPHY_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09477_ _09477_/A _09484_/Y vssd1 vssd1 vccd1 vccd1 _13677_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_169_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06689_ _06715_/CLK line[43] vssd1 vssd1 vccd1 vccd1 _06690_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_169_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08428_ _08430_/CLK line[56] vssd1 vssd1 vccd1 vccd1 _08429_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08359_ _08359_/A _08364_/Y vssd1 vssd1 vccd1 vccd1 _13679_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11350__D line[126] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[15\].VALID\[13\].FF_D A[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XOVHB\[25\].CG clk OVHB\[25\].CGAND/X vssd1 vssd1 vccd1 vccd1 OVHB\[25\].V/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_149_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06444__D line[59] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11370_ _11370_/CLK line[121] vssd1 vssd1 vccd1 vccd1 _11371_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_50_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10321_ _10321_/A _10324_/Y vssd1 vssd1 vccd1 vccd1 _13681_/Z sky130_fd_sc_hd__ebufn_2
X_13040_ _13050_/CLK line[116] vssd1 vssd1 vccd1 vccd1 _13041_/A sky130_fd_sc_hd__dfxtp_1
X_10252_ _10252_/CLK _10253_/X vssd1 vssd1 vccd1 vccd1 _10250_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08014__A _13912_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13277__D line[111] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10183_ _13922_/X wr vssd1 vssd1 vccd1 vccd1 _10183_/X sky130_fd_sc_hd__and2_1
XOVHB\[17\].VALID\[14\].TOBUF OVHB\[17\].VALID\[14\].FF/Q OVHB\[17\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__07275__D line[41] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_OVHB\[25\].VALID\[12\].FF_D A[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[5\].VALID\[0\].TOBUF OVHB\[5\].VALID\[0\].FF/Q OVHB\[5\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04924_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_47_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13942_ _13949_/A _13949_/B _13949_/C _13949_/D vssd1 vssd1 vccd1 vccd1 _13942_/Y
+ sky130_fd_sc_hd__nor4b_4
XFILLER_46_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13873_ _13873_/A _13894_/Y vssd1 vssd1 vccd1 vccd1 _13873_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_74_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11525__D line[78] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12824_ _12840_/CLK line[17] vssd1 vssd1 vccd1 vccd1 _12825_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06619__D line[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[1\].V_D TIE/HI vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05523__D line[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12755_ _12755_/A _12774_/Y vssd1 vssd1 vccd1 vccd1 _13875_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13740__D line[52] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[2\].CLKBUF\[5\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11706_ _11720_/CLK line[18] vssd1 vssd1 vccd1 vccd1 _11707_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08834__D line[113] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12686_ _12700_/CLK line[82] vssd1 vssd1 vccd1 vccd1 _12687_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11637_ _11637_/A _11654_/Y vssd1 vssd1 vccd1 vccd1 _13877_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[10\].VALID\[13\].TOBUF OVHB\[10\].VALID\[13\].FF/Q OVHB\[10\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04916_/B2 sky130_fd_sc_hd__ebufn_2
X_11568_ _11580_/CLK line[83] vssd1 vssd1 vccd1 vccd1 _11569_/A sky130_fd_sc_hd__dfxtp_1
X_13307_ _13307_/A _13334_/Y vssd1 vssd1 vccd1 vccd1 _13867_/Z sky130_fd_sc_hd__ebufn_2
X_10519_ _10519_/A _10534_/Y vssd1 vssd1 vccd1 vccd1 _13879_/Z sky130_fd_sc_hd__ebufn_2
X_11499_ _11499_/A _11514_/Y vssd1 vssd1 vccd1 vccd1 _13739_/Z sky130_fd_sc_hd__ebufn_2
X_13238_ _13260_/CLK line[93] vssd1 vssd1 vccd1 vccd1 _13239_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12091__D line[66] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13169_ _13169_/A _13194_/Y vssd1 vssd1 vccd1 vccd1 _13729_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07185__D line[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05991_ _06015_/CLK line[108] vssd1 vssd1 vccd1 vccd1 _05992_/A sky130_fd_sc_hd__dfxtp_1
X_07730_ _07730_/CLK line[121] vssd1 vssd1 vccd1 vccd1 _07731_/A sky130_fd_sc_hd__dfxtp_1
X_04942_ _04942_/A _04969_/Y vssd1 vssd1 vccd1 vccd1 _13622_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_65_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05283__A _13900_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07661_ _07661_/A _07664_/Y vssd1 vssd1 vccd1 vccd1 _13821_/Z sky130_fd_sc_hd__ebufn_2
X_09400_ _09410_/CLK line[116] vssd1 vssd1 vccd1 vccd1 _09401_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_1_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06612_ _06612_/CLK _06613_/X vssd1 vssd1 vccd1 vccd1 _06610_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_198_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07592_ _07592_/CLK _07593_/X vssd1 vssd1 vccd1 vccd1 _07590_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_34_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05433__D line[109] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09331_ _09331_/A _09344_/Y vssd1 vssd1 vccd1 vccd1 _13811_/Z sky130_fd_sc_hd__ebufn_2
X_06543_ _13904_/X wr vssd1 vssd1 vccd1 vccd1 _06543_/X sky130_fd_sc_hd__and2_1
XANTENNA__13650__D line[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09262_ _09270_/CLK line[53] vssd1 vssd1 vccd1 vccd1 _09263_/A sky130_fd_sc_hd__dfxtp_1
X_06474_ _13904_/X vssd1 vssd1 vccd1 vccd1 _06474_/Y sky130_fd_sc_hd__inv_2
XOVHB\[18\].VALID\[7\].FF OVHB\[18\].V/CLK A[14] vssd1 vssd1 vccd1 vccd1 OVHB\[18\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_08213_ _08213_/A _08224_/Y vssd1 vssd1 vccd1 vccd1 _13813_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_21_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12266__D line[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05425_ _05455_/CLK line[96] vssd1 vssd1 vccd1 vccd1 _05426_/A sky130_fd_sc_hd__dfxtp_1
X_09193_ _09193_/A _09204_/Y vssd1 vssd1 vccd1 vccd1 _13673_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_166_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12844__A _13937_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05356_ _05356_/A _05389_/Y vssd1 vssd1 vccd1 vccd1 _13756_/Z sky130_fd_sc_hd__ebufn_2
X_08144_ _08150_/CLK line[54] vssd1 vssd1 vccd1 vccd1 _08145_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_147_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12563__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08075_ _08075_/A _08084_/Y vssd1 vssd1 vccd1 vccd1 _13675_/Z sky130_fd_sc_hd__ebufn_2
X_05287_ _05315_/CLK line[42] vssd1 vssd1 vccd1 vccd1 _05288_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[20\].INV _13957_/X vssd1 vssd1 vccd1 vccd1 OVHB\[20\].INV/Y sky130_fd_sc_hd__inv_2
XANTENNA__09575__D line[68] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07026_ _07030_/CLK line[55] vssd1 vssd1 vccd1 vccd1 _07027_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05458__A _13900_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10514__D line[113] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05608__D line[61] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08977_ _08977_/A _08994_/Y vssd1 vssd1 vccd1 vccd1 _13737_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13825__D line[96] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07928_ _07940_/CLK line[83] vssd1 vssd1 vccd1 vccd1 _07929_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_28_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07823__D line[35] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07859_ _07859_/A _07874_/Y vssd1 vssd1 vccd1 vccd1 _13739_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_16_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10870_ _10880_/CLK line[20] vssd1 vssd1 vccd1 vccd1 _10871_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_28_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XOVHB\[30\].VALID\[13\].TOBUF OVHB\[30\].VALID\[13\].FF/Q OVHB\[30\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04916_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__12738__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09529_ _09529_/A _09554_/Y vssd1 vssd1 vccd1 vccd1 _13729_/Z sky130_fd_sc_hd__ebufn_2
XPHY_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12540_ _12560_/CLK line[30] vssd1 vssd1 vccd1 vccd1 _12541_/A sky130_fd_sc_hd__dfxtp_1
XPHY_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12471_ _12471_/A _12494_/Y vssd1 vssd1 vccd1 vccd1 _13871_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_200_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11080__D line[116] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[3\].VALID\[5\].TOBUF OVHB\[3\].VALID\[5\].FF/Q OVHB\[3\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04927_/B2 sky130_fd_sc_hd__ebufn_2
X_11422_ _11440_/CLK line[31] vssd1 vssd1 vccd1 vccd1 _11423_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06174__D line[49] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[28\].VALID\[8\].TOBUF OVHB\[28\].VALID\[8\].FF/Q OVHB\[28\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04931_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__12904__D line[54] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11353_ _11353_/A _11374_/Y vssd1 vssd1 vccd1 vccd1 _13873_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_4_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09485__D line[32] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10304_ _10320_/CLK line[17] vssd1 vssd1 vccd1 vccd1 _10305_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[16\].VALID\[9\].FF OVHB\[16\].V/CLK A[16] vssd1 vssd1 vccd1 vccd1 OVHB\[16\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_152_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11284_ _11300_/CLK line[81] vssd1 vssd1 vccd1 vccd1 _11285_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_112_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_OVHB\[20\].VALID\[4\].FF_D A[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13023_ _13023_/A _13054_/Y vssd1 vssd1 vccd1 vccd1 _13863_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_180_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10235_ _10235_/A _10254_/Y vssd1 vssd1 vccd1 vccd1 _13875_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_106_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08679__A _13914_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10166_ _10180_/CLK line[82] vssd1 vssd1 vccd1 vccd1 _10167_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08398__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10097_ _10097_/A _10114_/Y vssd1 vssd1 vccd1 vccd1 _13737_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_19_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13925_ _13927_/B _13927_/A _13927_/C _13927_/D vssd1 vssd1 vccd1 vccd1 _13925_/X
+ sky130_fd_sc_hd__and4b_4
XANTENNA_OVHB\[13\].VALID\[8\].FF_D A[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11255__D line[68] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06349__D line[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13856_ _13856_/A _13859_/Y vssd1 vssd1 vccd1 vccd1 _13856_/Z sky130_fd_sc_hd__ebufn_2
X_12807_ _12807_/CLK _12808_/X vssd1 vssd1 vccd1 vccd1 _12805_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_62_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13787_ _13787_/CLK _13788_/X vssd1 vssd1 vccd1 vccd1 _13785_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__13470__D line[57] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10999_ _10999_/A _11024_/Y vssd1 vssd1 vccd1 vccd1 _13799_/Z sky130_fd_sc_hd__ebufn_2
X_12738_ _13936_/X wr vssd1 vssd1 vccd1 vccd1 _12738_/X sky130_fd_sc_hd__and2_1
XANTENNA__08564__D line[118] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12669_ _13936_/X vssd1 vssd1 vccd1 vccd1 _12669_/Y sky130_fd_sc_hd__inv_2
XPHY_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05210_ _05210_/CLK line[121] vssd1 vssd1 vccd1 vccd1 _05211_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_175_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06190_ _06190_/CLK line[57] vssd1 vssd1 vccd1 vccd1 _06191_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[21\].CGAND_B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05141_ _05141_/A _05144_/Y vssd1 vssd1 vccd1 vccd1 _13821_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[3\].V OVHB\[3\].V/CLK TIE/HI rst_n vssd1 vssd1 vccd1 vccd1 OVHB\[3\].V/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12814__D line[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_DATA\[0\].CLKBUF\[7\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10184__A _13922_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09973__A _13921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05072_ _05072_/CLK _05073_/X vssd1 vssd1 vccd1 vccd1 _05070_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA_OVHB\[6\].CGAND_B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06812__D line[85] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[25\].CGAND_A _13921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08900_ _08920_/CLK line[30] vssd1 vssd1 vccd1 vccd1 _08901_/A sky130_fd_sc_hd__dfxtp_1
X_09880_ _09900_/CLK line[94] vssd1 vssd1 vccd1 vccd1 _09881_/A sky130_fd_sc_hd__dfxtp_1
X_08831_ _08831_/A _08854_/Y vssd1 vssd1 vccd1 vccd1 _13871_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[10\].VALID\[0\].TOBUF OVHB\[10\].VALID\[0\].FF/Q OVHB\[10\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04924_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_97_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13645__D line[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08739__D line[70] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08762_ _08780_/CLK line[95] vssd1 vssd1 vccd1 vccd1 _08763_/A sky130_fd_sc_hd__dfxtp_1
X_05974_ _05980_/CLK line[86] vssd1 vssd1 vccd1 vccd1 _05975_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[3\].VALID\[13\].FF OVHB\[3\].V/CLK A[20] vssd1 vssd1 vccd1 vccd1 OVHB\[3\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_07713_ _07713_/A _07734_/Y vssd1 vssd1 vccd1 vccd1 _13873_/Z sky130_fd_sc_hd__ebufn_2
X_04925_ A_h[9] _04925_/B2 A_h[9] _04925_/B2 vssd1 vssd1 vccd1 vccd1 _04928_/B sky130_fd_sc_hd__a2bb2oi_2
X_08693_ _08693_/A _08714_/Y vssd1 vssd1 vccd1 vccd1 _13733_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11165__D line[32] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07644_ _07660_/CLK line[81] vssd1 vssd1 vccd1 vccd1 _07645_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.M\[0\].MUX\[5\]_A2 _13778_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05163__D line[99] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07575_ _07575_/A _07594_/Y vssd1 vssd1 vccd1 vccd1 _13735_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13380__D line[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10359__A _13923_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09314_ _09340_/CLK line[91] vssd1 vssd1 vccd1 vccd1 _09315_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08474__D line[91] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06526_ _06540_/CLK line[82] vssd1 vssd1 vccd1 vccd1 _06527_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_179_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10078__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09245_ _09245_/A _09274_/Y vssd1 vssd1 vccd1 vccd1 _13725_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_193_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06457_ _06457_/A _06474_/Y vssd1 vssd1 vccd1 vccd1 _13737_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[1\].CLKBUF\[6\] clk vssd1 vssd1 vccd1 vccd1 _08257_/CLK sky130_fd_sc_hd__clkbuf_4
X_05408_ _05420_/CLK line[83] vssd1 vssd1 vccd1 vccd1 _05409_/A sky130_fd_sc_hd__dfxtp_1
X_09176_ _09200_/CLK line[28] vssd1 vssd1 vccd1 vccd1 _09177_/A sky130_fd_sc_hd__dfxtp_1
X_06388_ _06400_/CLK line[19] vssd1 vssd1 vccd1 vccd1 _06389_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_5_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08127_ _08127_/A _08154_/Y vssd1 vssd1 vccd1 vccd1 _13727_/Z sky130_fd_sc_hd__ebufn_2
X_05339_ _05339_/A _05354_/Y vssd1 vssd1 vccd1 vccd1 _13739_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_134_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06722__D line[58] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08058_ _08080_/CLK line[29] vssd1 vssd1 vccd1 vccd1 _08059_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10244__D line[118] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07009_ _07009_/A _07034_/Y vssd1 vssd1 vccd1 vccd1 _13729_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_162_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[31\].VOBUF OVHB\[31\].V/Q OVHB\[31\].INV/Y vssd1 vssd1 vccd1 vccd1 _04912_/B1
+ sky130_fd_sc_hd__ebufn_2
XFILLER_0_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05338__D line[51] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10020_ _10040_/CLK line[30] vssd1 vssd1 vccd1 vccd1 _10021_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13555__D line[110] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_OVHB\[26\].VALID\[8\].FF_D A[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08649__D line[43] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07553__D line[40] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XDATA\[31\].CLKBUF\[4\] clk vssd1 vssd1 vccd1 vccd1 _11827_/CLK sky130_fd_sc_hd__clkbuf_4
X_11971_ _11971_/A _12004_/Y vssd1 vssd1 vccd1 vccd1 _13651_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_56_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13710_ _13710_/A _13719_/Y vssd1 vssd1 vccd1 vccd1 _13710_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11653__A _13926_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10922_ _10950_/CLK line[58] vssd1 vssd1 vccd1 vccd1 _10923_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_72_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XOVHB\[27\].VALID\[11\].FF OVHB\[27\].V/CLK A[18] vssd1 vssd1 vccd1 vccd1 OVHB\[27\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_72_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13641_ _13645_/CLK line[7] vssd1 vssd1 vccd1 vccd1 _13642_/A sky130_fd_sc_hd__dfxtp_1
X_10853_ _10853_/A _10884_/Y vssd1 vssd1 vccd1 vccd1 _13653_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_31_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XOVHB\[4\].VALID\[10\].TOBUF OVHB\[4\].VALID\[10\].FF/Q OVHB\[4\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04932_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_13_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11803__D line[77] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13572_ _13572_/A _13579_/Y vssd1 vssd1 vccd1 vccd1 _13852_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_31_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10784_ _10810_/CLK line[123] vssd1 vssd1 vccd1 vccd1 _10785_/A sky130_fd_sc_hd__dfxtp_1
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05801__D line[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12523_ _12525_/CLK line[8] vssd1 vssd1 vccd1 vccd1 _12524_/A sky130_fd_sc_hd__dfxtp_1
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10419__D line[70] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12454_ _12454_/A _12459_/Y vssd1 vssd1 vccd1 vccd1 _13854_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_138_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11405_ _11405_/CLK line[9] vssd1 vssd1 vccd1 vccd1 _11406_/A sky130_fd_sc_hd__dfxtp_1
X_12385_ _12385_/CLK line[73] vssd1 vssd1 vccd1 vccd1 _12386_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_125_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XDATA\[0\].CLKBUF\[3\] clk vssd1 vssd1 vccd1 vccd1 _05072_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__07728__D line[120] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11336_ _11336_/A _11339_/Y vssd1 vssd1 vccd1 vccd1 _13856_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_4_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10154__D line[91] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11828__A _13927_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[9\].VALID\[2\].FF OVHB\[9\].V/CLK A[9] vssd1 vssd1 vccd1 vccd1 OVHB\[9\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_11267_ _11267_/CLK _11268_/X vssd1 vssd1 vccd1 vccd1 _11265_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_97_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13006_ _13006_/A _13019_/Y vssd1 vssd1 vccd1 vccd1 _13846_/Z sky130_fd_sc_hd__ebufn_2
X_10218_ _13922_/X wr vssd1 vssd1 vccd1 vccd1 _10218_/X sky130_fd_sc_hd__and2_1
XANTENNA_DATA\[21\].CLKBUF\[1\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11198_ _13933_/X wr vssd1 vssd1 vccd1 vccd1 _11198_/X sky130_fd_sc_hd__and2_1
XOVHB\[17\].VALID\[13\].FF OVHB\[17\].V/CLK A[20] vssd1 vssd1 vccd1 vccd1 OVHB\[17\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_10149_ _13922_/X vssd1 vssd1 vccd1 vccd1 _10149_/Y sky130_fd_sc_hd__inv_2
XANTENNA__07463__D line[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06079__D line[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13908_ A[4] vssd1 vssd1 vccd1 vccd1 _13916_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_62_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05690_ _05700_/CLK line[84] vssd1 vssd1 vccd1 vccd1 _05691_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_23_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13839_ _13855_/CLK line[97] vssd1 vssd1 vccd1 vccd1 _13840_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[30\].CLKBUF\[1\] clk vssd1 vssd1 vccd1 vccd1 _11442_/CLK sky130_fd_sc_hd__clkbuf_4
X_07360_ _07380_/CLK line[94] vssd1 vssd1 vccd1 vccd1 _07361_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05711__D line[108] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[7\].VALID\[3\].FF_D A[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06311_ _06311_/A _06334_/Y vssd1 vssd1 vccd1 vccd1 _13871_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_188_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10329__D line[43] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDATA\[20\].CLKBUF\[7\] clk vssd1 vssd1 vccd1 vccd1 _08572_/CLK sky130_fd_sc_hd__clkbuf_4
X_07291_ _07291_/A _07314_/Y vssd1 vssd1 vccd1 vccd1 _13731_/Z sky130_fd_sc_hd__ebufn_2
X_09030_ _09060_/CLK line[80] vssd1 vssd1 vccd1 vccd1 _09031_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07488__A _13911_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06242_ _06260_/CLK line[95] vssd1 vssd1 vccd1 vccd1 _06243_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[5\].INV _13980_/X vssd1 vssd1 vccd1 vccd1 OVHB\[5\].INV/Y sky130_fd_sc_hd__inv_2
XFILLER_175_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12544__D line[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06173_ _06173_/A _06194_/Y vssd1 vssd1 vccd1 vccd1 _13733_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_7_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07638__D line[93] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05124_ _05140_/CLK line[81] vssd1 vssd1 vccd1 vccd1 _05125_/A sky130_fd_sc_hd__dfxtp_1
XMUX.SEL1BUF\[0\] A[1] vssd1 vssd1 vccd1 vccd1 MUX.SEL1BUF\[0\]/X sky130_fd_sc_hd__clkbuf_2
XFILLER_117_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05055_ _05055_/A _05074_/Y vssd1 vssd1 vccd1 vccd1 _13735_/Z sky130_fd_sc_hd__ebufn_2
X_09932_ _09932_/A _09939_/Y vssd1 vssd1 vccd1 vccd1 _13852_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09853__D line[67] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09863_ _09865_/CLK line[72] vssd1 vssd1 vccd1 vccd1 _09864_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_97_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08814_ _08814_/A _08819_/Y vssd1 vssd1 vccd1 vccd1 _13854_/Z sky130_fd_sc_hd__ebufn_2
X_09794_ _09794_/A _09799_/Y vssd1 vssd1 vccd1 vccd1 _13714_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_39_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08745_ _08745_/CLK line[73] vssd1 vssd1 vccd1 vccd1 _08746_/A sky130_fd_sc_hd__dfxtp_1
X_05957_ _05957_/A _05984_/Y vssd1 vssd1 vccd1 vccd1 _13797_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_26_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[7\].VALID\[4\].FF OVHB\[7\].V/CLK A[11] vssd1 vssd1 vccd1 vccd1 OVHB\[7\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_08676_ _08676_/A _08679_/Y vssd1 vssd1 vccd1 vccd1 _13716_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_199_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05888_ _05910_/CLK line[61] vssd1 vssd1 vccd1 vccd1 _05889_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_198_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07627_ _07627_/CLK _07628_/X vssd1 vssd1 vccd1 vccd1 _07625_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__12719__D line[97] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07558_ _13911_/X wr vssd1 vssd1 vccd1 vccd1 _07558_/X sky130_fd_sc_hd__and2_1
XPHY_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06509_ _13904_/X vssd1 vssd1 vccd1 vccd1 _06509_/Y sky130_fd_sc_hd__inv_2
XOVHB\[27\].VALID\[12\].TOBUF OVHB\[27\].VALID\[12\].FF/Q OVHB\[27\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04929_/B2 sky130_fd_sc_hd__ebufn_2
X_07489_ _13911_/X vssd1 vssd1 vccd1 vccd1 _07489_/Y sky130_fd_sc_hd__inv_2
XFILLER_166_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09228_ _09228_/A _09239_/Y vssd1 vssd1 vccd1 vccd1 _13708_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_167_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09159_ _09165_/CLK line[6] vssd1 vssd1 vccd1 vccd1 _09160_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_182_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06452__D line[63] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12170_ _12170_/A _12179_/Y vssd1 vssd1 vccd1 vccd1 _13850_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11121_ _11125_/CLK line[7] vssd1 vssd1 vccd1 vccd1 _11122_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_89_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05068__D line[56] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11052_ _11052_/A _11059_/Y vssd1 vssd1 vccd1 vccd1 _13852_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13285__D line[100] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10003_ _10005_/CLK line[8] vssd1 vssd1 vccd1 vccd1 _10004_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08379__D line[33] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[17\].VALID\[0\].TOBUF OVHB\[17\].VALID\[0\].FF/Q OVHB\[17\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04924_/B2 sky130_fd_sc_hd__ebufn_2
X_11954_ _11954_/A _11969_/Y vssd1 vssd1 vccd1 vccd1 _13634_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[20\].VALID\[11\].TOBUF OVHB\[20\].VALID\[11\].FF/Q OVHB\[20\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04915_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_44_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10905_ _10915_/CLK line[36] vssd1 vssd1 vccd1 vccd1 _10906_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_44_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11885_ _11895_/CLK line[100] vssd1 vssd1 vccd1 vccd1 _11886_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_189_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11533__D line[67] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13624_ _13624_/A _13649_/Y vssd1 vssd1 vccd1 vccd1 _13624_/Z sky130_fd_sc_hd__ebufn_2
X_10836_ _10836_/A _10849_/Y vssd1 vssd1 vccd1 vccd1 _13636_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06627__D line[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09003__D line[77] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[5\].VALID\[6\].FF OVHB\[5\].V/CLK A[13] vssd1 vssd1 vccd1 vccd1 OVHB\[5\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_13555_ _13575_/CLK line[110] vssd1 vssd1 vccd1 vccd1 _13556_/A sky130_fd_sc_hd__dfxtp_1
X_10767_ _10775_/CLK line[101] vssd1 vssd1 vccd1 vccd1 _10768_/A sky130_fd_sc_hd__dfxtp_1
X_12506_ _12506_/A _12529_/Y vssd1 vssd1 vccd1 vccd1 _13626_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08842__D line[117] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13486_ _13486_/A _13509_/Y vssd1 vssd1 vccd1 vccd1 _13766_/Z sky130_fd_sc_hd__ebufn_2
X_10698_ _10698_/A _10709_/Y vssd1 vssd1 vccd1 vccd1 _13778_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_172_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12437_ _12455_/CLK line[111] vssd1 vssd1 vccd1 vccd1 _12438_/A sky130_fd_sc_hd__dfxtp_1
X_12368_ _12368_/A _12389_/Y vssd1 vssd1 vccd1 vccd1 _13768_/Z sky130_fd_sc_hd__ebufn_2
X_11319_ _11335_/CLK line[97] vssd1 vssd1 vccd1 vccd1 _11320_/A sky130_fd_sc_hd__dfxtp_1
X_12299_ _12315_/CLK line[33] vssd1 vssd1 vccd1 vccd1 _12300_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09028__A _13915_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11708__D line[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13195__D line[64] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06860_ _06890_/CLK line[112] vssd1 vssd1 vccd1 vccd1 _06861_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07193__D line[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05811_ _05811_/A _05844_/Y vssd1 vssd1 vccd1 vccd1 _13651_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_83_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06791_ _06791_/A _06824_/Y vssd1 vssd1 vccd1 vccd1 _13791_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12389__A _13935_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08530_ _08530_/A _08539_/Y vssd1 vssd1 vccd1 vccd1 _13850_/Z sky130_fd_sc_hd__ebufn_2
X_05742_ _05770_/CLK line[122] vssd1 vssd1 vccd1 vccd1 _05743_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_35_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08461_ _08465_/CLK line[71] vssd1 vssd1 vccd1 vccd1 _08462_/A sky130_fd_sc_hd__dfxtp_1
X_05673_ _05673_/A _05704_/Y vssd1 vssd1 vccd1 vccd1 _13793_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_50_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07412_ _07412_/A _07419_/Y vssd1 vssd1 vccd1 vccd1 _13852_/Z sky130_fd_sc_hd__ebufn_2
X_08392_ _08392_/A _08399_/Y vssd1 vssd1 vccd1 vccd1 _13712_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05441__D line[98] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07343_ _07345_/CLK line[72] vssd1 vssd1 vccd1 vccd1 _07344_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10059__D line[33] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08752__D line[90] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07274_ _07274_/A _07279_/Y vssd1 vssd1 vccd1 vccd1 _13714_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[20\].CG_CLK clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09013_ _09025_/CLK line[67] vssd1 vssd1 vccd1 vccd1 _09014_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12274__D line[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06225_ _06225_/CLK line[73] vssd1 vssd1 vccd1 vccd1 _06226_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_117_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XOVHB\[13\].VALID\[11\].FF OVHB\[13\].V/CLK A[18] vssd1 vssd1 vccd1 vccd1 OVHB\[13\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07368__D line[83] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06156_ _06156_/A _06159_/Y vssd1 vssd1 vccd1 vccd1 _13716_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[3\].VALID\[8\].FF OVHB\[3\].V/CLK A[15] vssd1 vssd1 vccd1 vccd1 OVHB\[3\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_05107_ _05107_/CLK _05108_/X vssd1 vssd1 vccd1 vccd1 _05105_/CLK sky130_fd_sc_hd__dlclkp_1
X_06087_ _06087_/CLK _06088_/X vssd1 vssd1 vccd1 vccd1 _06085_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__09583__D line[72] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05038_ _13931_/Y wr vssd1 vssd1 vccd1 vccd1 _05038_/X sky130_fd_sc_hd__and2_1
X_09915_ _09935_/CLK line[110] vssd1 vssd1 vccd1 vccd1 _09916_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13683__A _13899_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10522__D line[117] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09846_ _09846_/A _09869_/Y vssd1 vssd1 vccd1 vccd1 _13766_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05616__D line[50] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09777_ _09795_/CLK line[47] vssd1 vssd1 vccd1 vccd1 _09778_/A sky130_fd_sc_hd__dfxtp_1
X_06989_ _06995_/CLK line[38] vssd1 vssd1 vccd1 vccd1 _06990_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13833__D line[109] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08728_ _08728_/A _08749_/Y vssd1 vssd1 vccd1 vccd1 _13768_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05913__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08927__D line[42] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[2\].VALID\[12\].FF_D A[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07831__D line[39] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08659_ _08675_/CLK line[33] vssd1 vssd1 vccd1 vccd1 _08660_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12449__D line[102] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11670_ _11670_/A _11689_/Y vssd1 vssd1 vccd1 vccd1 _13630_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10621_ _10635_/CLK line[34] vssd1 vssd1 vccd1 vccd1 _10622_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09758__D line[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13340_ _13340_/A _13369_/Y vssd1 vssd1 vccd1 vccd1 _13620_/Z sky130_fd_sc_hd__ebufn_2
X_10552_ _10552_/A _10569_/Y vssd1 vssd1 vccd1 vccd1 _13632_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12184__D line[123] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13271_ _13295_/CLK line[108] vssd1 vssd1 vccd1 vccd1 _13272_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13858__A _13899_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10483_ _10495_/CLK line[99] vssd1 vssd1 vccd1 vccd1 _10484_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[15\].VALID\[5\].TOBUF OVHB\[15\].VALID\[5\].FF/Q OVHB\[15\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04927_/B2 sky130_fd_sc_hd__ebufn_2
XOVHB\[31\].VALID\[2\].FF OVHB\[31\].V/CLK A[9] vssd1 vssd1 vccd1 vccd1 OVHB\[31\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_12222_ _12222_/A _12249_/Y vssd1 vssd1 vccd1 vccd1 _13622_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06182__D line[53] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12153_ _12175_/CLK line[109] vssd1 vssd1 vccd1 vccd1 _12154_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_78_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09493__D line[45] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11104_ _11104_/A _11129_/Y vssd1 vssd1 vccd1 vccd1 _13624_/Z sky130_fd_sc_hd__ebufn_2
X_12084_ _12084_/A _12109_/Y vssd1 vssd1 vccd1 vccd1 _13764_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_123_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10432__D line[90] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11035_ _11055_/CLK line[110] vssd1 vssd1 vccd1 vccd1 _11036_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_76_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[9\].V_RESET_B rst_n vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[18\].CLKBUF\[4\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12986_ _12986_/A _13019_/Y vssd1 vssd1 vccd1 vccd1 _13826_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07741__D line[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12359__D line[75] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11937_ _11965_/CLK line[10] vssd1 vssd1 vccd1 vccd1 _11938_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[3\].VALID\[6\].FF_D A[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11263__D line[72] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06357__D line[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11868_ _11868_/A _11899_/Y vssd1 vssd1 vccd1 vccd1 _13828_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_32_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10819_ _10845_/CLK line[11] vssd1 vssd1 vccd1 vccd1 _10820_/A sky130_fd_sc_hd__dfxtp_1
X_13607_ _13607_/A _13614_/Y vssd1 vssd1 vccd1 vccd1 _13887_/Z sky130_fd_sc_hd__ebufn_2
X_11799_ _11825_/CLK line[75] vssd1 vssd1 vccd1 vccd1 _11800_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09668__D line[125] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13538_ _13540_/CLK line[88] vssd1 vssd1 vccd1 vccd1 _13539_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10607__D line[42] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13469_ _13469_/A _13474_/Y vssd1 vssd1 vccd1 vccd1 _13749_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06092__D line[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06010_ _06010_/A _06019_/Y vssd1 vssd1 vccd1 vccd1 _13850_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_145_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12822__D line[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[8\].VALID\[13\].FF OVHB\[8\].V/CLK A[20] vssd1 vssd1 vccd1 vccd1 OVHB\[8\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XOVHB\[12\].VALID\[0\].FF OVHB\[12\].V/CLK A[7] vssd1 vssd1 vccd1 vccd1 OVHB\[12\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07916__D line[92] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06820__D line[89] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07961_ _07975_/CLK line[98] vssd1 vssd1 vccd1 vccd1 _07962_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11438__D line[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09700_ _09700_/A _09729_/Y vssd1 vssd1 vccd1 vccd1 _13620_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.M\[1\].MUX\[7\]_A2 _13768_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06912_ _06912_/A _06929_/Y vssd1 vssd1 vccd1 vccd1 _13632_/Z sky130_fd_sc_hd__ebufn_2
X_07892_ _07892_/A _07909_/Y vssd1 vssd1 vccd1 vccd1 _13772_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_95_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XOVHB\[21\].VALID\[4\].TOBUF OVHB\[21\].VALID\[4\].FF/Q OVHB\[21\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04925_/B2 sky130_fd_sc_hd__ebufn_2
X_09631_ _09655_/CLK line[108] vssd1 vssd1 vccd1 vccd1 _09632_/A sky130_fd_sc_hd__dfxtp_1
X_06843_ _06855_/CLK line[99] vssd1 vssd1 vccd1 vccd1 _06844_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_67_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09562_ _09562_/A _09589_/Y vssd1 vssd1 vccd1 vccd1 _13762_/Z sky130_fd_sc_hd__ebufn_2
X_06774_ _06774_/A _06789_/Y vssd1 vssd1 vccd1 vccd1 _13774_/Z sky130_fd_sc_hd__ebufn_2
X_08513_ _08535_/CLK line[109] vssd1 vssd1 vccd1 vccd1 _08514_/A sky130_fd_sc_hd__dfxtp_1
X_05725_ _05735_/CLK line[100] vssd1 vssd1 vccd1 vccd1 _05726_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_36_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09493_ _09515_/CLK line[45] vssd1 vssd1 vccd1 vccd1 _09494_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11173__D line[45] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08444_ _08444_/A _08469_/Y vssd1 vssd1 vccd1 vccd1 _13764_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06267__D line[106] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05656_ _05656_/A _05669_/Y vssd1 vssd1 vccd1 vccd1 _13776_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05171__D line[103] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08375_ _08395_/CLK line[46] vssd1 vssd1 vccd1 vccd1 _08376_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_149_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05587_ _05595_/CLK line[37] vssd1 vssd1 vccd1 vccd1 _05588_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_177_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07326_ _07326_/A _07349_/Y vssd1 vssd1 vccd1 vccd1 _13766_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08482__D line[95] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07257_ _07275_/CLK line[47] vssd1 vssd1 vccd1 vccd1 _07258_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07098__D line[88] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[18\].VALID\[3\].FF_D A[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06208_ _06208_/A _06229_/Y vssd1 vssd1 vccd1 vccd1 _13768_/Z sky130_fd_sc_hd__ebufn_2
X_07188_ _07188_/A _07209_/Y vssd1 vssd1 vccd1 vccd1 _13628_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_3_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11198__A _13933_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06139_ _06155_/CLK line[33] vssd1 vssd1 vccd1 vccd1 _06140_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_132_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[28\].VALID\[5\].FF OVHB\[28\].V/CLK A[12] vssd1 vssd1 vccd1 vccd1 OVHB\[28\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06730__D line[62] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11348__D line[125] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05346__D line[55] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09829_ _09829_/A _09834_/Y vssd1 vssd1 vccd1 vccd1 _13749_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_73_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13563__D line[99] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12840_ _12840_/CLK line[25] vssd1 vssd1 vccd1 vccd1 _12841_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_74_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08657__D line[47] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[10\].VALID\[2\].FF OVHB\[10\].V/CLK A[9] vssd1 vssd1 vccd1 vccd1 OVHB\[10\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_12771_ _12771_/A _12774_/Y vssd1 vssd1 vccd1 vccd1 _13891_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11722_ _11722_/CLK _11723_/X vssd1 vssd1 vccd1 vccd1 _11720_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_70_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05081__D line[76] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XOVHB\[17\].VALID\[10\].TOBUF OVHB\[17\].VALID\[10\].FF/Q OVHB\[17\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04932_/B2 sky130_fd_sc_hd__ebufn_2
XPHY_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11653_ _13926_/X wr vssd1 vssd1 vccd1 vccd1 _11653_/X sky130_fd_sc_hd__and2_1
XPHY_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11811__D line[66] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTIE vssd1 vssd1 vccd1 vccd1 TIE/HI TIE/LO sky130_fd_sc_hd__conb_1
X_10604_ _13924_/X vssd1 vssd1 vccd1 vccd1 _10604_/Y sky130_fd_sc_hd__inv_2
XPHY_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06905__D line[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11584_ _13926_/X vssd1 vssd1 vccd1 vccd1 _11584_/Y sky130_fd_sc_hd__inv_2
XPHY_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13323_ _13323_/A _13334_/Y vssd1 vssd1 vccd1 vccd1 _13883_/Z sky130_fd_sc_hd__ebufn_2
X_10535_ _10565_/CLK line[0] vssd1 vssd1 vccd1 vccd1 _10536_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_13_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__04924__A1_N A_h[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13254_ _13260_/CLK line[86] vssd1 vssd1 vccd1 vccd1 _13255_/A sky130_fd_sc_hd__dfxtp_1
X_10466_ _10466_/A _10499_/Y vssd1 vssd1 vccd1 vccd1 _13826_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13738__D line[51] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12205_ _12205_/A _12214_/Y vssd1 vssd1 vccd1 vccd1 _13885_/Z sky130_fd_sc_hd__ebufn_2
X_13185_ _13185_/A _13194_/Y vssd1 vssd1 vccd1 vccd1 _13745_/Z sky130_fd_sc_hd__ebufn_2
X_10397_ _10425_/CLK line[74] vssd1 vssd1 vccd1 vccd1 _10398_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_151_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12136_ _12140_/CLK line[87] vssd1 vssd1 vccd1 vccd1 _12137_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10162__D line[95] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12067_ _12067_/A _12074_/Y vssd1 vssd1 vccd1 vccd1 _13747_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05256__D line[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11018_ _11020_/CLK line[88] vssd1 vssd1 vccd1 vccd1 _11019_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_37_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[26\].VALID\[7\].FF OVHB\[26\].V/CLK A[14] vssd1 vssd1 vccd1 vccd1 OVHB\[26\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07471__D line[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12089__D line[65] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12969_ _12969_/A _12984_/Y vssd1 vssd1 vccd1 vccd1 _13809_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_18_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05510_ _05510_/A _05529_/Y vssd1 vssd1 vccd1 vccd1 _13630_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_61_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06490_ _06490_/A _06509_/Y vssd1 vssd1 vccd1 vccd1 _13770_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_205_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_OVHB\[9\].VALID\[12\].FF_D A[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05441_ _05455_/CLK line[98] vssd1 vssd1 vccd1 vccd1 _05442_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[16\].CLKBUF\[6\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09398__D line[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08160_ _08160_/A _08189_/Y vssd1 vssd1 vccd1 vccd1 _13760_/Z sky130_fd_sc_hd__ebufn_2
X_05372_ _05372_/A _05389_/Y vssd1 vssd1 vccd1 vccd1 _13772_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_159_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07111_ _07135_/CLK line[108] vssd1 vssd1 vccd1 vccd1 _07112_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10337__D line[47] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08091_ _08115_/CLK line[44] vssd1 vssd1 vccd1 vccd1 _08092_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_158_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07042_ _07042_/A _07069_/Y vssd1 vssd1 vccd1 vccd1 _13762_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__04913__A A_h[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12552__D line[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07646__D line[82] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08993_ _13915_/X wr vssd1 vssd1 vccd1 vccd1 _08993_/X sky130_fd_sc_hd__and2_1
XFILLER_125_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07944_ _13912_/X vssd1 vssd1 vccd1 vccd1 _07944_/Y sky130_fd_sc_hd__inv_2
XANTENNA__07943__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09861__D line[71] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[9\].CLKBUF\[6\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07875_ _07905_/CLK line[64] vssd1 vssd1 vccd1 vccd1 _07876_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_110_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13961__A A_h[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09614_ _09620_/CLK line[86] vssd1 vssd1 vccd1 vccd1 _09615_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10800__D line[116] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06826_ _06826_/A _06859_/Y vssd1 vssd1 vccd1 vccd1 _13826_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_141_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09545_ _09545_/A _09554_/Y vssd1 vssd1 vccd1 vccd1 _13745_/Z sky130_fd_sc_hd__ebufn_2
X_06757_ _06785_/CLK line[74] vssd1 vssd1 vccd1 vccd1 _06758_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_52_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05708_ _05708_/A _05739_/Y vssd1 vssd1 vccd1 vccd1 _13828_/Z sky130_fd_sc_hd__ebufn_2
X_09476_ _09480_/CLK line[23] vssd1 vssd1 vccd1 vccd1 _09477_/A sky130_fd_sc_hd__dfxtp_1
XPHY_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06688_ _06688_/A _06719_/Y vssd1 vssd1 vccd1 vccd1 _13688_/Z sky130_fd_sc_hd__ebufn_2
XPHY_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08427_ _08427_/A _08434_/Y vssd1 vssd1 vccd1 vccd1 _13747_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_169_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12727__D line[101] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05639_ _05665_/CLK line[75] vssd1 vssd1 vccd1 vccd1 _05640_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_24_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[24\].VALID\[9\].FF OVHB\[24\].V/CLK A[16] vssd1 vssd1 vccd1 vccd1 OVHB\[24\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08358_ _08360_/CLK line[24] vssd1 vssd1 vccd1 vccd1 _08359_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[4\].VALID\[11\].FF OVHB\[4\].V/CLK A[18] vssd1 vssd1 vccd1 vccd1 OVHB\[4\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07309_ _07309_/A _07314_/Y vssd1 vssd1 vccd1 vccd1 _13749_/Z sky130_fd_sc_hd__ebufn_2
X_08289_ _08289_/A _08294_/Y vssd1 vssd1 vccd1 vccd1 _13889_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_166_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10320_ _10320_/CLK line[25] vssd1 vssd1 vccd1 vccd1 _10321_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10251_ _10251_/A _10254_/Y vssd1 vssd1 vccd1 vccd1 _13891_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12462__D line[122] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06460__D line[52] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10182_ _10182_/CLK _10183_/X vssd1 vssd1 vccd1 vccd1 _10180_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_182_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11078__D line[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09771__D line[44] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13941_ A_h[2] vssd1 vssd1 vccd1 vccd1 _13949_/C sky130_fd_sc_hd__clkbuf_2
XOVHB\[3\].VALID\[1\].TOBUF OVHB\[3\].VALID\[1\].FF/Q OVHB\[3\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04926_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__13293__D line[104] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10710__D line[80] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08387__D line[37] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13872_ _13890_/CLK line[127] vssd1 vssd1 vccd1 vccd1 _13873_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[28\].VALID\[4\].TOBUF OVHB\[28\].VALID\[4\].FF/Q OVHB\[28\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04925_/B2 sky130_fd_sc_hd__ebufn_2
X_12823_ _12823_/A _12844_/Y vssd1 vssd1 vccd1 vccd1 _13663_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_15_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12754_ _12770_/CLK line[113] vssd1 vssd1 vccd1 vccd1 _12755_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[26\].VOBUF OVHB\[26\].V/Q OVHB\[26\].INV/Y vssd1 vssd1 vccd1 vccd1 _04912_/B1
+ sky130_fd_sc_hd__ebufn_2
X_11705_ _11705_/A _11724_/Y vssd1 vssd1 vccd1 vccd1 _13665_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12637__D line[74] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12685_ _12685_/A _12704_/Y vssd1 vssd1 vccd1 vccd1 _13805_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11541__D line[71] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11636_ _11650_/CLK line[114] vssd1 vssd1 vccd1 vccd1 _11637_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06635__D line[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09011__D line[66] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11567_ _11567_/A _11584_/Y vssd1 vssd1 vccd1 vccd1 _13807_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09946__D line[124] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13306_ _13330_/CLK line[124] vssd1 vssd1 vccd1 vccd1 _13307_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08850__D line[121] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10518_ _10530_/CLK line[115] vssd1 vssd1 vccd1 vccd1 _10519_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_6_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11498_ _11510_/CLK line[51] vssd1 vssd1 vccd1 vccd1 _11499_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_170_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13468__D line[56] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13237_ _13237_/A _13264_/Y vssd1 vssd1 vccd1 vccd1 _13797_/Z sky130_fd_sc_hd__ebufn_2
X_10449_ _10449_/A _10464_/Y vssd1 vssd1 vccd1 vccd1 _13809_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06370__D line[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13168_ _13190_/CLK line[61] vssd1 vssd1 vccd1 vccd1 _13169_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_123_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12119_ _12119_/A _12144_/Y vssd1 vssd1 vccd1 vccd1 _13799_/Z sky130_fd_sc_hd__ebufn_2
X_13099_ _13099_/A _13124_/Y vssd1 vssd1 vccd1 vccd1 _13659_/Z sky130_fd_sc_hd__ebufn_2
X_05990_ _05990_/A _06019_/Y vssd1 vssd1 vccd1 vccd1 _13830_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05564__A _13901_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_04941_ _04965_/CLK line[12] vssd1 vssd1 vccd1 vccd1 _04942_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11716__D line[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05283__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08297__D line[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07660_ _07660_/CLK line[89] vssd1 vssd1 vccd1 vccd1 _07661_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_92_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06611_ _06611_/A _06614_/Y vssd1 vssd1 vccd1 vccd1 _13891_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[21\].VALID\[2\].FF_D A[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07591_ _07591_/A _07594_/Y vssd1 vssd1 vccd1 vccd1 _13751_/Z sky130_fd_sc_hd__ebufn_2
X_09330_ _09340_/CLK line[84] vssd1 vssd1 vccd1 vccd1 _09331_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_206_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06542_ _06542_/CLK _06543_/X vssd1 vssd1 vccd1 vccd1 _06540_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_179_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09261_ _09261_/A _09274_/Y vssd1 vssd1 vccd1 vccd1 _13741_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[18\].VALID\[11\].FF OVHB\[18\].V/CLK A[18] vssd1 vssd1 vccd1 vccd1 OVHB\[18\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_06473_ _13904_/X wr vssd1 vssd1 vccd1 vccd1 _06473_/X sky130_fd_sc_hd__and2_1
XANTENNA__11451__D line[44] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08212_ _08220_/CLK line[85] vssd1 vssd1 vccd1 vccd1 _08213_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06545__D line[96] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05424_ _13900_/X vssd1 vssd1 vccd1 vccd1 _05424_/Y sky130_fd_sc_hd__inv_2
X_09192_ _09200_/CLK line[21] vssd1 vssd1 vccd1 vccd1 _09193_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[14\].VALID\[6\].FF_D A[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08143_ _08143_/A _08154_/Y vssd1 vssd1 vccd1 vccd1 _13743_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10067__D line[37] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05355_ _05385_/CLK line[64] vssd1 vssd1 vccd1 vccd1 _05356_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05739__A _13901_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08760__D line[94] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08074_ _08080_/CLK line[22] vssd1 vssd1 vccd1 vccd1 _08075_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_119_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05286_ _05286_/A _05319_/Y vssd1 vssd1 vccd1 vccd1 _13686_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_174_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13378__D line[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07025_ _07025_/A _07034_/Y vssd1 vssd1 vccd1 vccd1 _13745_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05458__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07376__D line[87] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08976_ _08990_/CLK line[50] vssd1 vssd1 vccd1 vccd1 _08977_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_29_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07927_ _07927_/A _07944_/Y vssd1 vssd1 vccd1 vccd1 _13807_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_69_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11626__D line[124] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[11\].VALID\[10\].FF_D A[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10530__D line[121] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07858_ _07870_/CLK line[51] vssd1 vssd1 vccd1 vccd1 _07859_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_28_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05624__D line[54] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08000__D line[116] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06809_ _06809_/A _06824_/Y vssd1 vssd1 vccd1 vccd1 _13809_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_43_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07789_ _07789_/A _07804_/Y vssd1 vssd1 vccd1 vccd1 _13669_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13841__D line[98] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08935__D line[46] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09528_ _09550_/CLK line[61] vssd1 vssd1 vccd1 vccd1 _09529_/A sky130_fd_sc_hd__dfxtp_1
XPHY_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09459_ _09459_/A _09484_/Y vssd1 vssd1 vccd1 vccd1 _13659_/Z sky130_fd_sc_hd__ebufn_2
XPHY_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12470_ _12490_/CLK line[126] vssd1 vssd1 vccd1 vccd1 _12471_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[30\].V_D TIE/HI vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11421_ _11421_/A _11444_/Y vssd1 vssd1 vccd1 vccd1 _13661_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_177_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XOVHB\[1\].VALID\[6\].TOBUF OVHB\[1\].VALID\[6\].FF/Q OVHB\[1\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04923_/A2 sky130_fd_sc_hd__ebufn_2
X_11352_ _11370_/CLK line[127] vssd1 vssd1 vccd1 vccd1 _11353_/A sky130_fd_sc_hd__dfxtp_1
X_10303_ _10303_/A _10324_/Y vssd1 vssd1 vccd1 vccd1 _13663_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12192__D line[127] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[26\].VALID\[9\].TOBUF OVHB\[26\].VALID\[9\].FF/Q OVHB\[26\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04914_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__10705__D line[73] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11283_ _11283_/A _11304_/Y vssd1 vssd1 vccd1 vccd1 _13803_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_106_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07286__D line[60] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06190__D line[57] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13022_ _13050_/CLK line[122] vssd1 vssd1 vccd1 vccd1 _13023_/A sky130_fd_sc_hd__dfxtp_1
X_10234_ _10250_/CLK line[113] vssd1 vssd1 vccd1 vccd1 _10235_/A sky130_fd_sc_hd__dfxtp_1
X_10165_ _10165_/A _10184_/Y vssd1 vssd1 vccd1 vccd1 _13805_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_86_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10096_ _10110_/CLK line[50] vssd1 vssd1 vccd1 vccd1 _10097_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10440__D line[94] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13924_ _13927_/A _13927_/B _13927_/C _13927_/D vssd1 vssd1 vccd1 vccd1 _13924_/X
+ sky130_fd_sc_hd__and4bb_4
XANTENNA__05534__D line[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13855_ _13855_/CLK line[105] vssd1 vssd1 vccd1 vccd1 _13856_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_16_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12806_ _12806_/A _12809_/Y vssd1 vssd1 vccd1 vccd1 _13646_/Z sky130_fd_sc_hd__ebufn_2
X_13786_ _13786_/A _13789_/Y vssd1 vssd1 vccd1 vccd1 _13786_/Z sky130_fd_sc_hd__ebufn_2
X_10998_ _11020_/CLK line[93] vssd1 vssd1 vccd1 vccd1 _10999_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07104__A _13909_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12367__D line[79] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[27\].VALID\[6\].FF_D A[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12737_ _12737_/CLK _12738_/X vssd1 vssd1 vccd1 vccd1 _12735_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__06365__D line[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12668_ _13936_/X wr vssd1 vssd1 vccd1 vccd1 _12668_/X sky130_fd_sc_hd__and2_1
XPHY_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11619_ _13926_/X vssd1 vssd1 vccd1 vccd1 _11619_/Y sky130_fd_sc_hd__inv_2
XANTENNA__09676__D line[114] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12599_ _13936_/X vssd1 vssd1 vccd1 vccd1 _12599_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05140_ _05140_/CLK line[89] vssd1 vssd1 vccd1 vccd1 _05141_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09973__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05071_ _05071_/A _05074_/Y vssd1 vssd1 vccd1 vccd1 _13751_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10615__D line[46] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[25\].CGAND_B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05709__D line[107] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12830__D line[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08830_ _08850_/CLK line[126] vssd1 vssd1 vccd1 vccd1 _08831_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[29\].CGAND_A _13925_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07924__D line[81] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08761_ _08761_/A _08784_/Y vssd1 vssd1 vccd1 vccd1 _13801_/Z sky130_fd_sc_hd__ebufn_2
X_05973_ _05973_/A _05984_/Y vssd1 vssd1 vccd1 vccd1 _13813_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_66_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07712_ _07730_/CLK line[127] vssd1 vssd1 vccd1 vccd1 _07713_/A sky130_fd_sc_hd__dfxtp_1
X_04924_ A_h[5] _04924_/B2 A_h[5] _04924_/B2 vssd1 vssd1 vccd1 vccd1 _04928_/A sky130_fd_sc_hd__a2bb2oi_2
XOVHB\[15\].CG clk OVHB\[15\].CGAND/X vssd1 vssd1 vccd1 vccd1 OVHB\[15\].V/CLK sky130_fd_sc_hd__dlclkp_1
X_08692_ _08710_/CLK line[63] vssd1 vssd1 vccd1 vccd1 _08693_/A sky130_fd_sc_hd__dfxtp_1
X_07643_ _07643_/A _07664_/Y vssd1 vssd1 vccd1 vccd1 _13803_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_25_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_MUX.M\[0\].MUX\[5\]_A3 _13848_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07574_ _07590_/CLK line[49] vssd1 vssd1 vccd1 vccd1 _07575_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_41_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[7\].VALID\[12\].TOBUF OVHB\[7\].VALID\[12\].FF/Q OVHB\[7\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04929_/B2 sky130_fd_sc_hd__ebufn_2
X_09313_ _09313_/A _09344_/Y vssd1 vssd1 vccd1 vccd1 _13793_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_81_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06525_ _06525_/A _06544_/Y vssd1 vssd1 vccd1 vccd1 _13805_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11181__D line[34] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09244_ _09270_/CLK line[59] vssd1 vssd1 vccd1 vccd1 _09245_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06275__D line[110] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06456_ _06470_/CLK line[50] vssd1 vssd1 vccd1 vccd1 _06457_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_166_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05407_ _05407_/A _05424_/Y vssd1 vssd1 vccd1 vccd1 _13807_/Z sky130_fd_sc_hd__ebufn_2
X_09175_ _09175_/A _09204_/Y vssd1 vssd1 vccd1 vccd1 _13655_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_21_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06387_ _06387_/A _06404_/Y vssd1 vssd1 vccd1 vccd1 _13667_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[28\].CLKBUF\[2\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08126_ _08150_/CLK line[60] vssd1 vssd1 vccd1 vccd1 _08127_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08490__D line[84] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05338_ _05350_/CLK line[51] vssd1 vssd1 vccd1 vccd1 _05339_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[16\].VALID\[14\].FF_D A[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08057_ _08057_/A _08084_/Y vssd1 vssd1 vccd1 vccd1 _13657_/Z sky130_fd_sc_hd__ebufn_2
X_05269_ _05269_/A _05284_/Y vssd1 vssd1 vccd1 vccd1 _13669_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[0\].V_D TIE/HI vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07008_ _07030_/CLK line[61] vssd1 vssd1 vccd1 vccd1 _07009_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[8\].VALID\[1\].FF_D A[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12740__D line[112] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[0\].VALID\[11\].TOBUF OVHB\[0\].VALID\[11\].FF/Q OVHB\[0\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04915_/B2 sky130_fd_sc_hd__ebufn_2
X_08959_ _13915_/X vssd1 vssd1 vccd1 vccd1 _08959_/Y sky130_fd_sc_hd__inv_2
XANTENNA_DEC.DEC0.AND2_A_N A[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11356__D line[114] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11934__A _13927_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11970_ _12000_/CLK line[16] vssd1 vssd1 vccd1 vccd1 _11971_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[26\].VALID\[13\].FF_D A[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10921_ _10921_/A _10954_/Y vssd1 vssd1 vccd1 vccd1 _13721_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11653__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13571__D line[103] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10852_ _10880_/CLK line[26] vssd1 vssd1 vccd1 vccd1 _10853_/A sky130_fd_sc_hd__dfxtp_1
X_13640_ _13640_/A _13649_/Y vssd1 vssd1 vccd1 vccd1 _13640_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08665__D line[36] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10783_ _10783_/A _10814_/Y vssd1 vssd1 vccd1 vccd1 _13863_/Z sky130_fd_sc_hd__ebufn_2
X_13571_ _13575_/CLK line[103] vssd1 vssd1 vccd1 vccd1 _13572_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_12_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12522_ _12522_/A _12529_/Y vssd1 vssd1 vccd1 vccd1 _13642_/Z sky130_fd_sc_hd__ebufn_2
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12915__D line[64] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12453_ _12455_/CLK line[104] vssd1 vssd1 vccd1 vccd1 _12454_/A sky130_fd_sc_hd__dfxtp_1
X_11404_ _11404_/A _11409_/Y vssd1 vssd1 vccd1 vccd1 _13644_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06913__D line[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12384_ _12384_/A _12389_/Y vssd1 vssd1 vccd1 vccd1 _13784_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_126_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11335_ _11335_/CLK line[105] vssd1 vssd1 vccd1 vccd1 _11336_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[1\].CLKBUF\[1\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07594__A _13911_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11266_ _11266_/A _11269_/Y vssd1 vssd1 vccd1 vccd1 _13786_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11828__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13746__D line[55] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13005_ _13015_/CLK line[100] vssd1 vssd1 vccd1 vccd1 _13006_/A sky130_fd_sc_hd__dfxtp_1
X_10217_ _10217_/CLK _10218_/X vssd1 vssd1 vccd1 vccd1 _10215_/CLK sky130_fd_sc_hd__dlclkp_1
X_11197_ _11197_/CLK _11198_/X vssd1 vssd1 vccd1 vccd1 _11195_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_95_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10148_ _13922_/X wr vssd1 vssd1 vccd1 vccd1 _10148_/X sky130_fd_sc_hd__and2_1
XANTENNA__10170__D line[84] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10079_ _13922_/X vssd1 vssd1 vccd1 vccd1 _10079_/Y sky130_fd_sc_hd__inv_2
XANTENNA__05264__D line[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13907_ A[3] vssd1 vssd1 vccd1 vccd1 _13916_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_47_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13481__D line[76] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[18\].VALID\[10\].FF_D A[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08575__D line[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13838_ _13838_/A _13859_/Y vssd1 vssd1 vccd1 vccd1 _13838_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12097__D line[69] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[10\].VALID\[9\].FF_D A[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13769_ _13785_/CLK line[65] vssd1 vssd1 vccd1 vccd1 _13770_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06310_ _06330_/CLK line[126] vssd1 vssd1 vccd1 vccd1 _06311_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07769__A _13912_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07290_ _07310_/CLK line[62] vssd1 vssd1 vccd1 vccd1 _07291_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_188_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06241_ _06241_/A _06264_/Y vssd1 vssd1 vccd1 vccd1 _13801_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07488__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06172_ _06190_/CLK line[63] vssd1 vssd1 vccd1 vccd1 _06173_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_156_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XDATA\[19\].CLKBUF\[5\] clk vssd1 vssd1 vccd1 vccd1 _07942_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_172_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05123_ _05123_/A _05144_/Y vssd1 vssd1 vccd1 vccd1 _13803_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_7_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10345__D line[36] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05439__D line[97] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[8\].VALID\[6\].TOBUF OVHB\[8\].VALID\[6\].FF/Q OVHB\[8\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04923_/A2 sky130_fd_sc_hd__ebufn_2
X_05054_ _05070_/CLK line[49] vssd1 vssd1 vccd1 vccd1 _05055_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_104_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09931_ _09935_/CLK line[103] vssd1 vssd1 vccd1 vccd1 _09932_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13656__D line[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12560__D line[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09862_ _09862_/A _09869_/Y vssd1 vssd1 vccd1 vccd1 _13782_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07654__D line[86] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08813_ _08815_/CLK line[104] vssd1 vssd1 vccd1 vccd1 _08814_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_112_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09793_ _09795_/CLK line[40] vssd1 vssd1 vccd1 vccd1 _09794_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_100_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10080__D line[48] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08744_ _08744_/A _08749_/Y vssd1 vssd1 vccd1 vccd1 _13784_/Z sky130_fd_sc_hd__ebufn_2
X_05956_ _05980_/CLK line[92] vssd1 vssd1 vccd1 vccd1 _05957_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_26_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08675_ _08675_/CLK line[41] vssd1 vssd1 vccd1 vccd1 _08676_/A sky130_fd_sc_hd__dfxtp_1
X_05887_ _05887_/A _05914_/Y vssd1 vssd1 vccd1 vccd1 _13727_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[23\].VALID\[13\].TOBUF OVHB\[23\].VALID\[13\].FF/Q OVHB\[23\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04916_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__11904__D line[123] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[9\].VALID\[11\].FF OVHB\[9\].V/CLK A[18] vssd1 vssd1 vccd1 vccd1 OVHB\[9\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_07626_ _07626_/A _07629_/Y vssd1 vssd1 vccd1 vccd1 _13786_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05902__D line[53] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07557_ _07557_/CLK _07558_/X vssd1 vssd1 vccd1 vccd1 _07555_/CLK sky130_fd_sc_hd__dlclkp_1
XPHY_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06508_ _13904_/X wr vssd1 vssd1 vccd1 vccd1 _06508_/X sky130_fd_sc_hd__and2_1
X_07488_ _13911_/X wr vssd1 vssd1 vccd1 vccd1 _07488_/X sky130_fd_sc_hd__and2_1
XFILLER_21_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12735__D line[105] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06439_ _13904_/X vssd1 vssd1 vccd1 vccd1 _06439_/Y sky130_fd_sc_hd__inv_2
X_09227_ _09235_/CLK line[37] vssd1 vssd1 vccd1 vccd1 _09228_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_6_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07829__D line[38] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09158_ _09158_/A _09169_/Y vssd1 vssd1 vccd1 vccd1 _13638_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_181_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08109_ _08115_/CLK line[38] vssd1 vssd1 vccd1 vccd1 _08110_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10255__D line[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09089_ _09095_/CLK line[102] vssd1 vssd1 vccd1 vccd1 _09090_/A sky130_fd_sc_hd__dfxtp_1
X_11120_ _11120_/A _11129_/Y vssd1 vssd1 vccd1 vccd1 _13640_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[26\].CLKBUF\[4\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12470__D line[126] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11051_ _11055_/CLK line[103] vssd1 vssd1 vccd1 vccd1 _11052_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[18\].CLKBUF\[2\] clk vssd1 vssd1 vccd1 vccd1 _07557_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_88_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07564__D line[59] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[30\].VALID\[5\].FF_D A[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10002_ _10002_/A _10009_/Y vssd1 vssd1 vccd1 vccd1 _13642_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_49_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11086__D line[119] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[8\].V_RESET_B rst_n vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[15\].VALID\[1\].TOBUF OVHB\[15\].VALID\[1\].FF/Q OVHB\[15\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04926_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__09134__A _13915_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11953_ _11965_/CLK line[3] vssd1 vssd1 vccd1 vccd1 _11954_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_205_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[23\].VALID\[9\].FF_D A[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08395__D line[41] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10904_ _10904_/A _10919_/Y vssd1 vssd1 vccd1 vccd1 _13704_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_205_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11884_ _11884_/A _11899_/Y vssd1 vssd1 vccd1 vccd1 _13844_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05812__D line[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13623_ _13645_/CLK line[13] vssd1 vssd1 vccd1 vccd1 _13624_/A sky130_fd_sc_hd__dfxtp_1
X_10835_ _10845_/CLK line[4] vssd1 vssd1 vccd1 vccd1 _10836_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_198_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13554_ _13554_/A _13579_/Y vssd1 vssd1 vccd1 vccd1 _13834_/Z sky130_fd_sc_hd__ebufn_2
X_10766_ _10766_/A _10779_/Y vssd1 vssd1 vccd1 vccd1 _13846_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_13_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12505_ _12525_/CLK line[14] vssd1 vssd1 vccd1 vccd1 _12506_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12645__D line[78] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10697_ _10705_/CLK line[69] vssd1 vssd1 vccd1 vccd1 _10698_/A sky130_fd_sc_hd__dfxtp_1
X_13485_ _13505_/CLK line[78] vssd1 vssd1 vccd1 vccd1 _13486_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_173_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07739__D line[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[20\].VALID\[0\].FF OVHB\[20\].V/CLK A[7] vssd1 vssd1 vccd1 vccd1 OVHB\[20\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_145_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06643__D line[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12436_ _12436_/A _12459_/Y vssd1 vssd1 vccd1 vccd1 _13836_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_126_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10743__A _13924_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12367_ _12385_/CLK line[79] vssd1 vssd1 vccd1 vccd1 _12368_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09954__D line[113] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09309__A _13916_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11318_ _11318_/A _11339_/Y vssd1 vssd1 vccd1 vccd1 _13838_/Z sky130_fd_sc_hd__ebufn_2
X_12298_ _12298_/A _12319_/Y vssd1 vssd1 vccd1 vccd1 _13698_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_113_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11249_ _11265_/CLK line[65] vssd1 vssd1 vccd1 vccd1 _11250_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09028__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05810_ _05840_/CLK line[16] vssd1 vssd1 vccd1 vccd1 _05811_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_95_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06790_ _06820_/CLK line[80] vssd1 vssd1 vccd1 vccd1 _06791_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_55_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05741_ _05741_/A _05774_/Y vssd1 vssd1 vccd1 vccd1 _13861_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_36_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08460_ _08460_/A _08469_/Y vssd1 vssd1 vccd1 vccd1 _13780_/Z sky130_fd_sc_hd__ebufn_2
X_05672_ _05700_/CLK line[90] vssd1 vssd1 vccd1 vccd1 _05673_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06818__D line[88] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07411_ _07415_/CLK line[103] vssd1 vssd1 vccd1 vccd1 _07412_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_211_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08391_ _08395_/CLK line[39] vssd1 vssd1 vccd1 vccd1 _08392_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_189_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10918__A _13925_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07342_ _07342_/A _07349_/Y vssd1 vssd1 vccd1 vccd1 _13782_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_149_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[19\].VALID\[1\].FF OVHB\[19\].V/CLK A[8] vssd1 vssd1 vccd1 vccd1 OVHB\[19\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_07273_ _07275_/CLK line[40] vssd1 vssd1 vccd1 vccd1 _07274_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[21\].VALID\[0\].TOBUF OVHB\[21\].VALID\[0\].FF/Q OVHB\[21\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04924_/B2 sky130_fd_sc_hd__ebufn_2
X_09012_ _09012_/A _09029_/Y vssd1 vssd1 vccd1 vccd1 _13772_/Z sky130_fd_sc_hd__ebufn_2
X_06224_ _06224_/A _06229_/Y vssd1 vssd1 vccd1 vccd1 _13784_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06553__D line[109] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[4\].VALID\[4\].FF_D A[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10075__D line[41] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06155_ _06155_/CLK line[41] vssd1 vssd1 vccd1 vccd1 _06156_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05169__D line[102] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05106_ _05106_/A _05109_/Y vssd1 vssd1 vccd1 vccd1 _13786_/Z sky130_fd_sc_hd__ebufn_2
X_06086_ _06086_/A _06089_/Y vssd1 vssd1 vccd1 vccd1 _13646_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_104_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13386__D line[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05037_ _05037_/CLK _05038_/X vssd1 vssd1 vccd1 vccd1 _05035_/CLK sky130_fd_sc_hd__dlclkp_1
X_09914_ _09914_/A _09939_/Y vssd1 vssd1 vccd1 vccd1 _13834_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_86_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13683__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09845_ _09865_/CLK line[78] vssd1 vssd1 vccd1 vccd1 _09846_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_86_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09776_ _09776_/A _09799_/Y vssd1 vssd1 vccd1 vccd1 _13696_/Z sky130_fd_sc_hd__ebufn_2
X_06988_ _06988_/A _06999_/Y vssd1 vssd1 vccd1 vccd1 _13708_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06578__A _13904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08727_ _08745_/CLK line[79] vssd1 vssd1 vccd1 vccd1 _08728_/A sky130_fd_sc_hd__dfxtp_1
X_05939_ _05945_/CLK line[70] vssd1 vssd1 vccd1 vccd1 _05940_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11634__D line[113] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06728__D line[61] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08658_ _08658_/A _08679_/Y vssd1 vssd1 vccd1 vccd1 _13698_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09104__D line[123] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07609_ _07625_/CLK line[65] vssd1 vssd1 vccd1 vccd1 _07610_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08589_ _08605_/CLK line[1] vssd1 vssd1 vccd1 vccd1 _08590_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08943__D line[35] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10620_ _10620_/A _10639_/Y vssd1 vssd1 vccd1 vccd1 _13700_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10551_ _10565_/CLK line[2] vssd1 vssd1 vccd1 vccd1 _10552_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_139_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10482_ _10482_/A _10499_/Y vssd1 vssd1 vccd1 vccd1 _13842_/Z sky130_fd_sc_hd__ebufn_2
X_13270_ _13270_/A _13299_/Y vssd1 vssd1 vccd1 vccd1 _13830_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_185_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13858__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12221_ _12245_/CLK line[12] vssd1 vssd1 vccd1 vccd1 _12222_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[13\].VALID\[6\].TOBUF OVHB\[13\].VALID\[6\].FF/Q OVHB\[13\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04923_/A2 sky130_fd_sc_hd__ebufn_2
XANTENNA__05079__D line[75] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12152_ _12152_/A _12179_/Y vssd1 vssd1 vccd1 vccd1 _13832_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_108_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XOVHB\[17\].VALID\[3\].FF OVHB\[17\].V/CLK A[10] vssd1 vssd1 vccd1 vccd1 OVHB\[17\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_11103_ _11125_/CLK line[13] vssd1 vssd1 vccd1 vccd1 _11104_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11809__D line[65] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12083_ _12105_/CLK line[77] vssd1 vssd1 vccd1 vccd1 _12084_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07294__D line[49] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11034_ _11034_/A _11059_/Y vssd1 vssd1 vccd1 vccd1 _13834_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_150_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_OVHB\[19\].VALID\[1\].FF_D A[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[4\].INV _13979_/X vssd1 vssd1 vccd1 vccd1 OVHB\[4\].INV/Y sky130_fd_sc_hd__inv_2
XANTENNA_DATA\[24\].CLKBUF\[6\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12985_ _13015_/CLK line[96] vssd1 vssd1 vccd1 vccd1 _12986_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DEC.DEC0.AND0_A A[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09799__A _13921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11936_ _11936_/A _11969_/Y vssd1 vssd1 vccd1 vccd1 _13616_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05542__D line[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11867_ _11895_/CLK line[106] vssd1 vssd1 vccd1 vccd1 _11868_/A sky130_fd_sc_hd__dfxtp_1
X_13606_ _13610_/CLK line[119] vssd1 vssd1 vccd1 vccd1 _13607_/A sky130_fd_sc_hd__dfxtp_1
X_10818_ _10818_/A _10849_/Y vssd1 vssd1 vccd1 vccd1 _13618_/Z sky130_fd_sc_hd__ebufn_2
X_11798_ _11798_/A _11829_/Y vssd1 vssd1 vccd1 vccd1 _13758_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12375__D line[68] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13537_ _13537_/A _13544_/Y vssd1 vssd1 vccd1 vccd1 _13817_/Z sky130_fd_sc_hd__ebufn_2
X_10749_ _10775_/CLK line[107] vssd1 vssd1 vccd1 vccd1 _10750_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07469__D line[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13468_ _13470_/CLK line[56] vssd1 vssd1 vccd1 vccd1 _13469_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_173_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12419_ _12419_/A _12424_/Y vssd1 vssd1 vccd1 vccd1 _13819_/Z sky130_fd_sc_hd__ebufn_2
X_13399_ _13399_/A _13404_/Y vssd1 vssd1 vccd1 vccd1 _13679_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09684__D line[118] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10623__D line[35] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07960_ _07960_/A _07979_/Y vssd1 vssd1 vccd1 vccd1 _13840_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_68_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05717__D line[111] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MUX.M\[1\].MUX\[7\]_A3 _13838_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06911_ _06925_/CLK line[2] vssd1 vssd1 vccd1 vccd1 _06912_/A sky130_fd_sc_hd__dfxtp_1
X_07891_ _07905_/CLK line[66] vssd1 vssd1 vccd1 vccd1 _07892_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_68_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09630_ _09630_/A _09659_/Y vssd1 vssd1 vccd1 vccd1 _13830_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_56_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06842_ _06842_/A _06859_/Y vssd1 vssd1 vccd1 vccd1 _13842_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_55_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07932__D line[85] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[15\].VALID\[5\].FF OVHB\[15\].V/CLK A[12] vssd1 vssd1 vccd1 vccd1 OVHB\[15\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_09561_ _09585_/CLK line[76] vssd1 vssd1 vccd1 vccd1 _09562_/A sky130_fd_sc_hd__dfxtp_1
X_06773_ _06785_/CLK line[67] vssd1 vssd1 vccd1 vccd1 _06774_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_209_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08512_ _08512_/A _08539_/Y vssd1 vssd1 vccd1 vccd1 _13832_/Z sky130_fd_sc_hd__ebufn_2
X_05724_ _05724_/A _05739_/Y vssd1 vssd1 vccd1 vccd1 _13844_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_24_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09492_ _09492_/A _09519_/Y vssd1 vssd1 vccd1 vccd1 _13692_/Z sky130_fd_sc_hd__ebufn_2
XPHY_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05655_ _05665_/CLK line[68] vssd1 vssd1 vccd1 vccd1 _05656_/A sky130_fd_sc_hd__dfxtp_1
X_08443_ _08465_/CLK line[77] vssd1 vssd1 vccd1 vccd1 _08444_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[31\].VALID\[14\].FF OVHB\[31\].V/CLK A[21] vssd1 vssd1 vccd1 vccd1 OVHB\[31\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_211_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09859__D line[70] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08374_ _08374_/A _08399_/Y vssd1 vssd1 vccd1 vccd1 _13694_/Z sky130_fd_sc_hd__ebufn_2
X_05586_ _05586_/A _05599_/Y vssd1 vssd1 vccd1 vccd1 _13706_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08118__A _13932_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07325_ _07345_/CLK line[78] vssd1 vssd1 vccd1 vccd1 _07326_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12285__D line[32] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07256_ _07256_/A _07279_/Y vssd1 vssd1 vccd1 vccd1 _13696_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_149_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06283__D line[99] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06207_ _06225_/CLK line[79] vssd1 vssd1 vccd1 vccd1 _06208_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11479__A _13926_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07187_ _07205_/CLK line[15] vssd1 vssd1 vccd1 vccd1 _07188_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09594__D line[91] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06138_ _06138_/A _06159_/Y vssd1 vssd1 vccd1 vccd1 _13698_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11198__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06069_ _06085_/CLK line[1] vssd1 vssd1 vccd1 vccd1 _06070_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_47_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09828_ _09830_/CLK line[56] vssd1 vssd1 vccd1 vccd1 _09829_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_171_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07842__D line[58] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XOVHB\[13\].VALID\[11\].TOBUF OVHB\[13\].VALID\[11\].FF/Q OVHB\[13\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04915_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_73_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09759_ _09759_/A _09764_/Y vssd1 vssd1 vccd1 vccd1 _13679_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_104_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11364__D line[118] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06458__D line[51] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12770_ _12770_/CLK line[121] vssd1 vssd1 vccd1 vccd1 _12771_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ _11721_/A _11724_/Y vssd1 vssd1 vccd1 vccd1 _13681_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09769__D line[43] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08673__D line[40] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[13\].VALID\[7\].FF OVHB\[13\].V/CLK A[14] vssd1 vssd1 vccd1 vccd1 OVHB\[13\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_11652_ _11652_/CLK _11653_/X vssd1 vssd1 vccd1 vccd1 _11650_/CLK sky130_fd_sc_hd__dlclkp_1
XPHY_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMUX.M\[0\].MUX\[0\] _13616_/Z _13686_/Z _13756_/Z _13826_/Z MUX.SEL0BUF\[0\]/X MUX.SEL1BUF\[0\]/X
+ vssd1 vssd1 vccd1 vccd1 Do[0] sky130_fd_sc_hd__mux4_1
XPHY_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10603_ _13924_/X wr vssd1 vssd1 vccd1 vccd1 _10603_/X sky130_fd_sc_hd__and2_1
XPHY_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11583_ _13926_/X wr vssd1 vssd1 vccd1 vccd1 _11583_/X sky130_fd_sc_hd__and2_1
XPHY_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12773__A _13936_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13322_ _13330_/CLK line[117] vssd1 vssd1 vccd1 vccd1 _13323_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_182_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10534_ _13923_/X vssd1 vssd1 vccd1 vccd1 _10534_/Y sky130_fd_sc_hd__inv_2
XPHY_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10465_ _10495_/CLK line[96] vssd1 vssd1 vccd1 vccd1 _10466_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[28\].VALID\[0\].TOBUF OVHB\[28\].VALID\[0\].FF/Q OVHB\[28\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04924_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__12923__D line[77] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13253_ _13253_/A _13264_/Y vssd1 vssd1 vccd1 vccd1 _13813_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_182_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12204_ _12210_/CLK line[118] vssd1 vssd1 vccd1 vccd1 _12205_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06921__D line[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13184_ _13190_/CLK line[54] vssd1 vssd1 vccd1 vccd1 _13185_/A sky130_fd_sc_hd__dfxtp_1
X_10396_ _10396_/A _10429_/Y vssd1 vssd1 vccd1 vccd1 _13756_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[9\].CLKBUF\[6\] clk vssd1 vssd1 vccd1 vccd1 _13857_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_151_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11539__D line[70] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12135_ _12135_/A _12144_/Y vssd1 vssd1 vccd1 vccd1 _13815_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[22\].VOBUF OVHB\[22\].V/Q OVHB\[22\].INV/Y vssd1 vssd1 vccd1 vccd1 _04912_/B1
+ sky130_fd_sc_hd__ebufn_2
XANTENNA__09009__D line[65] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12066_ _12070_/CLK line[55] vssd1 vssd1 vccd1 vccd1 _12067_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_77_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11017_ _11017_/A _11024_/Y vssd1 vssd1 vccd1 vccd1 _13817_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_38_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08848__D line[120] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11274__D line[91] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12948__A _13937_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05272__D line[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12968_ _12980_/CLK line[83] vssd1 vssd1 vccd1 vccd1 _12969_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_73_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11919_ _11919_/A _11934_/Y vssd1 vssd1 vccd1 vccd1 _13879_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_206_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12899_ _12899_/A _12914_/Y vssd1 vssd1 vccd1 vccd1 _13739_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_21_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05440_ _05440_/A _05459_/Y vssd1 vssd1 vccd1 vccd1 _13840_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_178_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08583__D line[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05371_ _05385_/CLK line[66] vssd1 vssd1 vccd1 vccd1 _05372_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[0\].VALID\[7\].FF_D A[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07199__D line[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07110_ _07110_/A _07139_/Y vssd1 vssd1 vccd1 vccd1 _13830_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_186_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08090_ _08090_/A _08119_/Y vssd1 vssd1 vccd1 vccd1 _13690_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_146_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07041_ _07065_/CLK line[76] vssd1 vssd1 vccd1 vccd1 _07042_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_146_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[11\].VALID\[9\].FF OVHB\[11\].V/CLK A[16] vssd1 vssd1 vccd1 vccd1 OVHB\[11\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_173_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06831__D line[108] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11449__D line[43] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10353__D line[40] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08992_ _08992_/CLK _08993_/X vssd1 vssd1 vccd1 vccd1 _08990_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__05447__D line[101] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07943_ _13912_/X wr vssd1 vssd1 vccd1 vccd1 _07943_/X sky130_fd_sc_hd__and2_1
XANTENNA__13664__D line[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDATA\[8\].CLKBUF\[3\] clk vssd1 vssd1 vccd1 vccd1 _13472_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__13019__A _13937_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08758__D line[93] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07874_ _13912_/X vssd1 vssd1 vccd1 vccd1 _07874_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09613_ _09613_/A _09624_/Y vssd1 vssd1 vccd1 vccd1 _13813_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_55_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06825_ _06855_/CLK line[96] vssd1 vssd1 vccd1 vccd1 _06826_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_83_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09544_ _09550_/CLK line[54] vssd1 vssd1 vccd1 vccd1 _09545_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_71_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06756_ _06756_/A _06789_/Y vssd1 vssd1 vccd1 vccd1 _13756_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05182__D line[122] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[3\].VALID\[13\].FF_D A[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05707_ _05735_/CLK line[106] vssd1 vssd1 vccd1 vccd1 _05708_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_197_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09475_ _09475_/A _09484_/Y vssd1 vssd1 vccd1 vccd1 _13675_/Z sky130_fd_sc_hd__ebufn_2
X_06687_ _06715_/CLK line[42] vssd1 vssd1 vccd1 vccd1 _06688_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11912__D line[127] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08426_ _08430_/CLK line[55] vssd1 vssd1 vccd1 vccd1 _08427_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_211_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05638_ _05638_/A _05669_/Y vssd1 vssd1 vccd1 vccd1 _13758_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05910__D line[57] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10528__D line[120] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08357_ _08357_/A _08364_/Y vssd1 vssd1 vccd1 vccd1 _13677_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05569_ _05595_/CLK line[43] vssd1 vssd1 vccd1 vccd1 _05570_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_20_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07308_ _07310_/CLK line[56] vssd1 vssd1 vccd1 vccd1 _07309_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_109_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_OVHB\[22\].VALID\[0\].FF_D A[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08288_ _08290_/CLK line[120] vssd1 vssd1 vccd1 vccd1 _08289_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13839__D line[97] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07239_ _07239_/A _07244_/Y vssd1 vssd1 vccd1 vccd1 _13679_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_152_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10250_ _10250_/CLK line[121] vssd1 vssd1 vccd1 vccd1 _10251_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[28\].CLKBUF\[7\] clk vssd1 vssd1 vccd1 vccd1 _10812_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_133_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10263__D line[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10181_ _10181_/A _10184_/Y vssd1 vssd1 vccd1 vccd1 _13821_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05357__D line[74] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[15\].VALID\[4\].FF_D A[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13940_ A_h[1] vssd1 vssd1 vccd1 vccd1 _13949_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_19_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07572__D line[63] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[1\].VALID\[2\].TOBUF OVHB\[1\].VALID\[2\].FF/Q OVHB\[1\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04930_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_46_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13871_ _13871_/A _13894_/Y vssd1 vssd1 vccd1 vccd1 _13871_/Z sky130_fd_sc_hd__ebufn_2
X_12822_ _12840_/CLK line[31] vssd1 vssd1 vccd1 vccd1 _12823_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06188__D line[56] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XDATA\[7\].CLKBUF\[0\] clk vssd1 vssd1 vccd1 vccd1 _13087_/CLK sky130_fd_sc_hd__clkbuf_4
XOVHB\[26\].VALID\[5\].TOBUF OVHB\[26\].VALID\[5\].FF/Q OVHB\[26\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04927_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_43_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12753_ _12753_/A _12774_/Y vssd1 vssd1 vccd1 vccd1 _13873_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10288__A _13923_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09499__D line[33] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11704_ _11720_/CLK line[17] vssd1 vssd1 vccd1 vccd1 _11705_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12684_ _12700_/CLK line[81] vssd1 vssd1 vccd1 vccd1 _12685_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_30_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05820__D line[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11635_ _11635_/A _11654_/Y vssd1 vssd1 vccd1 vccd1 _13875_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10438__D line[93] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[6\].VALID\[0\].FF OVHB\[6\].V/CLK A[7] vssd1 vssd1 vccd1 vccd1 OVHB\[6\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_DATA\[17\].CLKBUF\[0\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11566_ _11580_/CLK line[82] vssd1 vssd1 vccd1 vccd1 _11567_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13305_ _13305_/A _13334_/Y vssd1 vssd1 vccd1 vccd1 _13865_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12653__D line[67] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10517_ _10517_/A _10534_/Y vssd1 vssd1 vccd1 vccd1 _13877_/Z sky130_fd_sc_hd__ebufn_2
X_11497_ _11497_/A _11514_/Y vssd1 vssd1 vccd1 vccd1 _13737_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07747__D line[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13236_ _13260_/CLK line[92] vssd1 vssd1 vccd1 vccd1 _13237_/A sky130_fd_sc_hd__dfxtp_1
X_10448_ _10460_/CLK line[83] vssd1 vssd1 vccd1 vccd1 _10449_/A sky130_fd_sc_hd__dfxtp_1
X_13167_ _13167_/A _13194_/Y vssd1 vssd1 vccd1 vccd1 _13727_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_97_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10379_ _10379_/A _10394_/Y vssd1 vssd1 vccd1 vccd1 _13739_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09962__D line[117] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12118_ _12140_/CLK line[93] vssd1 vssd1 vccd1 vccd1 _12119_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[29\].CGAND _13925_/X wr vssd1 vssd1 vccd1 vccd1 OVHB\[29\].CGAND/X sky130_fd_sc_hd__and2_4
X_13098_ _13120_/CLK line[29] vssd1 vssd1 vccd1 vccd1 _13099_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[27\].CLKBUF\[4\] clk vssd1 vssd1 vccd1 vccd1 _10427_/CLK sky130_fd_sc_hd__clkbuf_4
XMUX.M\[3\].MUX\[5\] _13659_/Z _13729_/Z _13799_/Z _13869_/Z MUX.SEL0BUF\[3\]/X MUX.SEL1BUF\[3\]/X
+ vssd1 vssd1 vccd1 vccd1 Do[29] sky130_fd_sc_hd__mux4_1
X_04940_ _04940_/A _04969_/Y vssd1 vssd1 vccd1 vccd1 _13620_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10901__D line[34] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12049_ _12049_/A _12074_/Y vssd1 vssd1 vccd1 vccd1 _13729_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_38_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06098__D line[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06610_ _06610_/CLK line[121] vssd1 vssd1 vccd1 vccd1 _06611_/A sky130_fd_sc_hd__dfxtp_1
X_07590_ _07590_/CLK line[57] vssd1 vssd1 vccd1 vccd1 _07591_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_80_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06541_ _06541_/A _06544_/Y vssd1 vssd1 vccd1 vccd1 _13821_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12828__D line[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06472_ _06472_/CLK _06473_/X vssd1 vssd1 vccd1 vccd1 _06470_/CLK sky130_fd_sc_hd__dlclkp_1
X_09260_ _09270_/CLK line[52] vssd1 vssd1 vccd1 vccd1 _09261_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_61_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05423_ _13900_/X wr vssd1 vssd1 vccd1 vccd1 _05423_/X sky130_fd_sc_hd__and2_1
X_08211_ _08211_/A _08224_/Y vssd1 vssd1 vccd1 vccd1 _13811_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_194_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09191_ _09191_/A _09204_/Y vssd1 vssd1 vccd1 vccd1 _13671_/Z sky130_fd_sc_hd__ebufn_2
X_05354_ _13900_/X vssd1 vssd1 vccd1 vccd1 _05354_/Y sky130_fd_sc_hd__inv_2
X_08142_ _08150_/CLK line[53] vssd1 vssd1 vccd1 vccd1 _08143_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_146_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08073_ _08073_/A _08084_/Y vssd1 vssd1 vccd1 vccd1 _13673_/Z sky130_fd_sc_hd__ebufn_2
X_05285_ _05315_/CLK line[32] vssd1 vssd1 vccd1 vccd1 _05286_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_161_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07024_ _07030_/CLK line[54] vssd1 vssd1 vccd1 vccd1 _07025_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06561__D line[98] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_OVHB\[28\].VALID\[4\].FF_D A[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11179__D line[33] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[4\].VALID\[2\].FF OVHB\[4\].V/CLK A[9] vssd1 vssd1 vccd1 vccd1 OVHB\[4\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09872__D line[90] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08975_ _08975_/A _08994_/Y vssd1 vssd1 vccd1 vccd1 _13735_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_76_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13394__D line[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13972__A A_h[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08488__D line[83] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07926_ _07940_/CLK line[82] vssd1 vssd1 vccd1 vccd1 _07927_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_28_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07857_ _07857_/A _07874_/Y vssd1 vssd1 vccd1 vccd1 _13737_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_29_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XDATA\[26\].CLKBUF\[1\] clk vssd1 vssd1 vccd1 vccd1 _10042_/CLK sky130_fd_sc_hd__clkbuf_4
X_06808_ _06820_/CLK line[83] vssd1 vssd1 vccd1 vccd1 _06809_/A sky130_fd_sc_hd__dfxtp_1
X_07788_ _07800_/CLK line[19] vssd1 vssd1 vccd1 vccd1 _07789_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_45_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09527_ _09527_/A _09554_/Y vssd1 vssd1 vccd1 vccd1 _13727_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__04931__B1 A_h[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06739_ _06739_/A _06754_/Y vssd1 vssd1 vccd1 vccd1 _13739_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11642__D line[117] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDATA\[16\].CLKBUF\[7\] clk vssd1 vssd1 vccd1 vccd1 _07172_/CLK sky130_fd_sc_hd__clkbuf_4
XPHY_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06736__D line[50] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09458_ _09480_/CLK line[29] vssd1 vssd1 vccd1 vccd1 _09459_/A sky130_fd_sc_hd__dfxtp_1
XPHY_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09112__D line[127] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08409_ _08409_/A _08434_/Y vssd1 vssd1 vccd1 vccd1 _13729_/Z sky130_fd_sc_hd__ebufn_2
XMUX.M\[2\].MUX\[7\] _13677_/Z _13747_/Z _13817_/Z _13887_/Z MUX.SEL0BUF\[2\]/X MUX.SEL1BUF\[2\]/X
+ vssd1 vssd1 vccd1 vccd1 Do[23] sky130_fd_sc_hd__mux4_1
X_09389_ _09389_/A _09414_/Y vssd1 vssd1 vccd1 vccd1 _13869_/Z sky130_fd_sc_hd__ebufn_2
X_11420_ _11440_/CLK line[30] vssd1 vssd1 vccd1 vccd1 _11421_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_137_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08951__D line[39] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13569__D line[102] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11351_ _11351_/A _11374_/Y vssd1 vssd1 vccd1 vccd1 _13871_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_153_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10302_ _10320_/CLK line[31] vssd1 vssd1 vccd1 vccd1 _10303_/A sky130_fd_sc_hd__dfxtp_1
X_11282_ _11300_/CLK line[95] vssd1 vssd1 vccd1 vccd1 _11283_/A sky130_fd_sc_hd__dfxtp_1
X_13021_ _13021_/A _13054_/Y vssd1 vssd1 vccd1 vccd1 _13861_/Z sky130_fd_sc_hd__ebufn_2
X_10233_ _10233_/A _10254_/Y vssd1 vssd1 vccd1 vccd1 _13873_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05087__D line[79] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XOVHB\[30\].CGAND _13926_/X wr vssd1 vssd1 vccd1 vccd1 OVHB\[30\].CGAND/X sky130_fd_sc_hd__and2_4
X_10164_ _10180_/CLK line[81] vssd1 vssd1 vccd1 vccd1 _10165_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_79_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11817__D line[69] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10095_ _10095_/A _10114_/Y vssd1 vssd1 vccd1 vccd1 _13735_/Z sky130_fd_sc_hd__ebufn_2
X_13923_ _13927_/C _13927_/B _13927_/A _13927_/D vssd1 vssd1 vccd1 vccd1 _13923_/X
+ sky130_fd_sc_hd__and4b_4
XOVHB\[2\].VALID\[4\].FF OVHB\[2\].V/CLK A[11] vssd1 vssd1 vccd1 vccd1 OVHB\[2\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13854_ _13854_/A _13859_/Y vssd1 vssd1 vccd1 vccd1 _13854_/Z sky130_fd_sc_hd__ebufn_2
X_12805_ _12805_/CLK line[9] vssd1 vssd1 vccd1 vccd1 _12806_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_188_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13785_ _13785_/CLK line[73] vssd1 vssd1 vccd1 vccd1 _13786_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11552__D line[90] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10997_ _10997_/A _11024_/Y vssd1 vssd1 vccd1 vccd1 _13797_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_203_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12736_ _12736_/A _12739_/Y vssd1 vssd1 vccd1 vccd1 _13856_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05550__D line[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10168__D line[83] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12667_ _12667_/CLK _12668_/X vssd1 vssd1 vccd1 vccd1 _12665_/CLK sky130_fd_sc_hd__dlclkp_1
XPHY_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08861__D line[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDATA\[15\].CLKBUF\[4\] clk vssd1 vssd1 vccd1 vccd1 _06787_/CLK sky130_fd_sc_hd__clkbuf_4
X_11618_ _13926_/X wr vssd1 vssd1 vccd1 vccd1 _11618_/X sky130_fd_sc_hd__and2_1
XPHY_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12598_ _13936_/X wr vssd1 vssd1 vccd1 vccd1 _12598_/X sky130_fd_sc_hd__and2_1
XANTENNA__13479__D line[75] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12383__D line[72] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11549_ _13926_/X vssd1 vssd1 vccd1 vccd1 _11549_/Y sky130_fd_sc_hd__inv_2
XFILLER_144_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07477__D line[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05070_ _05070_/CLK line[57] vssd1 vssd1 vccd1 vccd1 _05071_/A sky130_fd_sc_hd__dfxtp_1
X_13219_ _13225_/CLK line[70] vssd1 vssd1 vccd1 vccd1 _13220_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[15\].CLKBUF\[2\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[29\].CGAND_B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11727__D line[42] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10631__D line[39] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08760_ _08780_/CLK line[94] vssd1 vssd1 vccd1 vccd1 _08761_/A sky130_fd_sc_hd__dfxtp_1
X_05972_ _05980_/CLK line[85] vssd1 vssd1 vccd1 vccd1 _05973_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[3\].VALID\[13\].TOBUF OVHB\[3\].VALID\[13\].FF/Q OVHB\[3\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04916_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__05725__D line[100] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08101__D line[34] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07711_ _07711_/A _07734_/Y vssd1 vssd1 vccd1 vccd1 _13871_/Z sky130_fd_sc_hd__ebufn_2
X_04923_ _04918_/Y _04923_/A2 _04919_/X _04921_/Y _04922_/X vssd1 vssd1 vccd1 vccd1
+ _04934_/B sky130_fd_sc_hd__o2111ai_2
X_08691_ _08691_/A _08714_/Y vssd1 vssd1 vccd1 vccd1 _13731_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[30\].VALID\[9\].TOBUF OVHB\[30\].VALID\[9\].FF/Q OVHB\[30\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04914_/B2 sky130_fd_sc_hd__ebufn_2
X_07642_ _07660_/CLK line[95] vssd1 vssd1 vccd1 vccd1 _07643_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_202_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07940__D line[89] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[14\].CG_CLK clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12558__D line[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[8\].VALID\[2\].TOBUF OVHB\[8\].VALID\[2\].FF/Q OVHB\[8\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04930_/B2 sky130_fd_sc_hd__ebufn_2
X_07573_ _07573_/A _07594_/Y vssd1 vssd1 vccd1 vccd1 _13733_/Z sky130_fd_sc_hd__ebufn_2
X_09312_ _09340_/CLK line[90] vssd1 vssd1 vccd1 vccd1 _09313_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_15_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06524_ _06540_/CLK line[81] vssd1 vssd1 vccd1 vccd1 _06525_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_80_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XOVHB\[0\].VALID\[6\].FF OVHB\[0\].V/CLK A[13] vssd1 vssd1 vccd1 vccd1 OVHB\[0\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[8\].CLKBUF\[2\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05460__D line[112] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09243_ _09243_/A _09274_/Y vssd1 vssd1 vccd1 vccd1 _13723_/Z sky130_fd_sc_hd__ebufn_2
X_06455_ _06455_/A _06474_/Y vssd1 vssd1 vccd1 vccd1 _13735_/Z sky130_fd_sc_hd__ebufn_2
X_05406_ _05420_/CLK line[82] vssd1 vssd1 vccd1 vccd1 _05407_/A sky130_fd_sc_hd__dfxtp_1
X_09174_ _09200_/CLK line[27] vssd1 vssd1 vccd1 vccd1 _09175_/A sky130_fd_sc_hd__dfxtp_1
X_06386_ _06400_/CLK line[18] vssd1 vssd1 vccd1 vccd1 _06387_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_182_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05337_ _05337_/A _05354_/Y vssd1 vssd1 vccd1 vccd1 _13737_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12293__D line[45] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08125_ _08125_/A _08154_/Y vssd1 vssd1 vccd1 vccd1 _13725_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10806__D line[119] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07387__D line[106] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06291__D line[103] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08056_ _08080_/CLK line[28] vssd1 vssd1 vccd1 vccd1 _08057_/A sky130_fd_sc_hd__dfxtp_1
X_05268_ _05280_/CLK line[19] vssd1 vssd1 vccd1 vccd1 _05269_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[11\].VALID\[7\].FF_D A[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDATA\[14\].CLKBUF\[1\] clk vssd1 vssd1 vccd1 vccd1 _06402_/CLK sky130_fd_sc_hd__clkbuf_4
X_07007_ _07007_/A _07034_/Y vssd1 vssd1 vccd1 vccd1 _13727_/Z sky130_fd_sc_hd__ebufn_2
X_05199_ _05199_/A _05214_/Y vssd1 vssd1 vccd1 vccd1 _13879_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_0_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10541__D line[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[7\].V_RESET_B rst_n vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08958_ _13915_/X wr vssd1 vssd1 vccd1 vccd1 _08958_/X sky130_fd_sc_hd__and2_1
XANTENNA__05635__D line[64] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07909_ _13912_/X vssd1 vssd1 vccd1 vccd1 _07909_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08889_ _13915_/X vssd1 vssd1 vccd1 vccd1 _08889_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10920_ _10950_/CLK line[48] vssd1 vssd1 vccd1 vccd1 _10921_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07850__D line[62] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10851_ _10851_/A _10884_/Y vssd1 vssd1 vccd1 vccd1 _13651_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12468__D line[125] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06466__D line[55] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13570_ _13570_/A _13579_/Y vssd1 vssd1 vccd1 vccd1 _13850_/Z sky130_fd_sc_hd__ebufn_2
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10782_ _10810_/CLK line[122] vssd1 vssd1 vccd1 vccd1 _10783_/A sky130_fd_sc_hd__dfxtp_1
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12521_ _12525_/CLK line[7] vssd1 vssd1 vccd1 vccd1 _12522_/A sky130_fd_sc_hd__dfxtp_1
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09777__D line[47] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12452_ _12452_/A _12459_/Y vssd1 vssd1 vccd1 vccd1 _13852_/Z sky130_fd_sc_hd__ebufn_2
X_11403_ _11405_/CLK line[8] vssd1 vssd1 vccd1 vccd1 _11404_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10716__D line[92] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12383_ _12385_/CLK line[72] vssd1 vssd1 vccd1 vccd1 _12384_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09039__TE_B _09064_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11334_ _11334_/A _11339_/Y vssd1 vssd1 vccd1 vccd1 _13854_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_21_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12931__D line[66] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11265_ _11265_/CLK line[73] vssd1 vssd1 vccd1 vccd1 _11266_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_180_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13004_ _13004_/A _13019_/Y vssd1 vssd1 vccd1 vccd1 _13844_/Z sky130_fd_sc_hd__ebufn_2
X_10216_ _10216_/A _10219_/Y vssd1 vssd1 vccd1 vccd1 _13856_/Z sky130_fd_sc_hd__ebufn_2
X_11196_ _11196_/A _11199_/Y vssd1 vssd1 vccd1 vccd1 _13716_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_97_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10147_ _10147_/CLK _10148_/X vssd1 vssd1 vccd1 vccd1 _10145_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_0_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09017__D line[69] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[20\].VALID\[14\].FF_D A[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10078_ _13922_/X wr vssd1 vssd1 vccd1 vccd1 _10078_/X sky130_fd_sc_hd__and2_1
XFILLER_63_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13906_ A[2] vssd1 vssd1 vccd1 vccd1 _13916_/A sky130_fd_sc_hd__clkbuf_2
XOVHB\[27\].VALID\[1\].FF OVHB\[27\].V/CLK A[8] vssd1 vssd1 vccd1 vccd1 OVHB\[27\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_13837_ _13855_/CLK line[111] vssd1 vssd1 vccd1 vccd1 _13838_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11282__D line[95] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_OVHB\[31\].VALID\[3\].FF_D A[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06376__D line[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05280__D line[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13768_ _13768_/A _13789_/Y vssd1 vssd1 vccd1 vccd1 _13768_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_204_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12719_ _12735_/CLK line[97] vssd1 vssd1 vccd1 vccd1 _12720_/A sky130_fd_sc_hd__dfxtp_1
X_13699_ _13715_/CLK line[33] vssd1 vssd1 vccd1 vccd1 _13700_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06240_ _06260_/CLK line[94] vssd1 vssd1 vccd1 vccd1 _06241_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08591__D line[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_OVHB\[30\].VALID\[13\].FF_D A[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_OVHB\[24\].VALID\[7\].FF_D A[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06171_ _06171_/A _06194_/Y vssd1 vssd1 vccd1 vccd1 _13731_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05122_ _05140_/CLK line[95] vssd1 vssd1 vccd1 vccd1 _05123_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_117_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07000__D line[48] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05053_ _05053_/A _05074_/Y vssd1 vssd1 vccd1 vccd1 _13733_/Z sky130_fd_sc_hd__ebufn_2
X_09930_ _09930_/A _09939_/Y vssd1 vssd1 vccd1 vccd1 _13850_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[6\].VALID\[7\].TOBUF OVHB\[6\].VALID\[7\].FF/Q OVHB\[6\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/A2 sky130_fd_sc_hd__ebufn_2
XFILLER_131_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09861_ _09865_/CLK line[71] vssd1 vssd1 vccd1 vccd1 _09862_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11457__D line[47] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08812_ _08812_/A _08819_/Y vssd1 vssd1 vccd1 vccd1 _13852_/Z sky130_fd_sc_hd__ebufn_2
X_09792_ _09792_/A _09799_/Y vssd1 vssd1 vccd1 vccd1 _13712_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05455__D line[105] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08743_ _08745_/CLK line[72] vssd1 vssd1 vccd1 vccd1 _08744_/A sky130_fd_sc_hd__dfxtp_1
X_05955_ _05955_/A _05984_/Y vssd1 vssd1 vccd1 vccd1 _13795_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13672__D line[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[13\].CLKBUF\[4\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08766__D line[82] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08674_ _08674_/A _08679_/Y vssd1 vssd1 vccd1 vccd1 _13714_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05886_ _05910_/CLK line[60] vssd1 vssd1 vccd1 vccd1 _05887_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[12\].VALID\[11\].FF_D A[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07625_ _07625_/CLK line[73] vssd1 vssd1 vccd1 vccd1 _07626_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_14_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07556_ _07556_/A _07559_/Y vssd1 vssd1 vccd1 vccd1 _13716_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05190__D line[126] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06507_ _06507_/CLK _06508_/X vssd1 vssd1 vccd1 vccd1 _06505_/CLK sky130_fd_sc_hd__dlclkp_1
X_07487_ _07487_/CLK _07488_/X vssd1 vssd1 vccd1 vccd1 _07485_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__11920__D line[116] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09226_ _09226_/A _09239_/Y vssd1 vssd1 vccd1 vccd1 _13706_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[25\].VALID\[3\].FF OVHB\[25\].V/CLK A[10] vssd1 vssd1 vccd1 vccd1 OVHB\[25\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_06438_ _13904_/X wr vssd1 vssd1 vccd1 vccd1 _06438_/X sky130_fd_sc_hd__and2_1
XFILLER_194_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09157_ _09165_/CLK line[5] vssd1 vssd1 vccd1 vccd1 _09158_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_181_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06369_ _13904_/X vssd1 vssd1 vccd1 vccd1 _06369_/Y sky130_fd_sc_hd__inv_2
XFILLER_107_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_OVHB\[22\].VALID\[10\].FF_D A[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08108_ _08108_/A _08119_/Y vssd1 vssd1 vccd1 vccd1 _13708_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[6\].CLKBUF\[4\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08006__D line[119] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09088_ _09088_/A _09099_/Y vssd1 vssd1 vccd1 vccd1 _13848_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13847__D line[101] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08039_ _08045_/CLK line[6] vssd1 vssd1 vccd1 vccd1 _08040_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_150_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11050_ _11050_/A _11059_/Y vssd1 vssd1 vccd1 vccd1 _13850_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10271__D line[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10001_ _10005_/CLK line[7] vssd1 vssd1 vccd1 vccd1 _10002_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_191_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05365__D line[78] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[5\].VALID\[2\].FF_D A[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_OVHB\[11\].CGAND_A _13901_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13582__D line[122] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11952_ _11952_/A _11969_/Y vssd1 vssd1 vccd1 vccd1 _13632_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07580__D line[52] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[13\].VALID\[2\].TOBUF OVHB\[13\].VALID\[2\].FF/Q OVHB\[13\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04930_/B2 sky130_fd_sc_hd__ebufn_2
X_10903_ _10915_/CLK line[35] vssd1 vssd1 vccd1 vccd1 _10904_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12198__D line[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11883_ _11895_/CLK line[99] vssd1 vssd1 vccd1 vccd1 _11884_/A sky130_fd_sc_hd__dfxtp_1
X_13622_ _13622_/A _13649_/Y vssd1 vssd1 vccd1 vccd1 _13622_/Z sky130_fd_sc_hd__ebufn_2
X_10834_ _10834_/A _10849_/Y vssd1 vssd1 vccd1 vccd1 _13634_/Z sky130_fd_sc_hd__ebufn_2
X_13553_ _13575_/CLK line[109] vssd1 vssd1 vccd1 vccd1 _13554_/A sky130_fd_sc_hd__dfxtp_1
X_10765_ _10775_/CLK line[100] vssd1 vssd1 vccd1 vccd1 _10766_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[22\].VALID\[14\].FF OVHB\[22\].V/CLK A[21] vssd1 vssd1 vccd1 vccd1 OVHB\[22\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11830__D line[80] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12504_ _12504_/A _12529_/Y vssd1 vssd1 vccd1 vccd1 _13624_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_8_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13484_ _13484_/A _13509_/Y vssd1 vssd1 vccd1 vccd1 _13764_/Z sky130_fd_sc_hd__ebufn_2
X_10696_ _10696_/A _10709_/Y vssd1 vssd1 vccd1 vccd1 _13776_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_8_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12435_ _12455_/CLK line[110] vssd1 vssd1 vccd1 vccd1 _12436_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10446__D line[82] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12366_ _12366_/A _12389_/Y vssd1 vssd1 vccd1 vccd1 _13766_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13757__D line[74] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10743__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12661__D line[71] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11317_ _11335_/CLK line[111] vssd1 vssd1 vccd1 vccd1 _11318_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_181_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12297_ _12315_/CLK line[47] vssd1 vssd1 vccd1 vccd1 _12298_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07755__D line[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[23\].VALID\[5\].FF OVHB\[23\].V/CLK A[12] vssd1 vssd1 vccd1 vccd1 OVHB\[23\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_11248_ _11248_/A _11269_/Y vssd1 vssd1 vccd1 vccd1 _13768_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_141_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11179_ _11195_/CLK line[33] vssd1 vssd1 vccd1 vccd1 _11180_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09970__D line[121] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05740_ _05770_/CLK line[112] vssd1 vssd1 vccd1 vccd1 _05741_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07490__D line[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05671_ _05671_/A _05704_/Y vssd1 vssd1 vccd1 vccd1 _13791_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_35_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07410_ _07410_/A _07419_/Y vssd1 vssd1 vccd1 vccd1 _13850_/Z sky130_fd_sc_hd__ebufn_2
X_08390_ _08390_/A _08399_/Y vssd1 vssd1 vccd1 vccd1 _13710_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_211_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06684__A _13905_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10918__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07341_ _07345_/CLK line[71] vssd1 vssd1 vccd1 vccd1 _07342_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[17\].VOBUF OVHB\[17\].V/Q OVHB\[17\].INV/Y vssd1 vssd1 vccd1 vccd1 _04912_/B1
+ sky130_fd_sc_hd__ebufn_2
XANTENNA__12836__D line[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07272_ _07272_/A _07279_/Y vssd1 vssd1 vccd1 vccd1 _13712_/Z sky130_fd_sc_hd__ebufn_2
X_09011_ _09025_/CLK line[66] vssd1 vssd1 vccd1 vccd1 _09012_/A sky130_fd_sc_hd__dfxtp_1
X_06223_ _06225_/CLK line[72] vssd1 vssd1 vccd1 vccd1 _06224_/A sky130_fd_sc_hd__dfxtp_1
X_06154_ _06154_/A _06159_/Y vssd1 vssd1 vccd1 vccd1 _13714_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_117_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05105_ _05105_/CLK line[73] vssd1 vssd1 vccd1 vccd1 _05106_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12571__D line[44] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06085_ _06085_/CLK line[9] vssd1 vssd1 vccd1 vccd1 _06086_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_132_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07665__D line[96] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05036_ _05036_/A _05039_/Y vssd1 vssd1 vccd1 vccd1 _13716_/Z sky130_fd_sc_hd__ebufn_2
X_09913_ _09935_/CLK line[109] vssd1 vssd1 vccd1 vccd1 _09914_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11187__D line[37] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09844_ _09844_/A _09869_/Y vssd1 vssd1 vccd1 vccd1 _13764_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_112_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09880__D line[94] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06859__A _13905_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09775_ _09795_/CLK line[46] vssd1 vssd1 vccd1 vccd1 _09776_/A sky130_fd_sc_hd__dfxtp_1
X_06987_ _06995_/CLK line[37] vssd1 vssd1 vccd1 vccd1 _06988_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_100_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06578__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08726_ _08726_/A _08749_/Y vssd1 vssd1 vccd1 vccd1 _13766_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08496__D line[87] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[21\].VALID\[7\].FF OVHB\[21\].V/CLK A[14] vssd1 vssd1 vccd1 vccd1 OVHB\[21\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_05938_ _05938_/A _05949_/Y vssd1 vssd1 vccd1 vccd1 _13778_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_100_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_OVHB\[27\].VALID\[14\].FF_D A[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08657_ _08675_/CLK line[47] vssd1 vssd1 vccd1 vccd1 _08658_/A sky130_fd_sc_hd__dfxtp_1
X_05869_ _05875_/CLK line[38] vssd1 vssd1 vccd1 vccd1 _05870_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07608_ _07608_/A _07629_/Y vssd1 vssd1 vccd1 vccd1 _13768_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08588_ _08588_/A _08609_/Y vssd1 vssd1 vccd1 vccd1 _13628_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_DATA\[11\].CLKBUF\[6\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07539_ _07555_/CLK line[33] vssd1 vssd1 vccd1 vccd1 _07540_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12746__D line[124] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11650__D line[121] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[28\].CG clk OVHB\[28\].CGAND/X vssd1 vssd1 vccd1 vccd1 OVHB\[28\].V/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_139_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10550_ _10550_/A _10569_/Y vssd1 vssd1 vccd1 vccd1 _13630_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06744__D line[54] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09120__D line[116] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05003__A _13931_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09209_ _09235_/CLK line[43] vssd1 vssd1 vccd1 vccd1 _09210_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_155_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10481_ _10495_/CLK line[98] vssd1 vssd1 vccd1 vccd1 _10482_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_5_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XDATA\[5\].CLKBUF\[5\] clk vssd1 vssd1 vccd1 vccd1 _12702_/CLK sky130_fd_sc_hd__clkbuf_4
X_12220_ _12220_/A _12249_/Y vssd1 vssd1 vccd1 vccd1 _13620_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_204_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XOVHB\[11\].VALID\[7\].TOBUF OVHB\[11\].VALID\[7\].FF/Q OVHB\[11\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/A2 sky130_fd_sc_hd__ebufn_2
X_12151_ _12175_/CLK line[108] vssd1 vssd1 vccd1 vccd1 _12152_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_123_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11102_ _11102_/A _11129_/Y vssd1 vssd1 vccd1 vccd1 _13622_/Z sky130_fd_sc_hd__ebufn_2
X_12082_ _12082_/A _12109_/Y vssd1 vssd1 vccd1 vccd1 _13762_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11097__D line[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11033_ _11055_/CLK line[109] vssd1 vssd1 vccd1 vccd1 _11034_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[4\].CLKBUF\[6\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05095__D line[68] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11825__D line[73] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06919__D line[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12984_ _13937_/X vssd1 vssd1 vccd1 vccd1 _12984_/Y sky130_fd_sc_hd__inv_2
XFILLER_94_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_DEC.DEC0.AND0_B A[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11935_ _11965_/CLK line[0] vssd1 vssd1 vccd1 vccd1 _11936_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_72_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11866_ _11866_/A _11899_/Y vssd1 vssd1 vccd1 vccd1 _13826_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[19\].VALID\[11\].FF_D A[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13605_ _13605_/A _13614_/Y vssd1 vssd1 vccd1 vccd1 _13885_/Z sky130_fd_sc_hd__ebufn_2
X_10817_ _10845_/CLK line[10] vssd1 vssd1 vccd1 vccd1 _10818_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11560__D line[94] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11797_ _11825_/CLK line[74] vssd1 vssd1 vccd1 vccd1 _11798_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06654__D line[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13536_ _13540_/CLK line[87] vssd1 vssd1 vccd1 vccd1 _13537_/A sky130_fd_sc_hd__dfxtp_1
X_10748_ _10748_/A _10779_/Y vssd1 vssd1 vccd1 vccd1 _13828_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09030__D line[80] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10176__D line[87] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13467_ _13467_/A _13474_/Y vssd1 vssd1 vccd1 vccd1 _13747_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_146_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10679_ _10705_/CLK line[75] vssd1 vssd1 vccd1 vccd1 _10680_/A sky130_fd_sc_hd__dfxtp_1
X_12418_ _12420_/CLK line[88] vssd1 vssd1 vccd1 vccd1 _12419_/A sky130_fd_sc_hd__dfxtp_1
X_13398_ _13400_/CLK line[24] vssd1 vssd1 vccd1 vccd1 _13399_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08224__A _13932_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13487__D line[79] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12349_ _12349_/A _12354_/Y vssd1 vssd1 vccd1 vccd1 _13749_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_99_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07485__D line[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[29\].VALID\[10\].FF_D A[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XDATA\[4\].CLKBUF\[2\] clk vssd1 vssd1 vccd1 vccd1 _12317_/CLK sky130_fd_sc_hd__clkbuf_4
X_06910_ _06910_/A _06929_/Y vssd1 vssd1 vccd1 vccd1 _13630_/Z sky130_fd_sc_hd__ebufn_2
X_07890_ _07890_/A _07909_/Y vssd1 vssd1 vccd1 vccd1 _13770_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_95_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06841_ _06855_/CLK line[98] vssd1 vssd1 vccd1 vccd1 _06842_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_67_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11735__D line[46] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09560_ _09560_/A _09589_/Y vssd1 vssd1 vccd1 vccd1 _13760_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[16\].VALID\[13\].TOBUF OVHB\[16\].VALID\[13\].FF/Q OVHB\[16\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04916_/B2 sky130_fd_sc_hd__ebufn_2
X_06772_ _06772_/A _06789_/Y vssd1 vssd1 vccd1 vccd1 _13772_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06829__D line[107] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05733__D line[104] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09205__D line[32] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08511_ _08535_/CLK line[108] vssd1 vssd1 vccd1 vccd1 _08512_/A sky130_fd_sc_hd__dfxtp_1
X_05723_ _05735_/CLK line[99] vssd1 vssd1 vccd1 vccd1 _05724_/A sky130_fd_sc_hd__dfxtp_1
X_09491_ _09515_/CLK line[44] vssd1 vssd1 vccd1 vccd1 _09492_/A sky130_fd_sc_hd__dfxtp_1
X_08442_ _08442_/A _08469_/Y vssd1 vssd1 vccd1 vccd1 _13762_/Z sky130_fd_sc_hd__ebufn_2
X_05654_ _05654_/A _05669_/Y vssd1 vssd1 vccd1 vccd1 _13774_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_211_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08373_ _08395_/CLK line[45] vssd1 vssd1 vccd1 vccd1 _08374_/A sky130_fd_sc_hd__dfxtp_1
X_05585_ _05595_/CLK line[36] vssd1 vssd1 vccd1 vccd1 _05586_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_51_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08118__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07324_ _07324_/A _07349_/Y vssd1 vssd1 vccd1 vccd1 _13764_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_149_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10086__D line[60] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07255_ _07275_/CLK line[46] vssd1 vssd1 vccd1 vccd1 _07256_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[24\].CLKBUF\[6\] clk vssd1 vssd1 vccd1 vccd1 _09657_/CLK sky130_fd_sc_hd__clkbuf_4
X_06206_ _06206_/A _06229_/Y vssd1 vssd1 vccd1 vccd1 _13766_/Z sky130_fd_sc_hd__ebufn_2
X_07186_ _07186_/A _07209_/Y vssd1 vssd1 vccd1 vccd1 _13626_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_133_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MUX.M\[3\].MUX\[1\]_A0 _13681_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06137_ _06155_/CLK line[47] vssd1 vssd1 vccd1 vccd1 _06138_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_105_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07395__D line[110] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05908__D line[56] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06068_ _06068_/A _06089_/Y vssd1 vssd1 vccd1 vccd1 _13628_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_105_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[1\].VALID\[5\].FF_D A[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05019_ _05035_/CLK line[33] vssd1 vssd1 vccd1 vccd1 _05020_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_59_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MUX.SEL0BUF\[0\]_A A[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05493__A _13900_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09827_ _09827_/A _09834_/Y vssd1 vssd1 vccd1 vccd1 _13747_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_104_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09758_ _09760_/CLK line[24] vssd1 vssd1 vccd1 vccd1 _09759_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05643__D line[77] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08709_ _08709_/A _08714_/Y vssd1 vssd1 vccd1 vccd1 _13749_/Z sky130_fd_sc_hd__ebufn_2
X_09689_ _09689_/A _09694_/Y vssd1 vssd1 vccd1 vccd1 _13889_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_15_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_DATA\[25\].CLKBUF\[0\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13860__D line[112] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ _11720_/CLK line[25] vssd1 vssd1 vccd1 vccd1 _11721_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_15_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11651_ _11651_/A _11654_/Y vssd1 vssd1 vccd1 vccd1 _13891_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_14_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12476__D line[114] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10602_ _10602_/CLK _10603_/X vssd1 vssd1 vccd1 vccd1 _10600_/CLK sky130_fd_sc_hd__dlclkp_1
XPHY_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11582_ _11582_/CLK _11583_/X vssd1 vssd1 vccd1 vccd1 _11580_/CLK sky130_fd_sc_hd__dlclkp_1
XPHY_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12773__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13321_ _13321_/A _13334_/Y vssd1 vssd1 vccd1 vccd1 _13881_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_210_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10533_ _13923_/X wr vssd1 vssd1 vccd1 vccd1 _10533_/X sky130_fd_sc_hd__and2_1
XPHY_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09785__D line[36] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05668__A _13901_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13252_ _13260_/CLK line[85] vssd1 vssd1 vccd1 vccd1 _13253_/A sky130_fd_sc_hd__dfxtp_1
X_10464_ _13923_/X vssd1 vssd1 vccd1 vccd1 _10464_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12203_ _12203_/A _12214_/Y vssd1 vssd1 vccd1 vccd1 _13883_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[26\].VALID\[1\].TOBUF OVHB\[26\].VALID\[1\].FF/Q OVHB\[26\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04926_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__10724__D line[81] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13183_ _13183_/A _13194_/Y vssd1 vssd1 vccd1 vccd1 _13743_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13100__D line[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10395_ _10425_/CLK line[64] vssd1 vssd1 vccd1 vccd1 _10396_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05818__D line[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12134_ _12140_/CLK line[86] vssd1 vssd1 vccd1 vccd1 _12135_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[23\].CLKBUF\[3\] clk vssd1 vssd1 vccd1 vccd1 _09272_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_1_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12065_ _12065_/A _12074_/Y vssd1 vssd1 vccd1 vccd1 _13745_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_77_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11016_ _11020_/CLK line[87] vssd1 vssd1 vccd1 vccd1 _11017_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_77_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09025__D line[73] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12948__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12967_ _12967_/A _12984_/Y vssd1 vssd1 vccd1 vccd1 _13807_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_45_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[16\].VALID\[2\].FF_D A[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11918_ _11930_/CLK line[115] vssd1 vssd1 vccd1 vccd1 _11919_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_205_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12898_ _12910_/CLK line[51] vssd1 vssd1 vccd1 vccd1 _12899_/A sky130_fd_sc_hd__dfxtp_1
X_11849_ _11849_/A _11864_/Y vssd1 vssd1 vccd1 vccd1 _13809_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[25\].CGAND _13921_/X wr vssd1 vssd1 vccd1 vccd1 OVHB\[25\].CGAND/X sky130_fd_sc_hd__and2_4
XANTENNA__11290__D line[84] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06384__D line[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05370_ _05370_/A _05389_/Y vssd1 vssd1 vccd1 vccd1 _13770_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_9_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13519_ _13519_/A _13544_/Y vssd1 vssd1 vccd1 vccd1 _13799_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09695__D line[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07040_ _07040_/A _07069_/Y vssd1 vssd1 vccd1 vccd1 _13760_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08889__A _13915_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08991_ _08991_/A _08994_/Y vssd1 vssd1 vccd1 vccd1 _13751_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_130_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[18\].VALID\[7\].TOBUF OVHB\[18\].VALID\[7\].FF/Q OVHB\[18\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/A2 sky130_fd_sc_hd__ebufn_2
X_07942_ _07942_/CLK _07943_/X vssd1 vssd1 vccd1 vccd1 _07940_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_68_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07873_ _13912_/X wr vssd1 vssd1 vccd1 vccd1 _07873_/X sky130_fd_sc_hd__and2_1
XANTENNA__11465__D line[36] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[7\].VALID\[9\].FF_D A[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDATA\[22\].CLKBUF\[0\] clk vssd1 vssd1 vccd1 vccd1 _08887_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_95_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09612_ _09620_/CLK line[85] vssd1 vssd1 vccd1 vccd1 _09613_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_68_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06824_ _13905_/X vssd1 vssd1 vccd1 vccd1 _06824_/Y sky130_fd_sc_hd__inv_2
XANTENNA__06559__D line[97] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDATA\[12\].CLKBUF\[6\] clk vssd1 vssd1 vccd1 vccd1 _06017_/CLK sky130_fd_sc_hd__clkbuf_4
X_09543_ _09543_/A _09554_/Y vssd1 vssd1 vccd1 vccd1 _13743_/Z sky130_fd_sc_hd__ebufn_2
X_06755_ _06785_/CLK line[64] vssd1 vssd1 vccd1 vccd1 _06756_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_36_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13680__D line[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05706_ _05706_/A _05739_/Y vssd1 vssd1 vccd1 vccd1 _13826_/Z sky130_fd_sc_hd__ebufn_2
X_09474_ _09480_/CLK line[22] vssd1 vssd1 vccd1 vccd1 _09475_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08774__D line[86] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06686_ _06686_/A _06719_/Y vssd1 vssd1 vccd1 vccd1 _13686_/Z sky130_fd_sc_hd__ebufn_2
XPHY_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07033__A _13909_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08425_ _08425_/A _08434_/Y vssd1 vssd1 vccd1 vccd1 _13745_/Z sky130_fd_sc_hd__ebufn_2
X_05637_ _05665_/CLK line[74] vssd1 vssd1 vccd1 vccd1 _05638_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_51_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08356_ _08360_/CLK line[23] vssd1 vssd1 vccd1 vccd1 _08357_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05568_ _05568_/A _05599_/Y vssd1 vssd1 vccd1 vccd1 _13688_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_50_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07307_ _07307_/A _07314_/Y vssd1 vssd1 vccd1 vccd1 _13747_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_137_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10394__A _13923_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08287_ _08287_/A _08294_/Y vssd1 vssd1 vccd1 vccd1 _13887_/Z sky130_fd_sc_hd__ebufn_2
X_05499_ _05525_/CLK line[11] vssd1 vssd1 vccd1 vccd1 _05500_/A sky130_fd_sc_hd__dfxtp_1
X_07238_ _07240_/CLK line[24] vssd1 vssd1 vccd1 vccd1 _07239_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_166_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XOVHB\[3\].INV _13978_/X vssd1 vssd1 vccd1 vccd1 OVHB\[3\].INV/Y sky130_fd_sc_hd__inv_2
XFILLER_118_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07169_ _07169_/A _07174_/Y vssd1 vssd1 vccd1 vccd1 _13889_/Z sky130_fd_sc_hd__ebufn_2
X_10180_ _10180_/CLK line[89] vssd1 vssd1 vccd1 vccd1 _10181_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13855__D line[105] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08949__D line[38] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07208__A _13910_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11375__D line[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13870_ _13890_/CLK line[126] vssd1 vssd1 vccd1 vccd1 _13871_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[29\].VALID\[2\].FF_D A[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05373__D line[67] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[27\].VALID\[14\].FF OVHB\[27\].V/CLK A[21] vssd1 vssd1 vccd1 vccd1 OVHB\[27\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_12821_ _12821_/A _12844_/Y vssd1 vssd1 vccd1 vccd1 _13661_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13590__D line[126] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10569__A _13924_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[24\].VALID\[6\].TOBUF OVHB\[24\].VALID\[6\].FF/Q OVHB\[24\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04923_/A2 sky130_fd_sc_hd__ebufn_2
XFILLER_43_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08684__D line[59] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12752_ _12770_/CLK line[127] vssd1 vssd1 vccd1 vccd1 _12753_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10288__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11703_ _11703_/A _11724_/Y vssd1 vssd1 vccd1 vccd1 _13663_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12683_ _12683_/A _12704_/Y vssd1 vssd1 vccd1 vccd1 _13803_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XDATA\[11\].CLKBUF\[3\] clk vssd1 vssd1 vccd1 vccd1 _05632_/CLK sky130_fd_sc_hd__clkbuf_4
XPHY_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11634_ _11650_/CLK line[113] vssd1 vssd1 vccd1 vccd1 _11635_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_DATA\[23\].CLKBUF\[2\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11565_ _11565_/A _11584_/Y vssd1 vssd1 vccd1 vccd1 _13805_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13304_ _13330_/CLK line[123] vssd1 vssd1 vccd1 vccd1 _13305_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06932__D line[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10516_ _10530_/CLK line[114] vssd1 vssd1 vccd1 vccd1 _10517_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_156_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11496_ _11510_/CLK line[50] vssd1 vssd1 vccd1 vccd1 _11497_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10454__D line[86] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13235_ _13235_/A _13264_/Y vssd1 vssd1 vccd1 vccd1 _13795_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_143_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[9\].VALID\[5\].FF OVHB\[9\].V/CLK A[12] vssd1 vssd1 vccd1 vccd1 OVHB\[9\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_155_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10447_ _10447_/A _10464_/Y vssd1 vssd1 vccd1 vccd1 _13807_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_6_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05548__D line[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13166_ _13190_/CLK line[60] vssd1 vssd1 vccd1 vccd1 _13167_/A sky130_fd_sc_hd__dfxtp_1
X_10378_ _10390_/CLK line[51] vssd1 vssd1 vccd1 vccd1 _10379_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13765__D line[78] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12117_ _12117_/A _12144_/Y vssd1 vssd1 vccd1 vccd1 _13797_/Z sky130_fd_sc_hd__ebufn_2
X_13097_ _13097_/A _13124_/Y vssd1 vssd1 vccd1 vccd1 _13657_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08859__D line[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07763__D line[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12048_ _12070_/CLK line[61] vssd1 vssd1 vccd1 vccd1 _12049_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11863__A _13927_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06540_ _06540_/CLK line[89] vssd1 vssd1 vccd1 vccd1 _06541_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_179_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06471_ _06471_/A _06474_/Y vssd1 vssd1 vccd1 vccd1 _13751_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10629__D line[38] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13005__D line[100] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08210_ _08220_/CLK line[84] vssd1 vssd1 vccd1 vccd1 _08211_/A sky130_fd_sc_hd__dfxtp_1
X_05422_ _05422_/CLK _05423_/X vssd1 vssd1 vccd1 vccd1 _05420_/CLK sky130_fd_sc_hd__dlclkp_1
X_09190_ _09200_/CLK line[20] vssd1 vssd1 vccd1 vccd1 _09191_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_21_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08141_ _08141_/A _08154_/Y vssd1 vssd1 vccd1 vccd1 _13741_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[6\].V OVHB\[6\].V/CLK TIE/HI rst_n vssd1 vssd1 vccd1 vccd1 OVHB\[6\].V/Q sky130_fd_sc_hd__dfrtp_1
X_05353_ _13900_/X wr vssd1 vssd1 vccd1 vccd1 _05353_/X sky130_fd_sc_hd__and2_1
XANTENNA__07938__D line[88] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08072_ _08080_/CLK line[21] vssd1 vssd1 vccd1 vccd1 _08073_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[10\].CLKBUF\[0\] clk vssd1 vssd1 vccd1 vccd1 _05247_/CLK sky130_fd_sc_hd__clkbuf_4
X_05284_ _13900_/X vssd1 vssd1 vccd1 vccd1 _05284_/Y sky130_fd_sc_hd__inv_2
XOVHB\[30\].VALID\[5\].TOBUF OVHB\[30\].VALID\[5\].FF/Q OVHB\[30\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04927_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__10364__D line[59] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07023_ _07023_/A _07034_/Y vssd1 vssd1 vccd1 vccd1 _13743_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_162_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08974_ _08990_/CLK line[49] vssd1 vssd1 vccd1 vccd1 _08975_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[6\].V_RESET_B rst_n vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07673__D line[109] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07925_ _07925_/A _07944_/Y vssd1 vssd1 vccd1 vccd1 _13805_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_69_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11195__D line[41] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[7\].VALID\[7\].FF OVHB\[7\].V/CLK A[14] vssd1 vssd1 vccd1 vccd1 OVHB\[7\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06289__D line[102] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07856_ _07870_/CLK line[50] vssd1 vssd1 vccd1 vccd1 _07857_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_45_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06807_ _06807_/A _06824_/Y vssd1 vssd1 vccd1 vccd1 _13807_/Z sky130_fd_sc_hd__ebufn_2
X_07787_ _07787_/A _07804_/Y vssd1 vssd1 vccd1 vccd1 _13667_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_43_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_04999_ _04999_/A _05004_/Y vssd1 vssd1 vccd1 vccd1 _13679_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_71_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09526_ _09550_/CLK line[60] vssd1 vssd1 vccd1 vccd1 _09527_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_43_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06738_ _06750_/CLK line[51] vssd1 vssd1 vccd1 vccd1 _06739_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__04931__B2 _04931_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05921__D line[76] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10539__D line[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09457_ _09457_/A _09484_/Y vssd1 vssd1 vccd1 vccd1 _13657_/Z sky130_fd_sc_hd__ebufn_2
X_06669_ _06669_/A _06684_/Y vssd1 vssd1 vccd1 vccd1 _13669_/Z sky130_fd_sc_hd__ebufn_2
XPHY_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08408_ _08430_/CLK line[61] vssd1 vssd1 vccd1 vccd1 _08409_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07698__A _13911_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09388_ _09410_/CLK line[125] vssd1 vssd1 vccd1 vccd1 _09389_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[3\].CG_CLK clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08339_ _08339_/A _08364_/Y vssd1 vssd1 vccd1 vccd1 _13659_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12754__D line[113] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12109__A _13934_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07848__D line[61] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11350_ _11370_/CLK line[126] vssd1 vssd1 vccd1 vccd1 _11351_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_138_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10301_ _10301_/A _10324_/Y vssd1 vssd1 vccd1 vccd1 _13661_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_137_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11281_ _11281_/A _11304_/Y vssd1 vssd1 vccd1 vccd1 _13801_/Z sky130_fd_sc_hd__ebufn_2
X_13020_ _13050_/CLK line[112] vssd1 vssd1 vccd1 vccd1 _13021_/A sky130_fd_sc_hd__dfxtp_1
X_10232_ _10250_/CLK line[127] vssd1 vssd1 vccd1 vccd1 _10233_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_4_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10163_ _10163_/A _10184_/Y vssd1 vssd1 vccd1 vccd1 _13803_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_126_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10094_ _10110_/CLK line[49] vssd1 vssd1 vccd1 vccd1 _10095_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_47_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13922_ _13927_/C _13927_/A _13927_/B _13927_/D vssd1 vssd1 vccd1 vccd1 _13922_/X
+ sky130_fd_sc_hd__and4bb_4
XANTENNA__06199__D line[75] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[12\].VALID\[5\].FF_D A[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[20\].V OVHB\[20\].V/CLK TIE/HI rst_n vssd1 vssd1 vccd1 vccd1 OVHB\[20\].V/Q
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_19_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12929__D line[65] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13853_ _13855_/CLK line[104] vssd1 vssd1 vccd1 vccd1 _13854_/A sky130_fd_sc_hd__dfxtp_1
X_12804_ _12804_/A _12809_/Y vssd1 vssd1 vccd1 vccd1 _13644_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__04922__B2 _04922_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13784_ _13784_/A _13789_/Y vssd1 vssd1 vccd1 vccd1 _13784_/Z sky130_fd_sc_hd__ebufn_2
X_10996_ _11020_/CLK line[92] vssd1 vssd1 vccd1 vccd1 _10997_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09303__D line[72] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[5\].VALID\[9\].FF OVHB\[5\].V/CLK A[16] vssd1 vssd1 vccd1 vccd1 OVHB\[5\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12735_ _12735_/CLK line[105] vssd1 vssd1 vccd1 vccd1 _12736_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_203_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13403__A _13898_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12666_ _12666_/A _12669_/Y vssd1 vssd1 vccd1 vccd1 _13786_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11617_ _11617_/CLK _11618_/X vssd1 vssd1 vccd1 vccd1 _11615_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_187_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12597_ _12597_/CLK _12598_/X vssd1 vssd1 vccd1 vccd1 _12595_/CLK sky130_fd_sc_hd__dlclkp_1
XPHY_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06662__D line[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11548_ _13926_/X wr vssd1 vssd1 vccd1 vccd1 _11548_/X sky130_fd_sc_hd__and2_1
XOVHB\[26\].VALID\[11\].TOBUF OVHB\[26\].VALID\[11\].FF/Q OVHB\[26\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04915_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_143_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11479_ _13926_/X vssd1 vssd1 vccd1 vccd1 _11479_/Y sky130_fd_sc_hd__inv_2
XANTENNA__05278__D line[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13218_ _13218_/A _13229_/Y vssd1 vssd1 vccd1 vccd1 _13778_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_171_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_DATA\[21\].CLKBUF\[4\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13495__D line[68] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[23\].VALID\[12\].FF OVHB\[23\].V/CLK A[19] vssd1 vssd1 vccd1 vccd1 OVHB\[23\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08589__D line[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13149_ _13155_/CLK line[38] vssd1 vssd1 vccd1 vccd1 _13150_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05971_ _05971_/A _05984_/Y vssd1 vssd1 vccd1 vccd1 _13811_/Z sky130_fd_sc_hd__ebufn_2
X_07710_ _07730_/CLK line[126] vssd1 vssd1 vccd1 vccd1 _07711_/A sky130_fd_sc_hd__dfxtp_1
X_04922_ _04913_/Y _04922_/A2 _04920_/Y _04922_/B2 vssd1 vssd1 vccd1 vccd1 _04922_/X
+ sky130_fd_sc_hd__o22a_2
X_08690_ _08710_/CLK line[62] vssd1 vssd1 vccd1 vccd1 _08691_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_66_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XOVHB\[11\].V OVHB\[11\].V/CLK TIE/HI rst_n vssd1 vssd1 vccd1 vccd1 OVHB\[11\].V/Q
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09063__A _13915_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07641_ _07641_/A _07664_/Y vssd1 vssd1 vccd1 vccd1 _13801_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_65_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11743__D line[35] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07572_ _07590_/CLK line[63] vssd1 vssd1 vccd1 vccd1 _07573_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06837__D line[111] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09213__D line[45] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09311_ _09311_/A _09344_/Y vssd1 vssd1 vccd1 vccd1 _13791_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_80_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06523_ _06523_/A _06544_/Y vssd1 vssd1 vccd1 vccd1 _13803_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[6\].VALID\[3\].TOBUF OVHB\[6\].VALID\[3\].FF/Q OVHB\[6\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04919_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[4\].VALID\[14\].FF_D A[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09242_ _09270_/CLK line[58] vssd1 vssd1 vccd1 vccd1 _09243_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_194_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06454_ _06470_/CLK line[49] vssd1 vssd1 vccd1 vccd1 _06455_/A sky130_fd_sc_hd__dfxtp_1
X_05405_ _05405_/A _05424_/Y vssd1 vssd1 vccd1 vccd1 _13805_/Z sky130_fd_sc_hd__ebufn_2
X_09173_ _09173_/A _09204_/Y vssd1 vssd1 vccd1 vccd1 _13653_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_194_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06385_ _06385_/A _06404_/Y vssd1 vssd1 vccd1 vccd1 _13665_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[13\].VALID\[14\].FF OVHB\[13\].V/CLK A[21] vssd1 vssd1 vccd1 vccd1 OVHB\[13\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_31_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08124_ _08150_/CLK line[59] vssd1 vssd1 vccd1 vccd1 _08125_/A sky130_fd_sc_hd__dfxtp_1
X_05336_ _05350_/CLK line[50] vssd1 vssd1 vccd1 vccd1 _05337_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_174_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10094__D line[49] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08055_ _08055_/A _08084_/Y vssd1 vssd1 vccd1 vccd1 _13655_/Z sky130_fd_sc_hd__ebufn_2
X_05267_ _05267_/A _05284_/Y vssd1 vssd1 vccd1 vccd1 _13667_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05188__D line[125] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07006_ _07030_/CLK line[60] vssd1 vssd1 vccd1 vccd1 _07007_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09238__A _13916_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05198_ _05210_/CLK line[115] vssd1 vssd1 vccd1 vccd1 _05199_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11918__D line[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_OVHB\[25\].VALID\[5\].FF_D A[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08957_ _08957_/CLK _08958_/X vssd1 vssd1 vccd1 vccd1 _08955_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__12599__A _13936_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07908_ _13912_/X wr vssd1 vssd1 vccd1 vccd1 _07908_/X sky130_fd_sc_hd__and2_1
X_08888_ _13915_/X wr vssd1 vssd1 vccd1 vccd1 _08888_/X sky130_fd_sc_hd__and2_1
X_07839_ _13912_/X vssd1 vssd1 vccd1 vccd1 _07839_/Y sky130_fd_sc_hd__inv_2
X_10850_ _10880_/CLK line[16] vssd1 vssd1 vccd1 vccd1 _10851_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_112_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05651__D line[66] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[18\].VALID\[9\].FF_D A[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10269__D line[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09509_ _09515_/CLK line[38] vssd1 vssd1 vccd1 vccd1 _09510_/A sky130_fd_sc_hd__dfxtp_1
X_10781_ _10781_/A _10814_/Y vssd1 vssd1 vccd1 vccd1 _13861_/Z sky130_fd_sc_hd__ebufn_2
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12520_ _12520_/A _12529_/Y vssd1 vssd1 vccd1 vccd1 _13640_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08962__D line[58] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XOVHB\[14\].VALID\[1\].FF OVHB\[14\].V/CLK A[8] vssd1 vssd1 vccd1 vccd1 OVHB\[14\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_185_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12451_ _12455_/CLK line[103] vssd1 vssd1 vccd1 vccd1 _12452_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12484__D line[118] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07578__D line[51] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[31\].VALID\[5\].FF OVHB\[31\].V/CLK A[12] vssd1 vssd1 vccd1 vccd1 OVHB\[31\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_11402_ _11402_/A _11409_/Y vssd1 vssd1 vccd1 vccd1 _13642_/Z sky130_fd_sc_hd__ebufn_2
X_12382_ _12382_/A _12389_/Y vssd1 vssd1 vccd1 vccd1 _13782_/Z sky130_fd_sc_hd__ebufn_2
X_11333_ _11335_/CLK line[104] vssd1 vssd1 vccd1 vccd1 _11334_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09793__D line[40] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11264_ _11264_/A _11269_/Y vssd1 vssd1 vccd1 vccd1 _13784_/Z sky130_fd_sc_hd__ebufn_2
X_13003_ _13015_/CLK line[99] vssd1 vssd1 vccd1 vccd1 _13004_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10732__D line[85] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13893__A _13899_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10215_ _10215_/CLK line[105] vssd1 vssd1 vccd1 vccd1 _10216_/A sky130_fd_sc_hd__dfxtp_1
X_11195_ _11195_/CLK line[41] vssd1 vssd1 vccd1 vccd1 _11196_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05826__D line[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10146_ _10146_/A _10149_/Y vssd1 vssd1 vccd1 vccd1 _13786_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08202__D line[95] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_OVHB\[6\].VALID\[10\].FF_D A[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10077_ _10077_/CLK _10078_/X vssd1 vssd1 vccd1 vccd1 _10075_/CLK sky130_fd_sc_hd__dlclkp_1
X_13905_ _13905_/A _13905_/B _13905_/C _13905_/D vssd1 vssd1 vccd1 vccd1 _13905_/X
+ sky130_fd_sc_hd__and4_4
XANTENNA__12659__D line[70] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13836_ _13836_/A _13859_/Y vssd1 vssd1 vccd1 vccd1 _13836_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XDATA\[2\].CLKBUF\[7\] clk vssd1 vssd1 vccd1 vccd1 _11372_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_31_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10979_ _10985_/CLK line[70] vssd1 vssd1 vccd1 vccd1 _10980_/A sky130_fd_sc_hd__dfxtp_1
X_13767_ _13785_/CLK line[79] vssd1 vssd1 vccd1 vccd1 _13768_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_90_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09968__D line[120] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_OVHB\[6\].VALID\[0\].FF_D A[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12718_ _12718_/A _12739_/Y vssd1 vssd1 vccd1 vccd1 _13838_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_31_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13698_ _13698_/A _13719_/Y vssd1 vssd1 vccd1 vccd1 _13698_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12394__D line[91] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10907__D line[37] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12649_ _12665_/CLK line[65] vssd1 vssd1 vccd1 vccd1 _12650_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_176_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06392__D line[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06170_ _06190_/CLK line[62] vssd1 vssd1 vccd1 vccd1 _06171_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_172_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05121_ _05121_/A _05144_/Y vssd1 vssd1 vccd1 vccd1 _13801_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_172_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[12\].VALID\[3\].FF OVHB\[12\].V/CLK A[10] vssd1 vssd1 vccd1 vccd1 OVHB\[12\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_05052_ _05070_/CLK line[63] vssd1 vssd1 vccd1 vccd1 _05053_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_171_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09860_ _09860_/A _09869_/Y vssd1 vssd1 vccd1 vccd1 _13780_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10642__D line[58] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[4\].VALID\[8\].TOBUF OVHB\[4\].VALID\[8\].FF/Q OVHB\[4\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04931_/B2 sky130_fd_sc_hd__ebufn_2
XOVHB\[13\].VOBUF OVHB\[13\].V/Q OVHB\[13\].INV/Y vssd1 vssd1 vccd1 vccd1 _04912_/B1
+ sky130_fd_sc_hd__ebufn_2
X_08811_ _08815_/CLK line[103] vssd1 vssd1 vccd1 vccd1 _08812_/A sky130_fd_sc_hd__dfxtp_1
X_09791_ _09795_/CLK line[39] vssd1 vssd1 vccd1 vccd1 _09792_/A sky130_fd_sc_hd__dfxtp_1
X_08742_ _08742_/A _08749_/Y vssd1 vssd1 vccd1 vccd1 _13782_/Z sky130_fd_sc_hd__ebufn_2
X_05954_ _05980_/CLK line[91] vssd1 vssd1 vccd1 vccd1 _05955_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_66_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07951__D line[108] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08673_ _08675_/CLK line[40] vssd1 vssd1 vccd1 vccd1 _08674_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12569__D line[43] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05885_ _05885_/A _05914_/Y vssd1 vssd1 vccd1 vccd1 _13725_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11473__D line[40] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07624_ _07624_/A _07629_/Y vssd1 vssd1 vccd1 vccd1 _13784_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06567__D line[101] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07555_ _07555_/CLK line[41] vssd1 vssd1 vccd1 vccd1 _07556_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09878__D line[93] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06506_ _06506_/A _06509_/Y vssd1 vssd1 vccd1 vccd1 _13786_/Z sky130_fd_sc_hd__ebufn_2
X_07486_ _07486_/A _07489_/Y vssd1 vssd1 vccd1 vccd1 _13646_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09225_ _09235_/CLK line[36] vssd1 vssd1 vccd1 vccd1 _09226_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10817__D line[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06437_ _06437_/CLK _06438_/X vssd1 vssd1 vccd1 vccd1 _06435_/CLK sky130_fd_sc_hd__dlclkp_1
XDATA\[1\].CLKBUF\[4\] clk vssd1 vssd1 vccd1 vccd1 _08187_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_210_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09156_ _09156_/A _09169_/Y vssd1 vssd1 vccd1 vccd1 _13636_/Z sky130_fd_sc_hd__ebufn_2
X_06368_ _13904_/X wr vssd1 vssd1 vccd1 vccd1 _06368_/X sky130_fd_sc_hd__and2_1
X_08107_ _08115_/CLK line[37] vssd1 vssd1 vccd1 vccd1 _08108_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_135_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05319_ _13900_/X vssd1 vssd1 vccd1 vccd1 _05319_/Y sky130_fd_sc_hd__inv_2
X_09087_ _09095_/CLK line[101] vssd1 vssd1 vccd1 vccd1 _09088_/A sky130_fd_sc_hd__dfxtp_1
X_06299_ _13903_/X vssd1 vssd1 vccd1 vccd1 _06299_/Y sky130_fd_sc_hd__inv_2
XFILLER_190_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08038_ _08038_/A _08049_/Y vssd1 vssd1 vccd1 vccd1 _13638_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[28\].VALID\[8\].FF OVHB\[28\].V/CLK A[15] vssd1 vssd1 vccd1 vccd1 OVHB\[28\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11648__D line[120] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10000_ _10000_/A _10009_/Y vssd1 vssd1 vccd1 vccd1 _13640_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09118__D line[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09989_ _10005_/CLK line[1] vssd1 vssd1 vccd1 vccd1 _09990_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XOVHB\[10\].VALID\[5\].FF OVHB\[10\].V/CLK A[12] vssd1 vssd1 vccd1 vccd1 OVHB\[10\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_184_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_OVHB\[11\].CGAND_B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XDATA\[31\].CLKBUF\[2\] clk vssd1 vssd1 vccd1 vccd1 _11757_/CLK sky130_fd_sc_hd__clkbuf_4
X_11951_ _11965_/CLK line[2] vssd1 vssd1 vccd1 vccd1 _11952_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11383__D line[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06477__D line[74] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10902_ _10902_/A _10919_/Y vssd1 vssd1 vccd1 vccd1 _13702_/Z sky130_fd_sc_hd__ebufn_2
X_11882_ _11882_/A _11899_/Y vssd1 vssd1 vccd1 vccd1 _13842_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[11\].VALID\[3\].TOBUF OVHB\[11\].VALID\[3\].FF/Q OVHB\[11\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04919_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__05381__D line[71] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[15\].CGAND_A _13905_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10833_ _10845_/CLK line[3] vssd1 vssd1 vccd1 vccd1 _10834_/A sky130_fd_sc_hd__dfxtp_1
X_13621_ _13645_/CLK line[12] vssd1 vssd1 vccd1 vccd1 _13622_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08692__D line[63] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13552_ _13552_/A _13579_/Y vssd1 vssd1 vccd1 vccd1 _13832_/Z sky130_fd_sc_hd__ebufn_2
X_10764_ _10764_/A _10779_/Y vssd1 vssd1 vccd1 vccd1 _13844_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DECH.DEC0.AND3_A A_h[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12503_ _12525_/CLK line[13] vssd1 vssd1 vccd1 vccd1 _12504_/A sky130_fd_sc_hd__dfxtp_1
X_13483_ _13505_/CLK line[77] vssd1 vssd1 vccd1 vccd1 _13484_/A sky130_fd_sc_hd__dfxtp_1
X_10695_ _10705_/CLK line[68] vssd1 vssd1 vccd1 vccd1 _10696_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_200_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12434_ _12434_/A _12459_/Y vssd1 vssd1 vccd1 vccd1 _13834_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_157_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12365_ _12385_/CLK line[78] vssd1 vssd1 vccd1 vccd1 _12366_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[0\].CLKBUF\[1\] clk vssd1 vssd1 vccd1 vccd1 _05002_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__06940__D line[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11316_ _11316_/A _11339_/Y vssd1 vssd1 vccd1 vccd1 _13836_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_99_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12296_ _12296_/A _12319_/Y vssd1 vssd1 vccd1 vccd1 _13696_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11558__D line[93] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11247_ _11265_/CLK line[79] vssd1 vssd1 vccd1 vccd1 _11248_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05556__D line[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11178_ _11178_/A _11199_/Y vssd1 vssd1 vccd1 vccd1 _13698_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13773__D line[67] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10129_ _10145_/CLK line[65] vssd1 vssd1 vccd1 vccd1 _10130_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[18\].CLKBUF\[7\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08867__D line[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05670_ _05700_/CLK line[80] vssd1 vssd1 vccd1 vccd1 _05671_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05291__D line[44] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13819_ _13819_/A _13824_/Y vssd1 vssd1 vccd1 vccd1 _13819_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_189_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07340_ _07340_/A _07349_/Y vssd1 vssd1 vccd1 vccd1 _13780_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_148_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07271_ _07275_/CLK line[39] vssd1 vssd1 vccd1 vccd1 _07272_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[20\].CLKBUF\[5\] clk vssd1 vssd1 vccd1 vccd1 _08502_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__13013__D line[104] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09010_ _09010_/A _09029_/Y vssd1 vssd1 vccd1 vccd1 _13770_/Z sky130_fd_sc_hd__ebufn_2
X_06222_ _06222_/A _06229_/Y vssd1 vssd1 vccd1 vccd1 _13782_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_191_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08107__D line[37] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06153_ _06155_/CLK line[40] vssd1 vssd1 vccd1 vccd1 _06154_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_129_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05104_ _05104_/A _05109_/Y vssd1 vssd1 vccd1 vccd1 _13784_/Z sky130_fd_sc_hd__ebufn_2
X_06084_ _06084_/A _06089_/Y vssd1 vssd1 vccd1 vccd1 _13644_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_171_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05035_ _05035_/CLK line[41] vssd1 vssd1 vccd1 vccd1 _05036_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10372__D line[63] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[21\].VALID\[8\].FF_D A[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09912_ _09912_/A _09939_/Y vssd1 vssd1 vccd1 vccd1 _13832_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_113_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05466__D line[124] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09843_ _09865_/CLK line[77] vssd1 vssd1 vccd1 vccd1 _09844_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_140_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06986_ _06986_/A _06999_/Y vssd1 vssd1 vccd1 vccd1 _13706_/Z sky130_fd_sc_hd__ebufn_2
X_09774_ _09774_/A _09799_/Y vssd1 vssd1 vccd1 vccd1 _13694_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_37_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07681__D line[98] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12299__D line[33] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08725_ _08745_/CLK line[78] vssd1 vssd1 vccd1 vccd1 _08726_/A sky130_fd_sc_hd__dfxtp_1
X_05937_ _05945_/CLK line[69] vssd1 vssd1 vccd1 vccd1 _05938_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_160_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08656_ _08656_/A _08679_/Y vssd1 vssd1 vccd1 vccd1 _13696_/Z sky130_fd_sc_hd__ebufn_2
X_05868_ _05868_/A _05879_/Y vssd1 vssd1 vccd1 vccd1 _13708_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07607_ _07625_/CLK line[79] vssd1 vssd1 vccd1 vccd1 _07608_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08587_ _08605_/CLK line[15] vssd1 vssd1 vccd1 vccd1 _08588_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_54_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05799_ _05805_/CLK line[6] vssd1 vssd1 vccd1 vccd1 _05800_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07538_ _07538_/A _07559_/Y vssd1 vssd1 vccd1 vccd1 _13698_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[4\].VALID\[14\].FF OVHB\[4\].V/CLK A[21] vssd1 vssd1 vccd1 vccd1 OVHB\[4\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_169_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10547__D line[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07469_ _07485_/CLK line[1] vssd1 vssd1 vccd1 vccd1 _07470_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_194_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05003__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09208_ _09208_/A _09239_/Y vssd1 vssd1 vccd1 vccd1 _13688_/Z sky130_fd_sc_hd__ebufn_2
X_10480_ _10480_/A _10499_/Y vssd1 vssd1 vccd1 vccd1 _13840_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08017__D line[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09139_ _09165_/CLK line[11] vssd1 vssd1 vccd1 vccd1 _09140_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12762__D line[117] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07856__D line[50] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12150_ _12150_/A _12179_/Y vssd1 vssd1 vccd1 vccd1 _13830_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_2_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11101_ _11125_/CLK line[12] vssd1 vssd1 vccd1 vccd1 _11102_/A sky130_fd_sc_hd__dfxtp_1
X_12081_ _12105_/CLK line[76] vssd1 vssd1 vccd1 vccd1 _12082_/A sky130_fd_sc_hd__dfxtp_1
X_11032_ _11032_/A _11059_/Y vssd1 vssd1 vccd1 vccd1 _13832_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_78_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12983_ _13937_/X wr vssd1 vssd1 vccd1 vccd1 _12983_/X sky130_fd_sc_hd__and2_1
X_11934_ _13927_/X vssd1 vssd1 vccd1 vccd1 _11934_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[2\].VALID\[3\].FF_D A[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12937__D line[69] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11865_ _11895_/CLK line[96] vssd1 vssd1 vccd1 vccd1 _11866_/A sky130_fd_sc_hd__dfxtp_1
X_13604_ _13610_/CLK line[118] vssd1 vssd1 vccd1 vccd1 _13605_/A sky130_fd_sc_hd__dfxtp_1
X_10816_ _10816_/A _10849_/Y vssd1 vssd1 vccd1 vccd1 _13616_/Z sky130_fd_sc_hd__ebufn_2
X_11796_ _11796_/A _11829_/Y vssd1 vssd1 vccd1 vccd1 _13756_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_201_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13535_ _13535_/A _13544_/Y vssd1 vssd1 vccd1 vccd1 _13815_/Z sky130_fd_sc_hd__ebufn_2
X_10747_ _10775_/CLK line[106] vssd1 vssd1 vccd1 vccd1 _10748_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[28\].VALID\[12\].FF OVHB\[28\].V/CLK A[19] vssd1 vssd1 vccd1 vccd1 OVHB\[28\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_10678_ _10678_/A _10709_/Y vssd1 vssd1 vccd1 vccd1 _13758_/Z sky130_fd_sc_hd__ebufn_2
X_13466_ _13470_/CLK line[55] vssd1 vssd1 vccd1 vccd1 _13467_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_173_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12417_ _12417_/A _12424_/Y vssd1 vssd1 vccd1 vccd1 _13817_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12672__D line[90] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[31\].VALID\[14\].FF_D A[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13397_ _13397_/A _13404_/Y vssd1 vssd1 vccd1 vccd1 _13677_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06670__D line[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12348_ _12350_/CLK line[56] vssd1 vssd1 vccd1 vccd1 _12349_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11288__D line[83] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[12\].VALID\[14\].TOBUF OVHB\[12\].VALID\[14\].FF/Q OVHB\[12\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_4_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12279_ _12279_/A _12284_/Y vssd1 vssd1 vccd1 vccd1 _13679_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09981__D line[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[21\].CGAND _13914_/X wr vssd1 vssd1 vccd1 vccd1 OVHB\[21\].CGAND/X sky130_fd_sc_hd__and2_4
XANTENNA__10920__D line[48] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06840_ _06840_/A _06859_/Y vssd1 vssd1 vccd1 vccd1 _13840_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08597__D line[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06771_ _06785_/CLK line[66] vssd1 vssd1 vccd1 vccd1 _06772_/A sky130_fd_sc_hd__dfxtp_1
X_08510_ _08510_/A _08539_/Y vssd1 vssd1 vccd1 vccd1 _13830_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_209_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05722_ _05722_/A _05739_/Y vssd1 vssd1 vccd1 vccd1 _13842_/Z sky130_fd_sc_hd__ebufn_2
X_09490_ _09490_/A _09519_/Y vssd1 vssd1 vccd1 vccd1 _13690_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07006__D line[60] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08441_ _08465_/CLK line[76] vssd1 vssd1 vccd1 vccd1 _08442_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[18\].VALID\[14\].FF OVHB\[18\].V/CLK A[21] vssd1 vssd1 vccd1 vccd1 OVHB\[18\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_05653_ _05665_/CLK line[67] vssd1 vssd1 vccd1 vccd1 _05654_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12847__D line[42] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[13\].VALID\[12\].FF_D A[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11751__D line[39] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08372_ _08372_/A _08399_/Y vssd1 vssd1 vccd1 vccd1 _13692_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06845__D line[100] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05584_ _05584_/A _05599_/Y vssd1 vssd1 vccd1 vccd1 _13704_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[18\].VALID\[3\].TOBUF OVHB\[18\].VALID\[3\].FF/Q OVHB\[18\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04919_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__09221__D line[34] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XOVHB\[1\].VALID\[0\].FF OVHB\[1\].V/CLK A[7] vssd1 vssd1 vccd1 vccd1 OVHB\[1\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_07323_ _07345_/CLK line[77] vssd1 vssd1 vccd1 vccd1 _07324_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_149_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_DATA\[12\].CLKBUF\[0\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07254_ _07254_/A _07279_/Y vssd1 vssd1 vccd1 vccd1 _13694_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13678__D line[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06205_ _06225_/CLK line[78] vssd1 vssd1 vccd1 vccd1 _06206_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[17\].VALID\[0\].FF_D A[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07185_ _07205_/CLK line[14] vssd1 vssd1 vccd1 vccd1 _07186_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_145_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06136_ _06136_/A _06159_/Y vssd1 vssd1 vccd1 vccd1 _13696_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06580__D line[112] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MUX.M\[3\].MUX\[1\]_A1 _13751_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[23\].VALID\[11\].FF_D A[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06067_ _06085_/CLK line[15] vssd1 vssd1 vccd1 vccd1 _06068_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_160_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05196__D line[114] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05018_ _05018_/A _05039_/Y vssd1 vssd1 vccd1 vccd1 _13698_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05774__A _13901_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11926__D line[119] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09826_ _09830_/CLK line[55] vssd1 vssd1 vccd1 vccd1 _09827_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05493__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[5\].CLKBUF\[0\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09757_ _09757_/A _09764_/Y vssd1 vssd1 vccd1 vccd1 _13677_/Z sky130_fd_sc_hd__ebufn_2
X_06969_ _06995_/CLK line[43] vssd1 vssd1 vccd1 vccd1 _06970_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_104_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08708_ _08710_/CLK line[56] vssd1 vssd1 vccd1 vccd1 _08709_/A sky130_fd_sc_hd__dfxtp_1
X_09688_ _09690_/CLK line[120] vssd1 vssd1 vccd1 vccd1 _09689_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_54_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_DATA\[31\].CLKBUF\[2\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08639_ _08639_/A _08644_/Y vssd1 vssd1 vccd1 vccd1 _13679_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11661__D line[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11650_ _11650_/CLK line[121] vssd1 vssd1 vccd1 vccd1 _11651_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06755__D line[64] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[8\].VALID\[7\].FF_D A[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10277__D line[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10601_ _10601_/A _10604_/Y vssd1 vssd1 vccd1 vccd1 _13681_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11581_ _11581_/A _11584_/Y vssd1 vssd1 vccd1 vccd1 _13821_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08970__D line[62] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05949__A _13902_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10532_ _10532_/CLK _10533_/X vssd1 vssd1 vccd1 vccd1 _10530_/CLK sky130_fd_sc_hd__dlclkp_1
X_13320_ _13330_/CLK line[116] vssd1 vssd1 vccd1 vccd1 _13321_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13588__D line[125] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05668__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10463_ _13923_/X wr vssd1 vssd1 vccd1 vccd1 _10463_/X sky130_fd_sc_hd__and2_1
X_13251_ _13251_/A _13264_/Y vssd1 vssd1 vccd1 vccd1 _13811_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07586__D line[55] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12202_ _12210_/CLK line[117] vssd1 vssd1 vccd1 vccd1 _12203_/A sky130_fd_sc_hd__dfxtp_1
X_13182_ _13190_/CLK line[53] vssd1 vssd1 vccd1 vccd1 _13183_/A sky130_fd_sc_hd__dfxtp_1
X_10394_ _13923_/X vssd1 vssd1 vccd1 vccd1 _10394_/Y sky130_fd_sc_hd__inv_2
XOVHB\[24\].VALID\[2\].TOBUF OVHB\[24\].VALID\[2\].FF/Q OVHB\[24\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04930_/B2 sky130_fd_sc_hd__ebufn_2
X_12133_ _12133_/A _12144_/Y vssd1 vssd1 vccd1 vccd1 _13813_/Z sky130_fd_sc_hd__ebufn_2
X_12064_ _12070_/CLK line[54] vssd1 vssd1 vccd1 vccd1 _12065_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_1_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11836__D line[92] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11015_ _11015_/A _11024_/Y vssd1 vssd1 vccd1 vccd1 _13815_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10740__D line[89] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05834__D line[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[0\].VALID\[12\].FF OVHB\[0\].V/CLK A[19] vssd1 vssd1 vccd1 vccd1 OVHB\[0\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08210__D line[84] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12966_ _12980_/CLK line[82] vssd1 vssd1 vccd1 vccd1 _12967_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_206_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11917_ _11917_/A _11934_/Y vssd1 vssd1 vccd1 vccd1 _13877_/Z sky130_fd_sc_hd__ebufn_2
X_12897_ _12897_/A _12914_/Y vssd1 vssd1 vccd1 vccd1 _13737_/Z sky130_fd_sc_hd__ebufn_2
X_11848_ _11860_/CLK line[83] vssd1 vssd1 vccd1 vccd1 _11849_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10187__D line[106] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11779_ _11779_/A _11794_/Y vssd1 vssd1 vccd1 vccd1 _13739_/Z sky130_fd_sc_hd__ebufn_2
X_13518_ _13540_/CLK line[93] vssd1 vssd1 vccd1 vccd1 _13519_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_158_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10915__D line[41] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13449_ _13449_/A _13474_/Y vssd1 vssd1 vccd1 vccd1 _13729_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_174_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07496__D line[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08990_ _08990_/CLK line[57] vssd1 vssd1 vccd1 vccd1 _08991_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[5\].V_RESET_B rst_n vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07941_ _07941_/A _07944_/Y vssd1 vssd1 vccd1 vccd1 _13821_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[16\].VALID\[8\].TOBUF OVHB\[16\].VALID\[8\].FF/Q OVHB\[16\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04931_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_205_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10650__D line[62] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07872_ _07872_/CLK _07873_/X vssd1 vssd1 vccd1 vccd1 _07870_/CLK sky130_fd_sc_hd__dlclkp_1
XOVHB\[18\].CG clk OVHB\[18\].CGAND/X vssd1 vssd1 vccd1 vccd1 OVHB\[18\].V/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_110_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05744__D line[123] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09611_ _09611_/A _09624_/Y vssd1 vssd1 vccd1 vccd1 _13811_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_56_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08120__D line[48] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06823_ _13905_/X wr vssd1 vssd1 vccd1 vccd1 _06823_/X sky130_fd_sc_hd__and2_1
XFILLER_95_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[30\].VALID\[1\].TOBUF OVHB\[30\].VALID\[1\].FF/Q OVHB\[30\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04926_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_37_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06754_ _13905_/X vssd1 vssd1 vccd1 vccd1 _06754_/Y sky130_fd_sc_hd__inv_2
X_09542_ _09550_/CLK line[53] vssd1 vssd1 vccd1 vccd1 _09543_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07314__A _13910_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05705_ _05735_/CLK line[96] vssd1 vssd1 vccd1 vccd1 _05706_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12577__D line[47] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[24\].VALID\[10\].FF OVHB\[24\].V/CLK A[17] vssd1 vssd1 vccd1 vccd1 OVHB\[24\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_09473_ _09473_/A _09484_/Y vssd1 vssd1 vccd1 vccd1 _13673_/Z sky130_fd_sc_hd__ebufn_2
X_06685_ _06715_/CLK line[32] vssd1 vssd1 vccd1 vccd1 _06686_/A sky130_fd_sc_hd__dfxtp_1
XPHY_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05636_ _05636_/A _05669_/Y vssd1 vssd1 vccd1 vccd1 _13756_/Z sky130_fd_sc_hd__ebufn_2
X_08424_ _08430_/CLK line[54] vssd1 vssd1 vccd1 vccd1 _08425_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07033__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06575__D line[105] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08355_ _08355_/A _08364_/Y vssd1 vssd1 vccd1 vccd1 _13675_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05567_ _05595_/CLK line[42] vssd1 vssd1 vccd1 vccd1 _05568_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_211_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09886__D line[82] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07306_ _07310_/CLK line[55] vssd1 vssd1 vccd1 vccd1 _07307_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_165_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08286_ _08290_/CLK line[119] vssd1 vssd1 vccd1 vccd1 _08287_/A sky130_fd_sc_hd__dfxtp_1
X_05498_ _05498_/A _05529_/Y vssd1 vssd1 vccd1 vccd1 _13618_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10825__D line[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07237_ _07237_/A _07244_/Y vssd1 vssd1 vccd1 vccd1 _13677_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_192_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13201__D line[76] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05919__D line[75] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07168_ _07170_/CLK line[120] vssd1 vssd1 vccd1 vccd1 _07169_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[10\].CLKBUF\[2\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06119_ _06119_/A _06124_/Y vssd1 vssd1 vccd1 vccd1 _13679_/Z sky130_fd_sc_hd__ebufn_2
X_07099_ _07099_/A _07104_/Y vssd1 vssd1 vccd1 vccd1 _13819_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_59_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XOVHB\[14\].VALID\[12\].FF OVHB\[14\].V/CLK A[19] vssd1 vssd1 vccd1 vccd1 OVHB\[14\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07208__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09126__D line[119] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09809_ _09809_/A _09834_/Y vssd1 vssd1 vccd1 vccd1 _13729_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_46_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12820_ _12840_/CLK line[30] vssd1 vssd1 vccd1 vccd1 _12821_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_55_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12751_ _12751_/A _12774_/Y vssd1 vssd1 vccd1 vccd1 _13871_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11391__D line[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11702_ _11720_/CLK line[31] vssd1 vssd1 vccd1 vccd1 _11703_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_70_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06485__D line[78] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[3\].CLKBUF\[2\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[22\].VALID\[7\].TOBUF OVHB\[22\].VALID\[7\].FF/Q OVHB\[22\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/A2 sky130_fd_sc_hd__ebufn_2
XPHY_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12682_ _12700_/CLK line[95] vssd1 vssd1 vccd1 vccd1 _12683_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11633_ _11633_/A _11654_/Y vssd1 vssd1 vccd1 vccd1 _13873_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[6\].VALID\[11\].TOBUF OVHB\[6\].VALID\[11\].FF/Q OVHB\[6\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04915_/B2 sky130_fd_sc_hd__ebufn_2
X_11564_ _11580_/CLK line[81] vssd1 vssd1 vccd1 vccd1 _11565_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13303_ _13303_/A _13334_/Y vssd1 vssd1 vccd1 vccd1 _13863_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13896__A A[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10515_ _10515_/A _10534_/Y vssd1 vssd1 vccd1 vccd1 _13875_/Z sky130_fd_sc_hd__ebufn_2
X_11495_ _11495_/A _11514_/Y vssd1 vssd1 vccd1 vccd1 _13735_/Z sky130_fd_sc_hd__ebufn_2
X_10446_ _10460_/CLK line[82] vssd1 vssd1 vccd1 vccd1 _10447_/A sky130_fd_sc_hd__dfxtp_1
X_13234_ _13260_/CLK line[91] vssd1 vssd1 vccd1 vccd1 _13235_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_6_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12950__D line[80] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10377_ _10377_/A _10394_/Y vssd1 vssd1 vccd1 vccd1 _13737_/Z sky130_fd_sc_hd__ebufn_2
X_13165_ _13165_/A _13194_/Y vssd1 vssd1 vccd1 vccd1 _13725_/Z sky130_fd_sc_hd__ebufn_2
X_12116_ _12140_/CLK line[92] vssd1 vssd1 vccd1 vccd1 _12117_/A sky130_fd_sc_hd__dfxtp_1
X_13096_ _13120_/CLK line[28] vssd1 vssd1 vccd1 vccd1 _13097_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_69_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11566__D line[82] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12047_ _12047_/A _12074_/Y vssd1 vssd1 vccd1 vccd1 _13727_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09036__D line[92] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11863__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13781__D line[71] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08875__D line[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12949_ _13937_/X vssd1 vssd1 vccd1 vccd1 _12949_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06470_ _06470_/CLK line[57] vssd1 vssd1 vccd1 vccd1 _06471_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_61_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05421_ _05421_/A _05424_/Y vssd1 vssd1 vccd1 vccd1 _13821_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[13\].VALID\[3\].FF_D A[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08140_ _08150_/CLK line[52] vssd1 vssd1 vccd1 vccd1 _08141_/A sky130_fd_sc_hd__dfxtp_1
X_05352_ _05352_/CLK _05353_/X vssd1 vssd1 vccd1 vccd1 _05350_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_119_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08071_ _08071_/A _08084_/Y vssd1 vssd1 vccd1 vccd1 _13671_/Z sky130_fd_sc_hd__ebufn_2
X_05283_ _13900_/X wr vssd1 vssd1 vccd1 vccd1 _05283_/X sky130_fd_sc_hd__and2_1
XFILLER_146_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07022_ _07030_/CLK line[53] vssd1 vssd1 vccd1 vccd1 _07023_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08115__D line[41] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08973_ _08973_/A _08994_/Y vssd1 vssd1 vccd1 vccd1 _13733_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_29_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10380__D line[52] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07924_ _07940_/CLK line[81] vssd1 vssd1 vccd1 vccd1 _07925_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_68_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05474__D line[113] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07855_ _07855_/A _07874_/Y vssd1 vssd1 vccd1 vccd1 _13735_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_68_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13691__D line[44] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[9\].VALID\[14\].FF OVHB\[9\].V/CLK A[21] vssd1 vssd1 vccd1 vccd1 OVHB\[9\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08785__D line[96] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06806_ _06820_/CLK line[82] vssd1 vssd1 vccd1 vccd1 _06807_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[22\].VALID\[1\].FF OVHB\[22\].V/CLK A[8] vssd1 vssd1 vccd1 vccd1 OVHB\[22\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_45_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_04998_ _05000_/CLK line[24] vssd1 vssd1 vccd1 vccd1 _04999_/A sky130_fd_sc_hd__dfxtp_1
X_07786_ _07800_/CLK line[18] vssd1 vssd1 vccd1 vccd1 _07787_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_56_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09525_ _09525_/A _09554_/Y vssd1 vssd1 vccd1 vccd1 _13725_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_36_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06737_ _06737_/A _06754_/Y vssd1 vssd1 vccd1 vccd1 _13737_/Z sky130_fd_sc_hd__ebufn_2
XPHY_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07979__A _13912_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06668_ _06680_/CLK line[19] vssd1 vssd1 vccd1 vccd1 _06669_/A sky130_fd_sc_hd__dfxtp_1
X_09456_ _09480_/CLK line[28] vssd1 vssd1 vccd1 vccd1 _09457_/A sky130_fd_sc_hd__dfxtp_1
XPHY_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08407_ _08407_/A _08434_/Y vssd1 vssd1 vccd1 vccd1 _13727_/Z sky130_fd_sc_hd__ebufn_2
X_05619_ _05619_/A _05634_/Y vssd1 vssd1 vccd1 vccd1 _13739_/Z sky130_fd_sc_hd__ebufn_2
XPHY_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07698__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09387_ _09387_/A _09414_/Y vssd1 vssd1 vccd1 vccd1 _13867_/Z sky130_fd_sc_hd__ebufn_2
X_06599_ _06599_/A _06614_/Y vssd1 vssd1 vccd1 vccd1 _13879_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[28\].CLKBUF\[5\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08338_ _08360_/CLK line[29] vssd1 vssd1 vccd1 vccd1 _08339_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10555__D line[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08269_ _08269_/A _08294_/Y vssd1 vssd1 vccd1 vccd1 _13869_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05649__D line[65] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10300_ _10320_/CLK line[30] vssd1 vssd1 vccd1 vccd1 _10301_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_165_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08025__D line[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11280_ _11300_/CLK line[94] vssd1 vssd1 vccd1 vccd1 _11281_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[29\].VALID\[13\].TOBUF OVHB\[29\].VALID\[13\].FF/Q OVHB\[29\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04916_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_146_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13866__D line[124] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10231_ _10231_/A _10254_/Y vssd1 vssd1 vccd1 vccd1 _13871_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_10_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12770__D line[121] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07864__D line[54] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10162_ _10180_/CLK line[95] vssd1 vssd1 vccd1 vccd1 _10163_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06123__A _13903_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10290__D line[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10093_ _10093_/A _10114_/Y vssd1 vssd1 vccd1 vccd1 _13733_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_120_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13921_ _13927_/C _13927_/B _13927_/A _13927_/D vssd1 vssd1 vccd1 vccd1 _13921_/X
+ sky130_fd_sc_hd__and4bb_4
XFILLER_19_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13852_ _13852_/A _13859_/Y vssd1 vssd1 vccd1 vccd1 _13852_/Z sky130_fd_sc_hd__ebufn_2
X_12803_ _12805_/CLK line[8] vssd1 vssd1 vccd1 vccd1 _12804_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_62_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__04922__A2 _04922_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13783_ _13785_/CLK line[72] vssd1 vssd1 vccd1 vccd1 _13784_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13106__D line[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10995_ _10995_/A _11024_/Y vssd1 vssd1 vccd1 vccd1 _13795_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_27_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12734_ _12734_/A _12739_/Y vssd1 vssd1 vccd1 vccd1 _13854_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[26\].VALID\[3\].FF_D A[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13403__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12945__D line[73] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[22\].VALID\[12\].TOBUF OVHB\[22\].VALID\[12\].FF/Q OVHB\[22\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04929_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_42_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12665_ _12665_/CLK line[73] vssd1 vssd1 vccd1 vccd1 _12666_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[20\].VALID\[3\].FF OVHB\[20\].V/CLK A[10] vssd1 vssd1 vccd1 vccd1 OVHB\[20\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11616_ _11616_/A _11619_/Y vssd1 vssd1 vccd1 vccd1 _13856_/Z sky130_fd_sc_hd__ebufn_2
XPHY_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12596_ _12596_/A _12599_/Y vssd1 vssd1 vccd1 vccd1 _13716_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_156_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10465__D line[96] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11547_ _11547_/CLK _11548_/X vssd1 vssd1 vccd1 vccd1 _11545_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA_DATA\[1\].CLKBUF\[4\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[10\].VALID\[10\].FF OVHB\[10\].V/CLK A[17] vssd1 vssd1 vccd1 vccd1 OVHB\[10\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[19\].VALID\[7\].FF_D A[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11478_ _13926_/X wr vssd1 vssd1 vccd1 vccd1 _11478_/X sky130_fd_sc_hd__and2_1
XFILLER_109_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12680__D line[94] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13217_ _13225_/CLK line[69] vssd1 vssd1 vccd1 vccd1 _13218_/A sky130_fd_sc_hd__dfxtp_1
X_10429_ _13923_/X vssd1 vssd1 vccd1 vccd1 _10429_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07774__D line[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13148_ _13148_/A _13159_/Y vssd1 vssd1 vccd1 vccd1 _13708_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11296__D line[87] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05970_ _05980_/CLK line[84] vssd1 vssd1 vccd1 vccd1 _05971_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13079_ _13085_/CLK line[6] vssd1 vssd1 vccd1 vccd1 _13080_/A sky130_fd_sc_hd__dfxtp_1
X_04921_ _04920_/Y _04922_/B2 _04918_/Y _04923_/A2 vssd1 vssd1 vccd1 vccd1 _04921_/Y
+ sky130_fd_sc_hd__a22oi_2
XANTENNA__09344__A _13916_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09063__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07640_ _07660_/CLK line[94] vssd1 vssd1 vccd1 vccd1 _07641_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[2\].INV _13977_/X vssd1 vssd1 vccd1 vccd1 OVHB\[2\].INV/Y sky130_fd_sc_hd__inv_2
X_07571_ _07571_/A _07594_/Y vssd1 vssd1 vccd1 vccd1 _13731_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_207_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09310_ _09340_/CLK line[80] vssd1 vssd1 vccd1 vccd1 _09311_/A sky130_fd_sc_hd__dfxtp_1
X_06522_ _06540_/CLK line[95] vssd1 vssd1 vccd1 vccd1 _06523_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_202_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07014__D line[49] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[4\].VALID\[4\].TOBUF OVHB\[4\].VALID\[4\].FF/Q OVHB\[4\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04925_/B2 sky130_fd_sc_hd__ebufn_2
XOVHB\[19\].VALID\[4\].FF OVHB\[19\].V/CLK A[11] vssd1 vssd1 vccd1 vccd1 OVHB\[19\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_06453_ _06453_/A _06474_/Y vssd1 vssd1 vccd1 vccd1 _13733_/Z sky130_fd_sc_hd__ebufn_2
X_09241_ _09241_/A _09274_/Y vssd1 vssd1 vccd1 vccd1 _13721_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12855__D line[46] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[29\].VALID\[7\].TOBUF OVHB\[29\].VALID\[7\].FF/Q OVHB\[29\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/A2 sky130_fd_sc_hd__ebufn_2
X_05404_ _05420_/CLK line[81] vssd1 vssd1 vccd1 vccd1 _05405_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07949__D line[107] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09172_ _09200_/CLK line[26] vssd1 vssd1 vccd1 vccd1 _09173_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06853__D line[104] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06384_ _06400_/CLK line[17] vssd1 vssd1 vccd1 vccd1 _06385_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_178_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08123_ _08123_/A _08154_/Y vssd1 vssd1 vccd1 vccd1 _13723_/Z sky130_fd_sc_hd__ebufn_2
X_05335_ _05335_/A _05354_/Y vssd1 vssd1 vccd1 vccd1 _13735_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10953__A _13925_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08054_ _08080_/CLK line[27] vssd1 vssd1 vccd1 vccd1 _08055_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_135_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05266_ _05280_/CLK line[18] vssd1 vssd1 vccd1 vccd1 _05267_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09519__A _13920_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[23\].CG_CLK clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07005_ _07005_/A _07034_/Y vssd1 vssd1 vccd1 vccd1 _13725_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09238__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05197_ _05197_/A _05214_/Y vssd1 vssd1 vccd1 vccd1 _13877_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_1_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08956_ _08956_/A _08959_/Y vssd1 vssd1 vccd1 vccd1 _13716_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_69_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07907_ _07907_/CLK _07908_/X vssd1 vssd1 vccd1 vccd1 _07905_/CLK sky130_fd_sc_hd__dlclkp_1
X_08887_ _08887_/CLK _08888_/X vssd1 vssd1 vccd1 vccd1 _08885_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_186_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07838_ _13912_/X wr vssd1 vssd1 vccd1 vccd1 _07838_/X sky130_fd_sc_hd__and2_1
XANTENNA__09404__D line[118] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07769_ _13912_/X vssd1 vssd1 vccd1 vccd1 _07769_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09508_ _09508_/A _09519_/Y vssd1 vssd1 vccd1 vccd1 _13708_/Z sky130_fd_sc_hd__ebufn_2
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10780_ _10810_/CLK line[112] vssd1 vssd1 vccd1 vccd1 _10781_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_40_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09439_ _09445_/CLK line[6] vssd1 vssd1 vccd1 vccd1 _09440_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_40_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11024__A _13925_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06763__D line[77] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12450_ _12450_/A _12459_/Y vssd1 vssd1 vccd1 vccd1 _13850_/Z sky130_fd_sc_hd__ebufn_2
X_11401_ _11405_/CLK line[7] vssd1 vssd1 vccd1 vccd1 _11402_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10285__D line[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12381_ _12385_/CLK line[71] vssd1 vssd1 vccd1 vccd1 _12382_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05379__D line[70] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11332_ _11332_/A _11339_/Y vssd1 vssd1 vccd1 vccd1 _13852_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_138_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XOVHB\[17\].VALID\[6\].FF OVHB\[17\].V/CLK A[13] vssd1 vssd1 vccd1 vccd1 OVHB\[17\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13596__D line[114] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[26\].CLKBUF\[7\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11263_ _11265_/CLK line[72] vssd1 vssd1 vccd1 vccd1 _11264_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[5\].VALID\[12\].FF OVHB\[5\].V/CLK A[19] vssd1 vssd1 vccd1 vccd1 OVHB\[5\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_106_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13002_ _13002_/A _13019_/Y vssd1 vssd1 vccd1 vccd1 _13842_/Z sky130_fd_sc_hd__ebufn_2
X_10214_ _10214_/A _10219_/Y vssd1 vssd1 vccd1 vccd1 _13854_/Z sky130_fd_sc_hd__ebufn_2
X_11194_ _11194_/A _11199_/Y vssd1 vssd1 vccd1 vccd1 _13714_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13893__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10145_ _10145_/CLK line[73] vssd1 vssd1 vccd1 vccd1 _10146_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12005__D line[32] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06788__A _13905_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06003__D line[99] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10076_ _10076_/A _10079_/Y vssd1 vssd1 vccd1 vccd1 _13716_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11844__D line[81] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13904_ _13905_/A _13905_/B _13905_/C _13905_/D vssd1 vssd1 vccd1 vccd1 _13904_/X
+ sky130_fd_sc_hd__and4b_4
XANTENNA__06938__D line[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09314__D line[91] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13835_ _13855_/CLK line[110] vssd1 vssd1 vccd1 vccd1 _13836_/A sky130_fd_sc_hd__dfxtp_1
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13766_ _13766_/A _13789_/Y vssd1 vssd1 vccd1 vccd1 _13766_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_15_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10978_ _10978_/A _10989_/Y vssd1 vssd1 vccd1 vccd1 _13778_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_203_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12717_ _12735_/CLK line[111] vssd1 vssd1 vccd1 vccd1 _12718_/A sky130_fd_sc_hd__dfxtp_1
X_13697_ _13715_/CLK line[47] vssd1 vssd1 vccd1 vccd1 _13698_/A sky130_fd_sc_hd__dfxtp_1
XPHY_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12648_ _12648_/A _12669_/Y vssd1 vssd1 vccd1 vccd1 _13768_/Z sky130_fd_sc_hd__ebufn_2
XPHY_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10195__D line[110] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12579_ _12595_/CLK line[33] vssd1 vssd1 vccd1 vccd1 _12580_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_156_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05289__D line[43] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05120_ _05140_/CLK line[94] vssd1 vssd1 vccd1 vccd1 _05121_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_183_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05051_ _05051_/A _05074_/Y vssd1 vssd1 vccd1 vccd1 _13731_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_132_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08810_ _08810_/A _08819_/Y vssd1 vssd1 vccd1 vccd1 _13850_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[2\].VALID\[9\].TOBUF OVHB\[2\].VALID\[9\].FF/Q OVHB\[2\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04914_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[0\].VALID\[11\].FF_D A[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09790_ _09790_/A _09799_/Y vssd1 vssd1 vccd1 vccd1 _13710_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[15\].VALID\[8\].FF OVHB\[15\].V/CLK A[15] vssd1 vssd1 vccd1 vccd1 OVHB\[15\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__04919__A2_N _04919_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[29\].VALID\[10\].FF OVHB\[29\].V/CLK A[17] vssd1 vssd1 vccd1 vccd1 OVHB\[29\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_08741_ _08745_/CLK line[71] vssd1 vssd1 vccd1 vccd1 _08742_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_85_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05953_ _05953_/A _05984_/Y vssd1 vssd1 vccd1 vccd1 _13793_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_38_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05884_ _05910_/CLK line[59] vssd1 vssd1 vccd1 vccd1 _05885_/A sky130_fd_sc_hd__dfxtp_1
X_08672_ _08672_/A _08679_/Y vssd1 vssd1 vccd1 vccd1 _13712_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05752__D line[127] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07623_ _07625_/CLK line[72] vssd1 vssd1 vccd1 vccd1 _07624_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_198_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07554_ _07554_/A _07559_/Y vssd1 vssd1 vccd1 vccd1 _13714_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_22_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06505_ _06505_/CLK line[73] vssd1 vssd1 vccd1 vccd1 _06506_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12585__D line[36] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07485_ _07485_/CLK line[9] vssd1 vssd1 vccd1 vccd1 _07486_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_22_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07679__D line[97] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[16\].CGAND _13909_/Y wr vssd1 vssd1 vccd1 vccd1 OVHB\[16\].CGAND/X sky130_fd_sc_hd__and2_4
X_09224_ _09224_/A _09239_/Y vssd1 vssd1 vccd1 vccd1 _13704_/Z sky130_fd_sc_hd__ebufn_2
X_06436_ _06436_/A _06439_/Y vssd1 vssd1 vccd1 vccd1 _13716_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_158_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06367_ _06367_/CLK _06368_/X vssd1 vssd1 vccd1 vccd1 _06365_/CLK sky130_fd_sc_hd__dlclkp_1
X_09155_ _09165_/CLK line[4] vssd1 vssd1 vccd1 vccd1 _09156_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[0\].CG clk OVHB\[0\].CGAND/X vssd1 vssd1 vccd1 vccd1 OVHB\[0\].V/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__09894__D line[86] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05318_ _13900_/X wr vssd1 vssd1 vccd1 vccd1 _05318_/X sky130_fd_sc_hd__and2_1
X_08106_ _08106_/A _08119_/Y vssd1 vssd1 vccd1 vccd1 _13706_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_190_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08153__A _13932_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09086_ _09086_/A _09099_/Y vssd1 vssd1 vccd1 vccd1 _13846_/Z sky130_fd_sc_hd__ebufn_2
X_06298_ _13903_/X wr vssd1 vssd1 vccd1 vccd1 _06298_/X sky130_fd_sc_hd__and2_1
XOVHB\[19\].VALID\[12\].FF OVHB\[19\].V/CLK A[19] vssd1 vssd1 vccd1 vccd1 OVHB\[19\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_08037_ _08045_/CLK line[5] vssd1 vssd1 vccd1 vccd1 _08038_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10833__D line[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05249_ _13900_/X vssd1 vssd1 vccd1 vccd1 _05249_/Y sky130_fd_sc_hd__inv_2
XFILLER_190_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05927__D line[79] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08303__D line[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09988_ _09988_/A _10009_/Y vssd1 vssd1 vccd1 vccd1 _13628_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_67_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08939_ _08955_/CLK line[33] vssd1 vssd1 vccd1 vccd1 _08940_/A sky130_fd_sc_hd__dfxtp_1
X_11950_ _11950_/A _11969_/Y vssd1 vssd1 vccd1 vccd1 _13630_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_72_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10901_ _10915_/CLK line[34] vssd1 vssd1 vccd1 vccd1 _10902_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.M\[1\].MUX\[0\]_A0 _13644_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[22\].VALID\[6\].FF_D A[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11881_ _11895_/CLK line[98] vssd1 vssd1 vccd1 vccd1 _11882_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_45_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[15\].CGAND_B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13620_ _13620_/A _13649_/Y vssd1 vssd1 vccd1 vccd1 _13620_/Z sky130_fd_sc_hd__ebufn_2
X_10832_ _10832_/A _10849_/Y vssd1 vssd1 vccd1 vccd1 _13632_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08328__A _13913_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13551_ _13575_/CLK line[108] vssd1 vssd1 vccd1 vccd1 _13552_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12495__D line[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10763_ _10775_/CLK line[99] vssd1 vssd1 vccd1 vccd1 _10764_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[19\].CGAND_A _13912_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DECH.DEC0.AND3_B A_h[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12502_ _12502_/A _12529_/Y vssd1 vssd1 vccd1 vccd1 _13622_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06493__D line[67] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13482_ _13482_/A _13509_/Y vssd1 vssd1 vccd1 vccd1 _13762_/Z sky130_fd_sc_hd__ebufn_2
X_10694_ _10694_/A _10709_/Y vssd1 vssd1 vccd1 vccd1 _13774_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11689__A _13927_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12433_ _12455_/CLK line[109] vssd1 vssd1 vccd1 vccd1 _12434_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_172_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XOVHB\[19\].VALID\[11\].TOBUF OVHB\[19\].VALID\[11\].FF/Q OVHB\[19\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04915_/B2 sky130_fd_sc_hd__ebufn_2
X_12364_ _12364_/A _12389_/Y vssd1 vssd1 vccd1 vccd1 _13764_/Z sky130_fd_sc_hd__ebufn_2
X_11315_ _11335_/CLK line[110] vssd1 vssd1 vccd1 vccd1 _11316_/A sky130_fd_sc_hd__dfxtp_1
X_12295_ _12315_/CLK line[46] vssd1 vssd1 vccd1 vccd1 _12296_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_107_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11246_ _11246_/A _11269_/Y vssd1 vssd1 vccd1 vccd1 _13766_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_180_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11177_ _11195_/CLK line[47] vssd1 vssd1 vccd1 vccd1 _11178_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_67_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10128_ _10128_/A _10149_/Y vssd1 vssd1 vccd1 vccd1 _13768_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11574__D line[86] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06668__D line[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10059_ _10075_/CLK line[33] vssd1 vssd1 vccd1 vccd1 _10060_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_48_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09044__D line[81] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_DATA\[20\].CLKBUF\[0\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09979__D line[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08883__D line[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13818_ _13820_/CLK line[88] vssd1 vssd1 vccd1 vccd1 _13819_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[12\].VALID\[10\].TOBUF OVHB\[12\].VALID\[10\].FF/Q OVHB\[12\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04932_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_188_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13749_ _13749_/A _13754_/Y vssd1 vssd1 vccd1 vccd1 _13749_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12983__A _13937_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07270_ _07270_/A _07279_/Y vssd1 vssd1 vccd1 vccd1 _13710_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[1\].VALID\[10\].FF OVHB\[1\].V/CLK A[17] vssd1 vssd1 vccd1 vccd1 OVHB\[1\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_06221_ _06225_/CLK line[71] vssd1 vssd1 vccd1 vccd1 _06222_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[3\].VALID\[1\].FF_D A[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06152_ _06152_/A _06159_/Y vssd1 vssd1 vccd1 vccd1 _13712_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[19\].CLKBUF\[3\] clk vssd1 vssd1 vccd1 vccd1 _07872_/CLK sky130_fd_sc_hd__clkbuf_4
X_05103_ _05105_/CLK line[72] vssd1 vssd1 vccd1 vccd1 _05104_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11749__D line[38] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06083_ _06085_/CLK line[8] vssd1 vssd1 vccd1 vccd1 _06084_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10008__A _13922_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09219__D line[33] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05034_ _05034_/A _05039_/Y vssd1 vssd1 vccd1 vccd1 _13714_/Z sky130_fd_sc_hd__ebufn_2
X_09911_ _09935_/CLK line[108] vssd1 vssd1 vccd1 vccd1 _09912_/A sky130_fd_sc_hd__dfxtp_1
X_09842_ _09842_/A _09869_/Y vssd1 vssd1 vccd1 vccd1 _13762_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_112_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09773_ _09795_/CLK line[45] vssd1 vssd1 vccd1 vccd1 _09774_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11484__D line[59] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06985_ _06995_/CLK line[36] vssd1 vssd1 vccd1 vccd1 _06986_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[8\].VALID\[1\].FF OVHB\[8\].V/CLK A[8] vssd1 vssd1 vccd1 vccd1 OVHB\[8\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_37_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08724_ _08724_/A _08749_/Y vssd1 vssd1 vccd1 vccd1 _13764_/Z sky130_fd_sc_hd__ebufn_2
X_05936_ _05936_/A _05949_/Y vssd1 vssd1 vccd1 vccd1 _13776_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_66_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05482__D line[117] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08655_ _08675_/CLK line[46] vssd1 vssd1 vccd1 vccd1 _08656_/A sky130_fd_sc_hd__dfxtp_1
X_05867_ _05875_/CLK line[37] vssd1 vssd1 vccd1 vccd1 _05868_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_93_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07606_ _07606_/A _07629_/Y vssd1 vssd1 vccd1 vccd1 _13766_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_81_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08793__D line[109] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13054__A _13937_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08586_ _08586_/A _08609_/Y vssd1 vssd1 vccd1 vccd1 _13626_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_53_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05798_ _05798_/A _05809_/Y vssd1 vssd1 vccd1 vccd1 _13638_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07537_ _07555_/CLK line[47] vssd1 vssd1 vccd1 vccd1 _07538_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07468_ _07468_/A _07489_/Y vssd1 vssd1 vccd1 vccd1 _13628_/Z sky130_fd_sc_hd__ebufn_2
X_09207_ _09235_/CLK line[42] vssd1 vssd1 vccd1 vccd1 _09208_/A sky130_fd_sc_hd__dfxtp_1
X_06419_ _06435_/CLK line[33] vssd1 vssd1 vccd1 vccd1 _06420_/A sky130_fd_sc_hd__dfxtp_1
X_07399_ _07415_/CLK line[97] vssd1 vssd1 vccd1 vccd1 _07400_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_5_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09138_ _09138_/A _09169_/Y vssd1 vssd1 vccd1 vccd1 _13618_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_5_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11659__D line[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10563__D line[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09069_ _09095_/CLK line[107] vssd1 vssd1 vccd1 vccd1 _09070_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_163_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05657__D line[69] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11100_ _11100_/A _11129_/Y vssd1 vssd1 vccd1 vccd1 _13620_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08033__D line[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12080_ _12080_/A _12109_/Y vssd1 vssd1 vccd1 vccd1 _13760_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13874__D line[113] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13229__A _13938_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11031_ _11055_/CLK line[108] vssd1 vssd1 vccd1 vccd1 _11032_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[18\].CLKBUF\[0\] clk vssd1 vssd1 vccd1 vccd1 _07487_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__08968__D line[61] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[9\].VALID\[9\].TOBUF OVHB\[9\].VALID\[9\].FF/Q OVHB\[9\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04914_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[7\].VALID\[11\].FF_D A[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[19\].CLKBUF\[1\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05392__D line[90] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12982_ _12982_/CLK _12983_/X vssd1 vssd1 vccd1 vccd1 _12980_/CLK sky130_fd_sc_hd__dlclkp_1
X_11933_ _13927_/X wr vssd1 vssd1 vccd1 vccd1 _11933_/X sky130_fd_sc_hd__and2_1
XFILLER_17_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11864_ _13927_/X vssd1 vssd1 vccd1 vccd1 _11864_/Y sky130_fd_sc_hd__inv_2
XANTENNA_OVHB\[30\].CGAND_A _13926_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13603_ _13603_/A _13614_/Y vssd1 vssd1 vccd1 vccd1 _13883_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_60_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10738__D line[88] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10815_ _10845_/CLK line[0] vssd1 vssd1 vccd1 vccd1 _10816_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[15\].VALID\[10\].FF OVHB\[15\].V/CLK A[17] vssd1 vssd1 vccd1 vccd1 OVHB\[15\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XOVHB\[6\].VALID\[3\].FF OVHB\[6\].V/CLK A[10] vssd1 vssd1 vccd1 vccd1 OVHB\[6\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_11795_ _11825_/CLK line[64] vssd1 vssd1 vccd1 vccd1 _11796_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13114__D line[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13534_ _13540_/CLK line[86] vssd1 vssd1 vccd1 vccd1 _13535_/A sky130_fd_sc_hd__dfxtp_1
X_10746_ _10746_/A _10779_/Y vssd1 vssd1 vccd1 vccd1 _13826_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08208__D line[83] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13465_ _13465_/A _13474_/Y vssd1 vssd1 vccd1 vccd1 _13745_/Z sky130_fd_sc_hd__ebufn_2
X_10677_ _10705_/CLK line[74] vssd1 vssd1 vccd1 vccd1 _10678_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_173_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12416_ _12420_/CLK line[87] vssd1 vssd1 vccd1 vccd1 _12417_/A sky130_fd_sc_hd__dfxtp_1
X_13396_ _13400_/CLK line[23] vssd1 vssd1 vccd1 vccd1 _13397_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10473__D line[109] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12347_ _12347_/A _12354_/Y vssd1 vssd1 vccd1 vccd1 _13747_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05567__D line[42] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[9\].VALID\[5\].FF_D A[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[4\].V_RESET_B rst_n vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12278_ _12280_/CLK line[24] vssd1 vssd1 vccd1 vccd1 _12279_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_4_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11229_ _11229_/A _11234_/Y vssd1 vssd1 vccd1 vccd1 _13749_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07782__D line[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06398__D line[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06770_ _06770_/A _06789_/Y vssd1 vssd1 vccd1 vccd1 _13770_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_82_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05721_ _05735_/CLK line[98] vssd1 vssd1 vccd1 vccd1 _05722_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10498__A _13923_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08440_ _08440_/A _08469_/Y vssd1 vssd1 vccd1 vccd1 _13760_/Z sky130_fd_sc_hd__ebufn_2
X_05652_ _05652_/A _05669_/Y vssd1 vssd1 vccd1 vccd1 _13772_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_91_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05583_ _05595_/CLK line[35] vssd1 vssd1 vccd1 vccd1 _05584_/A sky130_fd_sc_hd__dfxtp_1
X_08371_ _08395_/CLK line[44] vssd1 vssd1 vccd1 vccd1 _08372_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10648__D line[61] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13024__D line[123] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[16\].VALID\[4\].TOBUF OVHB\[16\].VALID\[4\].FF/Q OVHB\[16\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04925_/B2 sky130_fd_sc_hd__ebufn_2
X_07322_ _07322_/A _07349_/Y vssd1 vssd1 vccd1 vccd1 _13762_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_149_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07022__D line[53] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07253_ _07275_/CLK line[45] vssd1 vssd1 vccd1 vccd1 _07254_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12863__D line[35] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07957__D line[111] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06204_ _06204_/A _06229_/Y vssd1 vssd1 vccd1 vccd1 _13764_/Z sky130_fd_sc_hd__ebufn_2
X_07184_ _07184_/A _07209_/Y vssd1 vssd1 vccd1 vccd1 _13624_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_145_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[4\].VALID\[5\].FF OVHB\[4\].V/CLK A[12] vssd1 vssd1 vccd1 vccd1 OVHB\[4\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_06135_ _06155_/CLK line[46] vssd1 vssd1 vccd1 vccd1 _06136_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.M\[3\].MUX\[1\]_A2 _13821_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06066_ _06066_/A _06089_/Y vssd1 vssd1 vccd1 vccd1 _13626_/Z sky130_fd_sc_hd__ebufn_2
X_05017_ _05035_/CLK line[47] vssd1 vssd1 vccd1 vccd1 _05018_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_59_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09825_ _09825_/A _09834_/Y vssd1 vssd1 vccd1 vccd1 _13745_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_86_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12103__D line[72] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09756_ _09760_/CLK line[23] vssd1 vssd1 vccd1 vccd1 _09757_/A sky130_fd_sc_hd__dfxtp_1
X_06968_ _06968_/A _06999_/Y vssd1 vssd1 vccd1 vccd1 _13688_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_64_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08707_ _08707_/A _08714_/Y vssd1 vssd1 vccd1 vccd1 _13747_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_104_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05919_ _05945_/CLK line[75] vssd1 vssd1 vccd1 vccd1 _05920_/A sky130_fd_sc_hd__dfxtp_1
X_09687_ _09687_/A _09694_/Y vssd1 vssd1 vccd1 vccd1 _13887_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_27_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06899_ _06925_/CLK line[11] vssd1 vssd1 vccd1 vccd1 _06900_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08638_ _08640_/CLK line[24] vssd1 vssd1 vccd1 vccd1 _08639_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_54_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08569_ _08569_/A _08574_/Y vssd1 vssd1 vccd1 vccd1 _13889_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10600_ _10600_/CLK line[25] vssd1 vssd1 vccd1 vccd1 _10601_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11580_ _11580_/CLK line[89] vssd1 vssd1 vccd1 vccd1 _11581_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10531_ _10531_/A _10534_/Y vssd1 vssd1 vccd1 vccd1 _13891_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06771__D line[66] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13250_ _13260_/CLK line[84] vssd1 vssd1 vccd1 vccd1 _13251_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_136_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10462_ _10462_/CLK _10463_/X vssd1 vssd1 vccd1 vccd1 _10460_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__11389__D line[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12201_ _12201_/A _12214_/Y vssd1 vssd1 vccd1 vccd1 _13881_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_182_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13181_ _13181_/A _13194_/Y vssd1 vssd1 vccd1 vccd1 _13741_/Z sky130_fd_sc_hd__ebufn_2
X_10393_ _13923_/X wr vssd1 vssd1 vccd1 vccd1 _10393_/X sky130_fd_sc_hd__and2_1
X_12132_ _12140_/CLK line[85] vssd1 vssd1 vccd1 vccd1 _12133_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[22\].VALID\[3\].TOBUF OVHB\[22\].VALID\[3\].FF/Q OVHB\[22\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04919_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__08698__D line[51] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12063_ _12063_/A _12074_/Y vssd1 vssd1 vccd1 vccd1 _13743_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_150_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11014_ _11020_/CLK line[86] vssd1 vssd1 vccd1 vccd1 _11015_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[2\].VALID\[7\].FF OVHB\[2\].V/CLK A[14] vssd1 vssd1 vccd1 vccd1 OVHB\[2\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_131_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12013__D line[45] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07107__D line[106] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06011__D line[103] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12965_ _12965_/A _12984_/Y vssd1 vssd1 vccd1 vccd1 _13805_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11852__D line[85] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11916_ _11930_/CLK line[114] vssd1 vssd1 vccd1 vccd1 _11917_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06946__D line[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12896_ _12910_/CLK line[50] vssd1 vssd1 vccd1 vccd1 _12897_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_205_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09322__D line[95] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11847_ _11847_/A _11864_/Y vssd1 vssd1 vccd1 vccd1 _13807_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_54_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_DATA\[17\].CLKBUF\[3\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11778_ _11790_/CLK line[51] vssd1 vssd1 vccd1 vccd1 _11779_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_41_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13779__D line[70] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13517_ _13517_/A _13544_/Y vssd1 vssd1 vccd1 vccd1 _13797_/Z sky130_fd_sc_hd__ebufn_2
X_10729_ _10729_/A _10744_/Y vssd1 vssd1 vccd1 vccd1 _13809_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12038__A _13934_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13448_ _13470_/CLK line[61] vssd1 vssd1 vccd1 vccd1 _13449_/A sky130_fd_sc_hd__dfxtp_1
X_13379_ _13379_/A _13404_/Y vssd1 vssd1 vccd1 vccd1 _13659_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05297__D line[47] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09037__TE_B _09064_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07940_ _07940_/CLK line[89] vssd1 vssd1 vccd1 vccd1 _07941_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[30\].VALID\[1\].FF OVHB\[30\].V/CLK A[8] vssd1 vssd1 vccd1 vccd1 OVHB\[30\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_130_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_OVHB\[31\].VALID\[9\].FF_D A[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07871_ _07871_/A _07874_/Y vssd1 vssd1 vccd1 vccd1 _13751_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[14\].VALID\[9\].TOBUF OVHB\[14\].VALID\[9\].FF/Q OVHB\[14\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04914_/B2 sky130_fd_sc_hd__ebufn_2
X_09610_ _09620_/CLK line[84] vssd1 vssd1 vccd1 vccd1 _09611_/A sky130_fd_sc_hd__dfxtp_1
X_06822_ _06822_/CLK _06823_/X vssd1 vssd1 vccd1 vccd1 _06820_/CLK sky130_fd_sc_hd__dlclkp_1
X_09541_ _09541_/A _09554_/Y vssd1 vssd1 vccd1 vccd1 _13741_/Z sky130_fd_sc_hd__ebufn_2
X_06753_ _13905_/X wr vssd1 vssd1 vccd1 vccd1 _06753_/X sky130_fd_sc_hd__and2_1
XANTENNA__11762__D line[58] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05704_ _13901_/X vssd1 vssd1 vccd1 vccd1 _05704_/Y sky130_fd_sc_hd__inv_2
X_09472_ _09480_/CLK line[21] vssd1 vssd1 vccd1 vccd1 _09473_/A sky130_fd_sc_hd__dfxtp_1
X_06684_ _13905_/X vssd1 vssd1 vccd1 vccd1 _06684_/Y sky130_fd_sc_hd__inv_2
XANTENNA__05760__D line[116] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[0\].VALID\[9\].FF OVHB\[0\].V/CLK A[16] vssd1 vssd1 vccd1 vccd1 OVHB\[0\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_197_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08423_ _08423_/A _08434_/Y vssd1 vssd1 vccd1 vccd1 _13743_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10378__D line[51] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05635_ _05665_/CLK line[64] vssd1 vssd1 vccd1 vccd1 _05636_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_211_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08354_ _08360_/CLK line[22] vssd1 vssd1 vccd1 vccd1 _08355_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05566_ _05566_/A _05599_/Y vssd1 vssd1 vccd1 vccd1 _13686_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13689__D line[43] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07305_ _07305_/A _07314_/Y vssd1 vssd1 vccd1 vccd1 _13745_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_165_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12593__D line[40] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05497_ _05525_/CLK line[10] vssd1 vssd1 vccd1 vccd1 _05498_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[9\].VALID\[13\].TOBUF OVHB\[9\].VALID\[13\].FF/Q OVHB\[9\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04916_/B2 sky130_fd_sc_hd__ebufn_2
X_08285_ _08285_/A _08294_/Y vssd1 vssd1 vccd1 vccd1 _13885_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07687__D line[101] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07236_ _07240_/CLK line[23] vssd1 vssd1 vccd1 vccd1 _07237_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_166_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07167_ _07167_/A _07174_/Y vssd1 vssd1 vccd1 vccd1 _13887_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11002__D line[95] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06118_ _06120_/CLK line[24] vssd1 vssd1 vccd1 vccd1 _06119_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_59_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XOVHB\[29\].VALID\[2\].FF OVHB\[29\].V/CLK A[9] vssd1 vssd1 vccd1 vccd1 OVHB\[29\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_07098_ _07100_/CLK line[88] vssd1 vssd1 vccd1 vccd1 _07099_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05000__D line[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11937__D line[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[14\].VALID\[1\].FF_D A[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10841__D line[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06049_ _06049_/A _06054_/Y vssd1 vssd1 vccd1 vccd1 _13889_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_160_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05935__D line[68] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MUX.M\[2\].MUX\[2\]_A0 _13667_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08311__D line[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09808_ _09830_/CLK line[61] vssd1 vssd1 vccd1 vccd1 _09809_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_75_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09739_ _09739_/A _09764_/Y vssd1 vssd1 vccd1 vccd1 _13659_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12768__D line[120] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[2\].VALID\[12\].TOBUF OVHB\[2\].VALID\[12\].FF/Q OVHB\[2\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04929_/B2 sky130_fd_sc_hd__ebufn_2
X_12750_ _12770_/CLK line[126] vssd1 vssd1 vccd1 vccd1 _12751_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_15_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05670__D line[80] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11701_ _11701_/A _11724_/Y vssd1 vssd1 vccd1 vccd1 _13661_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12681_ _12681_/A _12704_/Y vssd1 vssd1 vccd1 vccd1 _13801_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_15_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[20\].VALID\[8\].TOBUF OVHB\[20\].VALID\[8\].FF/Q OVHB\[20\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04931_/B2 sky130_fd_sc_hd__ebufn_2
XPHY_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11632_ _11650_/CLK line[127] vssd1 vssd1 vccd1 vccd1 _11633_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11563_ _11563_/A _11584_/Y vssd1 vssd1 vccd1 vccd1 _13803_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07597__D line[74] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13302_ _13330_/CLK line[122] vssd1 vssd1 vccd1 vccd1 _13303_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_7_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10514_ _10530_/CLK line[113] vssd1 vssd1 vccd1 vccd1 _10515_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_11_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11494_ _11510_/CLK line[49] vssd1 vssd1 vccd1 vccd1 _11495_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[5\].VALID\[8\].FF_D A[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13233_ _13233_/A _13264_/Y vssd1 vssd1 vccd1 vccd1 _13793_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_124_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10445_ _10445_/A _10464_/Y vssd1 vssd1 vccd1 vccd1 _13805_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_164_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13164_ _13190_/CLK line[59] vssd1 vssd1 vccd1 vccd1 _13165_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[9\].CLKBUF\[4\] clk vssd1 vssd1 vccd1 vccd1 _13787_/CLK sky130_fd_sc_hd__clkbuf_4
X_10376_ _10390_/CLK line[50] vssd1 vssd1 vccd1 vccd1 _10377_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10751__D line[108] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12115_ _12115_/A _12144_/Y vssd1 vssd1 vccd1 vccd1 _13795_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_112_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13095_ _13095_/A _13124_/Y vssd1 vssd1 vccd1 vccd1 _13655_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05845__D line[32] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12046_ _12070_/CLK line[60] vssd1 vssd1 vccd1 vccd1 _12047_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_37_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XOVHB\[27\].VALID\[4\].FF OVHB\[27\].V/CLK A[11] vssd1 vssd1 vccd1 vccd1 OVHB\[27\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12678__D line[93] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__04925__B1 A_h[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06676__D line[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12948_ _13937_/X wr vssd1 vssd1 vccd1 vccd1 _12948_/X sky130_fd_sc_hd__and2_1
XOVHB\[6\].VALID\[10\].FF OVHB\[6\].V/CLK A[17] vssd1 vssd1 vccd1 vccd1 OVHB\[6\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__09052__D line[85] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12879_ _13937_/X vssd1 vssd1 vccd1 vccd1 _12879_/Y sky130_fd_sc_hd__inv_2
XANTENNA__09987__D line[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[14\].VALID\[13\].FF_D A[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05420_ _05420_/CLK line[89] vssd1 vssd1 vccd1 vccd1 _05421_/A sky130_fd_sc_hd__dfxtp_1
X_05351_ _05351_/A _05354_/Y vssd1 vssd1 vccd1 vccd1 _13751_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10926__D line[60] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13302__D line[122] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08070_ _08080_/CLK line[20] vssd1 vssd1 vccd1 vccd1 _08071_/A sky130_fd_sc_hd__dfxtp_1
X_05282_ _05282_/CLK _05283_/X vssd1 vssd1 vccd1 vccd1 _05280_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__07300__D line[52] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07021_ _07021_/A _07034_/Y vssd1 vssd1 vccd1 vccd1 _13741_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[15\].CLKBUF\[5\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[27\].VALID\[1\].FF_D A[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XOVHB\[4\].VALID\[0\].TOBUF OVHB\[4\].VALID\[0\].FF/Q OVHB\[4\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04924_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[24\].VALID\[12\].FF_D A[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08972_ _08990_/CLK line[63] vssd1 vssd1 vccd1 vccd1 _08973_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_88_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09227__D line[37] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07923_ _07923_/A _07944_/Y vssd1 vssd1 vccd1 vccd1 _13803_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[29\].VALID\[3\].TOBUF OVHB\[29\].VALID\[3\].FF/Q OVHB\[29\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04919_/B2 sky130_fd_sc_hd__ebufn_2
XDATA\[8\].CLKBUF\[1\] clk vssd1 vssd1 vccd1 vccd1 _13402_/CLK sky130_fd_sc_hd__clkbuf_4
X_07854_ _07870_/CLK line[49] vssd1 vssd1 vccd1 vccd1 _07855_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_69_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06805_ _06805_/A _06824_/Y vssd1 vssd1 vccd1 vccd1 _13805_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__04916__B1 A_h[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07785_ _07785_/A _07804_/Y vssd1 vssd1 vccd1 vccd1 _13665_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11492__D line[63] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_04997_ _04997_/A _05004_/Y vssd1 vssd1 vccd1 vccd1 _13677_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_45_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09524_ _09550_/CLK line[59] vssd1 vssd1 vccd1 vccd1 _09525_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_83_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06736_ _06750_/CLK line[50] vssd1 vssd1 vccd1 vccd1 _06737_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06586__D line[124] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05490__D line[121] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_DATA\[8\].CLKBUF\[5\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09455_ _09455_/A _09484_/Y vssd1 vssd1 vccd1 vccd1 _13655_/Z sky130_fd_sc_hd__ebufn_2
XPHY_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06667_ _06667_/A _06684_/Y vssd1 vssd1 vccd1 vccd1 _13667_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_52_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08406_ _08430_/CLK line[60] vssd1 vssd1 vccd1 vccd1 _08407_/A sky130_fd_sc_hd__dfxtp_1
XPHY_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05618_ _05630_/CLK line[51] vssd1 vssd1 vccd1 vccd1 _05619_/A sky130_fd_sc_hd__dfxtp_1
X_09386_ _09410_/CLK line[124] vssd1 vssd1 vccd1 vccd1 _09387_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[25\].VALID\[6\].FF OVHB\[25\].V/CLK A[13] vssd1 vssd1 vccd1 vccd1 OVHB\[25\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XOVHB\[25\].VALID\[14\].TOBUF OVHB\[25\].VALID\[14\].FF/Q OVHB\[25\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_61_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06598_ _06610_/CLK line[115] vssd1 vssd1 vccd1 vccd1 _06599_/A sky130_fd_sc_hd__dfxtp_1
X_08337_ _08337_/A _08364_/Y vssd1 vssd1 vccd1 vccd1 _13657_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_138_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05549_ _05549_/A _05564_/Y vssd1 vssd1 vccd1 vccd1 _13669_/Z sky130_fd_sc_hd__ebufn_2
X_08268_ _08290_/CLK line[125] vssd1 vssd1 vccd1 vccd1 _08269_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07210__D line[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07219_ _07219_/A _07244_/Y vssd1 vssd1 vccd1 vccd1 _13659_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_146_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08199_ _08199_/A _08224_/Y vssd1 vssd1 vccd1 vccd1 _13799_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_193_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10230_ _10250_/CLK line[126] vssd1 vssd1 vccd1 vccd1 _10231_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[28\].CLKBUF\[5\] clk vssd1 vssd1 vccd1 vccd1 _10742_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__06404__A _13904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11667__D line[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10161_ _10161_/A _10184_/Y vssd1 vssd1 vccd1 vccd1 _13801_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06123__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05665__D line[73] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09137__D line[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08041__D line[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10092_ _10110_/CLK line[63] vssd1 vssd1 vccd1 vccd1 _10093_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_120_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13882__D line[117] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13920_ _13927_/A _13927_/B _13927_/C _13927_/D vssd1 vssd1 vccd1 vccd1 _13920_/Y
+ sky130_fd_sc_hd__nor4b_4
XANTENNA__08976__D line[50] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13851_ _13855_/CLK line[103] vssd1 vssd1 vccd1 vccd1 _13852_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_142_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12802_ _12802_/A _12809_/Y vssd1 vssd1 vccd1 vccd1 _13642_/Z sky130_fd_sc_hd__ebufn_2
X_13782_ _13782_/A _13789_/Y vssd1 vssd1 vccd1 vccd1 _13782_/Z sky130_fd_sc_hd__ebufn_2
X_10994_ _11020_/CLK line[91] vssd1 vssd1 vccd1 vccd1 _10995_/A sky130_fd_sc_hd__dfxtp_1
X_12733_ _12735_/CLK line[104] vssd1 vssd1 vccd1 vccd1 _12734_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_15_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12664_ _12664_/A _12669_/Y vssd1 vssd1 vccd1 vccd1 _13784_/Z sky130_fd_sc_hd__ebufn_2
XPHY_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09600__D line[94] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11615_ _11615_/CLK line[105] vssd1 vssd1 vccd1 vccd1 _11616_/A sky130_fd_sc_hd__dfxtp_1
XPHY_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12595_ _12595_/CLK line[41] vssd1 vssd1 vccd1 vccd1 _12596_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11546_ _11546_/A _11549_/Y vssd1 vssd1 vccd1 vccd1 _13786_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08216__D line[87] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11477_ _11477_/CLK _11478_/X vssd1 vssd1 vccd1 vccd1 _11475_/CLK sky130_fd_sc_hd__dlclkp_1
XOVHB\[23\].VALID\[8\].FF OVHB\[23\].V/CLK A[15] vssd1 vssd1 vccd1 vccd1 OVHB\[23\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_13216_ _13216_/A _13229_/Y vssd1 vssd1 vccd1 vccd1 _13776_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_143_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10428_ _13923_/X wr vssd1 vssd1 vccd1 vccd1 _10428_/X sky130_fd_sc_hd__and2_1
XANTENNA__10481__D line[98] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13147_ _13155_/CLK line[37] vssd1 vssd1 vccd1 vccd1 _13148_/A sky130_fd_sc_hd__dfxtp_1
X_10359_ _13923_/X vssd1 vssd1 vccd1 vccd1 _10359_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05575__D line[46] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13078_ _13078_/A _13089_/Y vssd1 vssd1 vccd1 vccd1 _13638_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[27\].CLKBUF\[2\] clk vssd1 vssd1 vccd1 vccd1 _10357_/CLK sky130_fd_sc_hd__clkbuf_4
XMUX.M\[3\].MUX\[3\] _13655_/Z _13725_/Z _13795_/Z _13865_/Z MUX.SEL0BUF\[3\]/X MUX.SEL1BUF\[3\]/X
+ vssd1 vssd1 vccd1 vccd1 Do[27] sky130_fd_sc_hd__mux4_1
XANTENNA__13792__D line[90] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_04920_ A_h[19] vssd1 vssd1 vccd1 vccd1 _04920_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12029_ _12035_/CLK line[38] vssd1 vssd1 vccd1 vccd1 _12030_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07790__D line[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XOVHB\[31\].INV _13971_/X vssd1 vssd1 vccd1 vccd1 OVHB\[31\].INV/Y sky130_fd_sc_hd__inv_2
XFILLER_80_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07570_ _07590_/CLK line[62] vssd1 vssd1 vccd1 vccd1 _07571_/A sky130_fd_sc_hd__dfxtp_1
X_06521_ _06521_/A _06544_/Y vssd1 vssd1 vccd1 vccd1 _13801_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_202_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09240_ _09270_/CLK line[48] vssd1 vssd1 vccd1 vccd1 _09241_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_178_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06452_ _06470_/CLK line[63] vssd1 vssd1 vccd1 vccd1 _06453_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[2\].VALID\[5\].TOBUF OVHB\[2\].VALID\[5\].FF/Q OVHB\[2\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04927_/B2 sky130_fd_sc_hd__ebufn_2
X_05403_ _05403_/A _05424_/Y vssd1 vssd1 vccd1 vccd1 _13803_/Z sky130_fd_sc_hd__ebufn_2
X_09171_ _09171_/A _09204_/Y vssd1 vssd1 vccd1 vccd1 _13651_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10656__D line[50] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06383_ _06383_/A _06404_/Y vssd1 vssd1 vccd1 vccd1 _13663_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13032__D line[127] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[27\].VALID\[8\].TOBUF OVHB\[27\].VALID\[8\].FF/Q OVHB\[27\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04931_/B2 sky130_fd_sc_hd__ebufn_2
X_08122_ _08150_/CLK line[58] vssd1 vssd1 vccd1 vccd1 _08123_/A sky130_fd_sc_hd__dfxtp_1
X_05334_ _05350_/CLK line[49] vssd1 vssd1 vccd1 vccd1 _05335_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08126__D line[60] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07030__D line[57] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10953__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08053_ _08053_/A _08084_/Y vssd1 vssd1 vccd1 vccd1 _13653_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12871__D line[39] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05265_ _05265_/A _05284_/Y vssd1 vssd1 vccd1 vccd1 _13665_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[10\].VALID\[4\].FF_D A[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07965__D line[100] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07004_ _07030_/CLK line[59] vssd1 vssd1 vccd1 vccd1 _07005_/A sky130_fd_sc_hd__dfxtp_1
X_05196_ _05210_/CLK line[114] vssd1 vssd1 vccd1 vccd1 _05197_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_142_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[12\].CGAND _13902_/X wr vssd1 vssd1 vccd1 vccd1 OVHB\[12\].CGAND/X sky130_fd_sc_hd__and2_4
X_08955_ _08955_/CLK line[41] vssd1 vssd1 vccd1 vccd1 _08956_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[13\].CLKBUF\[7\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07906_ _07906_/A _07909_/Y vssd1 vssd1 vccd1 vccd1 _13786_/Z sky130_fd_sc_hd__ebufn_2
X_08886_ _08886_/A _08889_/Y vssd1 vssd1 vccd1 vccd1 _13646_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07837_ _07837_/CLK _07838_/X vssd1 vssd1 vccd1 vccd1 _07835_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__13207__D line[79] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07768_ _13912_/X wr vssd1 vssd1 vccd1 vccd1 _07768_/X sky130_fd_sc_hd__and2_1
XANTENNA__06894__A _13905_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07205__D line[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09507_ _09515_/CLK line[37] vssd1 vssd1 vccd1 vccd1 _09508_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_112_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06719_ _13905_/X vssd1 vssd1 vccd1 vccd1 _06719_/Y sky130_fd_sc_hd__inv_2
XFILLER_197_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07699_ _13911_/X vssd1 vssd1 vccd1 vccd1 _07699_/Y sky130_fd_sc_hd__inv_2
XFILLER_188_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XDATA\[16\].CLKBUF\[5\] clk vssd1 vssd1 vccd1 vccd1 _07102_/CLK sky130_fd_sc_hd__clkbuf_4
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09438_ _09438_/A _09449_/Y vssd1 vssd1 vccd1 vccd1 _13638_/Z sky130_fd_sc_hd__ebufn_2
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMUX.M\[2\].MUX\[5\] _13673_/Z _13743_/Z _13813_/Z _13883_/Z MUX.SEL0BUF\[2\]/X MUX.SEL1BUF\[2\]/X
+ vssd1 vssd1 vccd1 vccd1 Do[21] sky130_fd_sc_hd__mux4_1
XFILLER_200_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09369_ _09375_/CLK line[102] vssd1 vssd1 vccd1 vccd1 _09370_/A sky130_fd_sc_hd__dfxtp_1
X_11400_ _11400_/A _11409_/Y vssd1 vssd1 vccd1 vccd1 _13640_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[6\].CLKBUF\[7\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12380_ _12380_/A _12389_/Y vssd1 vssd1 vccd1 vccd1 _13780_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_122_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12781__D line[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11331_ _11335_/CLK line[103] vssd1 vssd1 vccd1 vccd1 _11332_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_193_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07875__D line[64] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11262_ _11262_/A _11269_/Y vssd1 vssd1 vccd1 vccd1 _13782_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_106_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11397__D line[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13001_ _13015_/CLK line[98] vssd1 vssd1 vccd1 vccd1 _13002_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_4_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10213_ _10215_/CLK line[104] vssd1 vssd1 vccd1 vccd1 _10214_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_106_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11193_ _11195_/CLK line[40] vssd1 vssd1 vccd1 vccd1 _11194_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_121_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10144_ _10144_/A _10149_/Y vssd1 vssd1 vccd1 vccd1 _13784_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06788__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10075_ _10075_/CLK line[41] vssd1 vssd1 vccd1 vccd1 _10076_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_47_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13903_ _13905_/B _13905_/A _13905_/C _13905_/D vssd1 vssd1 vccd1 vccd1 _13903_/X
+ sky130_fd_sc_hd__and4b_4
XFILLER_48_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12021__D line[34] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13834_ _13834_/A _13859_/Y vssd1 vssd1 vccd1 vccd1 _13834_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07115__D line[110] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[30\].VALID\[0\].FF_D A[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13765_ _13785_/CLK line[78] vssd1 vssd1 vccd1 vccd1 _13766_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12956__D line[92] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11860__D line[89] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10977_ _10985_/CLK line[69] vssd1 vssd1 vccd1 vccd1 _10978_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_15_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12716_ _12716_/A _12739_/Y vssd1 vssd1 vccd1 vccd1 _13836_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06954__D line[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13696_ _13696_/A _13719_/Y vssd1 vssd1 vccd1 vccd1 _13696_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09330__D line[84] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05213__A _13931_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12647_ _12665_/CLK line[79] vssd1 vssd1 vccd1 vccd1 _12648_/A sky130_fd_sc_hd__dfxtp_1
XPHY_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XDATA\[15\].CLKBUF\[2\] clk vssd1 vssd1 vccd1 vccd1 _06717_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA_OVHB\[23\].VALID\[4\].FF_D A[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12578_ _12578_/A _12599_/Y vssd1 vssd1 vccd1 vccd1 _13698_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11529_ _11545_/CLK line[65] vssd1 vssd1 vccd1 vccd1 _11530_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_116_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05050_ _05070_/CLK line[62] vssd1 vssd1 vccd1 vccd1 _05051_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_194_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[16\].VALID\[8\].FF_D A[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMUX.M\[1\].MUX\[7\] _13628_/Z _13698_/Z _13768_/Z _13838_/Z MUX.SEL0BUF\[1\]/X MUX.SEL1BUF\[1\]/X
+ vssd1 vssd1 vccd1 vccd1 Do[15] sky130_fd_sc_hd__mux4_1
XFILLER_140_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08740_ _08740_/A _08749_/Y vssd1 vssd1 vccd1 vccd1 _13780_/Z sky130_fd_sc_hd__ebufn_2
X_05952_ _05980_/CLK line[90] vssd1 vssd1 vccd1 vccd1 _05953_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09505__D line[36] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08671_ _08675_/CLK line[39] vssd1 vssd1 vccd1 vccd1 _08672_/A sky130_fd_sc_hd__dfxtp_1
X_05883_ _05883_/A _05914_/Y vssd1 vssd1 vccd1 vccd1 _13723_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_38_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07622_ _07622_/A _07629_/Y vssd1 vssd1 vccd1 vccd1 _13782_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_66_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07553_ _07555_/CLK line[40] vssd1 vssd1 vccd1 vccd1 _07554_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_179_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11770__D line[62] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06504_ _06504_/A _06509_/Y vssd1 vssd1 vccd1 vccd1 _13784_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_179_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06864__D line[123] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07484_ _07484_/A _07489_/Y vssd1 vssd1 vccd1 vccd1 _13644_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_179_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09240__D line[48] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09223_ _09235_/CLK line[35] vssd1 vssd1 vccd1 vccd1 _09224_/A sky130_fd_sc_hd__dfxtp_1
X_06435_ _06435_/CLK line[41] vssd1 vssd1 vccd1 vccd1 _06436_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10386__D line[55] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09154_ _09154_/A _09169_/Y vssd1 vssd1 vccd1 vccd1 _13634_/Z sky130_fd_sc_hd__ebufn_2
X_06366_ _06366_/A _06369_/Y vssd1 vssd1 vccd1 vccd1 _13646_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08434__A _13913_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13697__D line[47] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08105_ _08115_/CLK line[36] vssd1 vssd1 vccd1 vccd1 _08106_/A sky130_fd_sc_hd__dfxtp_1
X_05317_ _05317_/CLK _05318_/X vssd1 vssd1 vccd1 vccd1 _05315_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA_MUX.M\[3\].MUX\[4\]_A0 _13657_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09085_ _09095_/CLK line[100] vssd1 vssd1 vccd1 vccd1 _09086_/A sky130_fd_sc_hd__dfxtp_1
X_06297_ _06297_/CLK _06298_/X vssd1 vssd1 vccd1 vccd1 _06295_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__08153__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07695__D line[105] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XOVHB\[6\].VOBUF OVHB\[6\].V/Q OVHB\[6\].INV/Y vssd1 vssd1 vccd1 vccd1 _04912_/B1
+ sky130_fd_sc_hd__ebufn_2
X_08036_ _08036_/A _08049_/Y vssd1 vssd1 vccd1 vccd1 _13636_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_107_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05248_ _13900_/X wr vssd1 vssd1 vccd1 vccd1 _05248_/X sky130_fd_sc_hd__and2_1
XFILLER_162_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_DATA\[27\].CLKBUF\[1\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11010__D line[84] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05179_ _13931_/Y vssd1 vssd1 vccd1 vccd1 _05179_/Y sky130_fd_sc_hd__inv_2
XANTENNA__06104__D line[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09987_ _10005_/CLK line[15] vssd1 vssd1 vccd1 vccd1 _09988_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_49_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11945__D line[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08938_ _08938_/A _08959_/Y vssd1 vssd1 vccd1 vccd1 _13698_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_76_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05943__D line[72] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09415__D line[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08869_ _08885_/CLK line[1] vssd1 vssd1 vccd1 vccd1 _08870_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_29_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10900_ _10900_/A _10919_/Y vssd1 vssd1 vccd1 vccd1 _13700_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_72_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11880_ _11880_/A _11899_/Y vssd1 vssd1 vccd1 vccd1 _13840_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.M\[1\].MUX\[0\]_A1 _13714_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08609__A _13914_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10831_ _10845_/CLK line[2] vssd1 vssd1 vccd1 vccd1 _10832_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_44_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XOVHB\[15\].VALID\[12\].TOBUF OVHB\[15\].VALID\[12\].FF/Q OVHB\[15\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04929_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__08328__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13550_ _13550_/A _13579_/Y vssd1 vssd1 vccd1 vccd1 _13830_/Z sky130_fd_sc_hd__ebufn_2
X_10762_ _10762_/A _10779_/Y vssd1 vssd1 vccd1 vccd1 _13842_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_12_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12501_ _12525_/CLK line[12] vssd1 vssd1 vccd1 vccd1 _12502_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10296__D line[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[19\].CGAND_B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13481_ _13505_/CLK line[76] vssd1 vssd1 vccd1 vccd1 _13482_/A sky130_fd_sc_hd__dfxtp_1
X_10693_ _10705_/CLK line[67] vssd1 vssd1 vccd1 vccd1 _10694_/A sky130_fd_sc_hd__dfxtp_1
X_12432_ _12432_/A _12459_/Y vssd1 vssd1 vccd1 vccd1 _13832_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_200_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XOVHB\[9\].VALID\[5\].TOBUF OVHB\[9\].VALID\[5\].FF/Q OVHB\[9\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04927_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_166_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12363_ _12385_/CLK line[77] vssd1 vssd1 vccd1 vccd1 _12364_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13400__D line[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11314_ _11314_/A _11339_/Y vssd1 vssd1 vccd1 vccd1 _13834_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_165_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_OVHB\[29\].VALID\[8\].FF_D A[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[3\].V_RESET_B rst_n vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12294_ _12294_/A _12319_/Y vssd1 vssd1 vccd1 vccd1 _13694_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[1\].INV _13976_/X vssd1 vssd1 vccd1 vccd1 OVHB\[1\].INV/Y sky130_fd_sc_hd__inv_2
X_11245_ _11265_/CLK line[78] vssd1 vssd1 vccd1 vccd1 _11246_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_79_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11176_ _11176_/A _11199_/Y vssd1 vssd1 vccd1 vccd1 _13696_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[0\].CLKBUF\[0\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10127_ _10145_/CLK line[79] vssd1 vssd1 vccd1 vccd1 _10128_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_67_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05853__D line[45] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10114__A _13922_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09903__A _13921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10058_ _10058_/A _10079_/Y vssd1 vssd1 vccd1 vccd1 _13698_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12686__D line[82] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13817_ _13817_/A _13824_/Y vssd1 vssd1 vccd1 vccd1 _13817_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_189_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13748_ _13750_/CLK line[56] vssd1 vssd1 vccd1 vccd1 _13749_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09060__D line[89] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12983__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13679_ _13679_/A _13684_/Y vssd1 vssd1 vccd1 vccd1 _13679_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09995__D line[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06220_ _06220_/A _06229_/Y vssd1 vssd1 vccd1 vccd1 _13780_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05878__A _13902_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06151_ _06155_/CLK line[39] vssd1 vssd1 vccd1 vccd1 _06152_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10934__D line[49] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13310__D line[126] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05102_ _05102_/A _05109_/Y vssd1 vssd1 vccd1 vccd1 _13782_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_172_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08404__D line[59] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06082_ _06082_/A _06089_/Y vssd1 vssd1 vccd1 vccd1 _13642_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10008__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05033_ _05035_/CLK line[40] vssd1 vssd1 vccd1 vccd1 _05034_/A sky130_fd_sc_hd__dfxtp_1
X_09910_ _09910_/A _09939_/Y vssd1 vssd1 vccd1 vccd1 _13830_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_144_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09841_ _09865_/CLK line[76] vssd1 vssd1 vccd1 vccd1 _09842_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[16\].VALID\[0\].TOBUF OVHB\[16\].VALID\[0\].FF/Q OVHB\[16\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04924_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_140_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09772_ _09772_/A _09799_/Y vssd1 vssd1 vccd1 vccd1 _13692_/Z sky130_fd_sc_hd__ebufn_2
X_06984_ _06984_/A _06999_/Y vssd1 vssd1 vccd1 vccd1 _13704_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09235__D line[41] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08723_ _08745_/CLK line[77] vssd1 vssd1 vccd1 vccd1 _08724_/A sky130_fd_sc_hd__dfxtp_1
X_05935_ _05945_/CLK line[68] vssd1 vssd1 vccd1 vccd1 _05936_/A sky130_fd_sc_hd__dfxtp_1
X_08654_ _08654_/A _08679_/Y vssd1 vssd1 vccd1 vccd1 _13694_/Z sky130_fd_sc_hd__ebufn_2
X_05866_ _05866_/A _05879_/Y vssd1 vssd1 vccd1 vccd1 _13706_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_93_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07605_ _07625_/CLK line[78] vssd1 vssd1 vccd1 vccd1 _07606_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08585_ _08605_/CLK line[14] vssd1 vssd1 vccd1 vccd1 _08586_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05797_ _05805_/CLK line[5] vssd1 vssd1 vccd1 vccd1 _05798_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_53_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07536_ _07536_/A _07559_/Y vssd1 vssd1 vccd1 vccd1 _13696_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06594__D line[113] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07467_ _07485_/CLK line[15] vssd1 vssd1 vccd1 vccd1 _07468_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_210_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09206_ _09206_/A _09239_/Y vssd1 vssd1 vccd1 vccd1 _13686_/Z sky130_fd_sc_hd__ebufn_2
X_06418_ _06418_/A _06439_/Y vssd1 vssd1 vccd1 vccd1 _13698_/Z sky130_fd_sc_hd__ebufn_2
X_07398_ _07398_/A _07419_/Y vssd1 vssd1 vccd1 vccd1 _13838_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_182_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09137_ _09165_/CLK line[10] vssd1 vssd1 vccd1 vccd1 _09138_/A sky130_fd_sc_hd__dfxtp_1
X_06349_ _06365_/CLK line[1] vssd1 vssd1 vccd1 vccd1 _06350_/A sky130_fd_sc_hd__dfxtp_1
X_09068_ _09068_/A _09099_/Y vssd1 vssd1 vccd1 vccd1 _13828_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_118_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08019_ _08045_/CLK line[11] vssd1 vssd1 vccd1 vccd1 _08020_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_190_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_MUX.SEL0BUF\[3\]_A A[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11030_ _11030_/A _11059_/Y vssd1 vssd1 vccd1 vccd1 _13830_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_150_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11675__D line[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06769__D line[65] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09145__D line[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12981_ _12981_/A _12984_/Y vssd1 vssd1 vccd1 vccd1 _13821_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13890__D line[121] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[25\].CLKBUF\[3\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11932_ _11932_/CLK _11933_/X vssd1 vssd1 vccd1 vccd1 _11930_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08984__D line[54] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07243__A _13910_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11863_ _13927_/X wr vssd1 vssd1 vccd1 vccd1 _11863_/X sky130_fd_sc_hd__and2_1
XANTENNA_OVHB\[30\].CGAND_B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10814_ _13924_/X vssd1 vssd1 vccd1 vccd1 _10814_/Y sky130_fd_sc_hd__inv_2
X_13602_ _13610_/CLK line[117] vssd1 vssd1 vccd1 vccd1 _13603_/A sky130_fd_sc_hd__dfxtp_1
X_11794_ _13927_/X vssd1 vssd1 vccd1 vccd1 _11794_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10745_ _10775_/CLK line[96] vssd1 vssd1 vccd1 vccd1 _10746_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_9_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13533_ _13533_/A _13544_/Y vssd1 vssd1 vccd1 vccd1 _13813_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_43_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13464_ _13470_/CLK line[54] vssd1 vssd1 vccd1 vccd1 _13465_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06009__D line[102] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10676_ _10676_/A _10709_/Y vssd1 vssd1 vccd1 vccd1 _13756_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_186_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12415_ _12415_/A _12424_/Y vssd1 vssd1 vccd1 vccd1 _13815_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_139_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13395_ _13395_/A _13404_/Y vssd1 vssd1 vccd1 vccd1 _13675_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[9\].VALID\[8\].FF OVHB\[9\].V/CLK A[15] vssd1 vssd1 vccd1 vccd1 OVHB\[9\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_154_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12346_ _12350_/CLK line[55] vssd1 vssd1 vccd1 vccd1 _12347_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_154_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12277_ _12277_/A _12284_/Y vssd1 vssd1 vccd1 vccd1 _13677_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_114_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11228_ _11230_/CLK line[56] vssd1 vssd1 vccd1 vccd1 _11229_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07418__A _13910_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11585__D line[96] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11159_ _11159_/A _11164_/Y vssd1 vssd1 vccd1 vccd1 _13679_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_122_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05583__D line[35] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_OVHB\[1\].VALID\[12\].FF_D A[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10779__A _13924_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05720_ _05720_/A _05739_/Y vssd1 vssd1 vccd1 vccd1 _13840_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08894__D line[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10498__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05651_ _05665_/CLK line[66] vssd1 vssd1 vccd1 vccd1 _05652_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08370_ _08370_/A _08399_/Y vssd1 vssd1 vccd1 vccd1 _13690_/Z sky130_fd_sc_hd__ebufn_2
X_05582_ _05582_/A _05599_/Y vssd1 vssd1 vccd1 vccd1 _13702_/Z sky130_fd_sc_hd__ebufn_2
X_07321_ _07345_/CLK line[76] vssd1 vssd1 vccd1 vccd1 _07322_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_204_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XDATA\[6\].CLKBUF\[6\] clk vssd1 vssd1 vccd1 vccd1 _13017_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_149_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XOVHB\[14\].VALID\[5\].TOBUF OVHB\[14\].VALID\[5\].FF/Q OVHB\[14\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04927_/B2 sky130_fd_sc_hd__ebufn_2
X_07252_ _07252_/A _07279_/Y vssd1 vssd1 vccd1 vccd1 _13692_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_137_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06203_ _06225_/CLK line[77] vssd1 vssd1 vccd1 vccd1 _06204_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10664__D line[54] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07183_ _07205_/CLK line[13] vssd1 vssd1 vccd1 vccd1 _07184_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13040__D line[116] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05758__D line[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06134_ _06134_/A _06159_/Y vssd1 vssd1 vccd1 vccd1 _13694_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08134__D line[49] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MUX.M\[3\].MUX\[1\]_A3 _13891_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06065_ _06085_/CLK line[14] vssd1 vssd1 vccd1 vccd1 _06066_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_99_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07973__D line[104] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[0\].VALID\[2\].FF_D A[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05016_ _05016_/A _05039_/Y vssd1 vssd1 vccd1 vccd1 _13696_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_98_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09824_ _09830_/CLK line[54] vssd1 vssd1 vccd1 vccd1 _09825_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_100_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09755_ _09755_/A _09764_/Y vssd1 vssd1 vccd1 vccd1 _13675_/Z sky130_fd_sc_hd__ebufn_2
X_06967_ _06995_/CLK line[42] vssd1 vssd1 vccd1 vccd1 _06968_/A sky130_fd_sc_hd__dfxtp_1
X_08706_ _08710_/CLK line[55] vssd1 vssd1 vccd1 vccd1 _08707_/A sky130_fd_sc_hd__dfxtp_1
X_05918_ _05918_/A _05949_/Y vssd1 vssd1 vccd1 vccd1 _13758_/Z sky130_fd_sc_hd__ebufn_2
X_09686_ _09690_/CLK line[119] vssd1 vssd1 vccd1 vccd1 _09687_/A sky130_fd_sc_hd__dfxtp_1
X_06898_ _06898_/A _06929_/Y vssd1 vssd1 vccd1 vccd1 _13618_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08637_ _08637_/A _08644_/Y vssd1 vssd1 vccd1 vccd1 _13677_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10839__D line[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05849_ _05875_/CLK line[43] vssd1 vssd1 vccd1 vccd1 _05850_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13215__D line[68] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08309__D line[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08568_ _08570_/CLK line[120] vssd1 vssd1 vccd1 vccd1 _08569_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07519_ _07519_/A _07524_/Y vssd1 vssd1 vccd1 vccd1 _13679_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_80_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08499_ _08499_/A _08504_/Y vssd1 vssd1 vccd1 vccd1 _13819_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10530_ _10530_/CLK line[121] vssd1 vssd1 vccd1 vccd1 _10531_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10574__D line[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10461_ _10461_/A _10464_/Y vssd1 vssd1 vccd1 vccd1 _13821_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_6_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12200_ _12210_/CLK line[116] vssd1 vssd1 vccd1 vccd1 _12201_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[5\].CLKBUF\[3\] clk vssd1 vssd1 vccd1 vccd1 _12632_/CLK sky130_fd_sc_hd__clkbuf_4
X_13180_ _13190_/CLK line[52] vssd1 vssd1 vccd1 vccd1 _13181_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_202_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10392_ _10392_/CLK _10393_/X vssd1 vssd1 vccd1 vccd1 _10390_/CLK sky130_fd_sc_hd__dlclkp_1
XOVHB\[18\].VALID\[0\].FF OVHB\[18\].V/CLK A[7] vssd1 vssd1 vccd1 vccd1 OVHB\[18\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_12131_ _12131_/A _12144_/Y vssd1 vssd1 vccd1 vccd1 _13811_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12144__A _13934_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07883__D line[77] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12062_ _12070_/CLK line[53] vssd1 vssd1 vccd1 vccd1 _12063_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[20\].VALID\[4\].TOBUF OVHB\[20\].VALID\[4\].FF/Q OVHB\[20\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04925_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_2_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11013_ _11013_/A _11024_/Y vssd1 vssd1 vccd1 vccd1 _13813_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_1_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06499__D line[70] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12964_ _12980_/CLK line[81] vssd1 vssd1 vccd1 vccd1 _12965_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10749__D line[107] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11915_ _11915_/A _11934_/Y vssd1 vssd1 vccd1 vccd1 _13875_/Z sky130_fd_sc_hd__ebufn_2
X_12895_ _12895_/A _12914_/Y vssd1 vssd1 vccd1 vccd1 _13735_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13125__D line[32] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11846_ _11860_/CLK line[82] vssd1 vssd1 vccd1 vccd1 _11847_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07123__D line[99] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDATA\[25\].CLKBUF\[7\] clk vssd1 vssd1 vccd1 vccd1 _09972_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA_DATA\[23\].CLKBUF\[5\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12964__D line[81] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11777_ _11777_/A _11794_/Y vssd1 vssd1 vccd1 vccd1 _13737_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_14_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12319__A _13935_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10728_ _10740_/CLK line[83] vssd1 vssd1 vccd1 vccd1 _10729_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_13_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13516_ _13540_/CLK line[92] vssd1 vssd1 vccd1 vccd1 _13517_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_159_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12038__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13447_ _13447_/A _13474_/Y vssd1 vssd1 vccd1 vccd1 _13727_/Z sky130_fd_sc_hd__ebufn_2
X_10659_ _10659_/A _10674_/Y vssd1 vssd1 vccd1 vccd1 _13739_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_173_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13378_ _13400_/CLK line[29] vssd1 vssd1 vccd1 vccd1 _13379_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_154_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12329_ _12329_/A _12354_/Y vssd1 vssd1 vccd1 vccd1 _13729_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_142_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XDATA\[4\].CLKBUF\[0\] clk vssd1 vssd1 vccd1 vccd1 _12247_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_68_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12204__D line[118] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07870_ _07870_/CLK line[57] vssd1 vssd1 vccd1 vccd1 _07871_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_68_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_OVHB\[6\].VALID\[6\].FF_D A[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06821_ _06821_/A _06824_/Y vssd1 vssd1 vccd1 vccd1 _13821_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[16\].VALID\[2\].FF OVHB\[16\].V/CLK A[9] vssd1 vssd1 vccd1 vccd1 OVHB\[16\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09540_ _09550_/CLK line[52] vssd1 vssd1 vccd1 vccd1 _09541_/A sky130_fd_sc_hd__dfxtp_1
X_06752_ _06752_/CLK _06753_/X vssd1 vssd1 vccd1 vccd1 _06750_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_209_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09513__D line[40] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05703_ _13901_/X wr vssd1 vssd1 vccd1 vccd1 _05703_/X sky130_fd_sc_hd__and2_1
X_09471_ _09471_/A _09484_/Y vssd1 vssd1 vccd1 vccd1 _13671_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[5\].VALID\[14\].TOBUF OVHB\[5\].VALID\[14\].FF/Q OVHB\[5\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/B2 sky130_fd_sc_hd__ebufn_2
X_06683_ _13905_/X wr vssd1 vssd1 vccd1 vccd1 _06683_/X sky130_fd_sc_hd__and2_1
X_08422_ _08430_/CLK line[53] vssd1 vssd1 vccd1 vccd1 _08423_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13613__A _13898_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05634_ _13901_/X vssd1 vssd1 vccd1 vccd1 _05634_/Y sky130_fd_sc_hd__inv_2
XANTENNA_OVHB\[17\].CG_CLK clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08353_ _08353_/A _08364_/Y vssd1 vssd1 vccd1 vccd1 _13673_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[9\].V OVHB\[9\].V/CLK TIE/HI rst_n vssd1 vssd1 vccd1 vccd1 OVHB\[9\].V/Q sky130_fd_sc_hd__dfrtp_1
XPHY_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05565_ _05595_/CLK line[32] vssd1 vssd1 vccd1 vccd1 _05566_/A sky130_fd_sc_hd__dfxtp_1
X_07304_ _07310_/CLK line[54] vssd1 vssd1 vccd1 vccd1 _07305_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06872__D line[127] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08284_ _08290_/CLK line[118] vssd1 vssd1 vccd1 vccd1 _08285_/A sky130_fd_sc_hd__dfxtp_1
X_05496_ _05496_/A _05529_/Y vssd1 vssd1 vccd1 vccd1 _13616_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_164_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07235_ _07235_/A _07244_/Y vssd1 vssd1 vccd1 vccd1 _13675_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[24\].CLKBUF\[4\] clk vssd1 vssd1 vccd1 vccd1 _09587_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__05488__D line[120] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07166_ _07170_/CLK line[119] vssd1 vssd1 vccd1 vccd1 _07167_/A sky130_fd_sc_hd__dfxtp_1
X_06117_ _06117_/A _06124_/Y vssd1 vssd1 vccd1 vccd1 _13677_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08799__D line[97] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07097_ _07097_/A _07104_/Y vssd1 vssd1 vccd1 vccd1 _13817_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_59_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06048_ _06050_/CLK line[120] vssd1 vssd1 vccd1 vccd1 _06049_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_133_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XOVHB\[25\].VALID\[10\].TOBUF OVHB\[25\].VALID\[10\].FF/Q OVHB\[25\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04932_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.M\[2\].MUX\[2\]_A1 _13737_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12114__D line[91] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09273__A _13916_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06112__D line[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09807_ _09807_/A _09834_/Y vssd1 vssd1 vccd1 vccd1 _13727_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_115_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07999_ _07999_/A _08014_/Y vssd1 vssd1 vccd1 vccd1 _13879_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11953__D line[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09738_ _09760_/CLK line[29] vssd1 vssd1 vccd1 vccd1 _09739_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09423__D line[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_OVHB\[8\].VALID\[12\].FF_D A[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_199_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09669_ _09669_/A _09694_/Y vssd1 vssd1 vccd1 vccd1 _13869_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11700_ _11720_/CLK line[30] vssd1 vssd1 vccd1 vccd1 _11701_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_27_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12680_ _12700_/CLK line[94] vssd1 vssd1 vccd1 vccd1 _12681_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08039__D line[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[14\].VALID\[4\].FF OVHB\[14\].V/CLK A[11] vssd1 vssd1 vccd1 vccd1 OVHB\[14\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11631_ _11631_/A _11654_/Y vssd1 vssd1 vccd1 vccd1 _13871_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_70_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[31\].VALID\[8\].FF OVHB\[31\].V/CLK A[15] vssd1 vssd1 vccd1 vccd1 OVHB\[31\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11562_ _11580_/CLK line[95] vssd1 vssd1 vccd1 vccd1 _11563_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10513_ _10513_/A _10534_/Y vssd1 vssd1 vccd1 vccd1 _13873_/Z sky130_fd_sc_hd__ebufn_2
X_13301_ _13301_/A _13334_/Y vssd1 vssd1 vccd1 vccd1 _13861_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11493_ _11493_/A _11514_/Y vssd1 vssd1 vccd1 vccd1 _13733_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05398__D line[93] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13232_ _13260_/CLK line[90] vssd1 vssd1 vccd1 vccd1 _13233_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09448__A _13920_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10444_ _10460_/CLK line[81] vssd1 vssd1 vccd1 vccd1 _10445_/A sky130_fd_sc_hd__dfxtp_1
X_13163_ _13163_/A _13194_/Y vssd1 vssd1 vccd1 vccd1 _13723_/Z sky130_fd_sc_hd__ebufn_2
X_10375_ _10375_/A _10394_/Y vssd1 vssd1 vccd1 vccd1 _13735_/Z sky130_fd_sc_hd__ebufn_2
X_12114_ _12140_/CLK line[91] vssd1 vssd1 vccd1 vccd1 _12115_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[23\].CLKBUF\[1\] clk vssd1 vssd1 vccd1 vccd1 _09202_/CLK sky130_fd_sc_hd__clkbuf_4
X_13094_ _13120_/CLK line[27] vssd1 vssd1 vccd1 vccd1 _13095_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_111_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12045_ _12045_/A _12074_/Y vssd1 vssd1 vccd1 vccd1 _13725_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_49_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XOVHB\[23\].V OVHB\[23\].V/CLK TIE/HI rst_n vssd1 vssd1 vccd1 vccd1 OVHB\[23\].V/Q
+ sky130_fd_sc_hd__dfrtp_1
XDATA\[13\].CLKBUF\[7\] clk vssd1 vssd1 vccd1 vccd1 _06332_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__06022__D line[122] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__04925__B2 _04925_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05861__D line[34] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10479__D line[97] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12947_ _12947_/CLK _12948_/X vssd1 vssd1 vccd1 vccd1 _12945_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_65_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12878_ _13937_/X wr vssd1 vssd1 vccd1 vccd1 _12878_/X sky130_fd_sc_hd__and2_1
XANTENNA__12694__D line[86] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11829_ _13927_/X vssd1 vssd1 vccd1 vccd1 _11829_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07788__D line[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05350_ _05350_/CLK line[57] vssd1 vssd1 vccd1 vccd1 _05351_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_186_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05281_ _05281_/A _05284_/Y vssd1 vssd1 vccd1 vccd1 _13681_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11103__D line[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07020_ _07030_/CLK line[52] vssd1 vssd1 vccd1 vccd1 _07021_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[12\].VALID\[6\].FF OVHB\[12\].V/CLK A[13] vssd1 vssd1 vccd1 vccd1 OVHB\[12\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__05101__D line[71] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[21\].CLKBUF\[7\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10942__D line[53] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08412__D line[63] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08971_ _08971_/A _08994_/Y vssd1 vssd1 vccd1 vccd1 _13731_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_102_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XOVHB\[2\].VALID\[1\].TOBUF OVHB\[2\].VALID\[1\].FF/Q OVHB\[2\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04926_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_114_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07922_ _07940_/CLK line[95] vssd1 vssd1 vccd1 vccd1 _07923_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[14\].V OVHB\[14\].V/CLK TIE/HI rst_n vssd1 vssd1 vccd1 vccd1 OVHB\[14\].V/Q
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07028__D line[56] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[27\].VALID\[4\].TOBUF OVHB\[27\].VALID\[4\].FF/Q OVHB\[27\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04925_/B2 sky130_fd_sc_hd__ebufn_2
X_07853_ _07853_/A _07874_/Y vssd1 vssd1 vccd1 vccd1 _13733_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12869__D line[38] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11128__A _13933_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06804_ _06820_/CLK line[81] vssd1 vssd1 vccd1 vccd1 _06805_/A sky130_fd_sc_hd__dfxtp_1
X_07784_ _07800_/CLK line[17] vssd1 vssd1 vccd1 vccd1 _07785_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__04916__B2 _04916_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_04996_ _05000_/CLK line[23] vssd1 vssd1 vccd1 vccd1 _04997_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[12\].CLKBUF\[4\] clk vssd1 vssd1 vccd1 vccd1 _05947_/CLK sky130_fd_sc_hd__clkbuf_4
X_09523_ _09523_/A _09554_/Y vssd1 vssd1 vccd1 vccd1 _13723_/Z sky130_fd_sc_hd__ebufn_2
X_06735_ _06735_/A _06754_/Y vssd1 vssd1 vccd1 vccd1 _13735_/Z sky130_fd_sc_hd__ebufn_2
X_09454_ _09480_/CLK line[27] vssd1 vssd1 vccd1 vccd1 _09455_/A sky130_fd_sc_hd__dfxtp_1
X_06666_ _06680_/CLK line[18] vssd1 vssd1 vccd1 vccd1 _06667_/A sky130_fd_sc_hd__dfxtp_1
XPHY_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08405_ _08405_/A _08434_/Y vssd1 vssd1 vccd1 vccd1 _13725_/Z sky130_fd_sc_hd__ebufn_2
X_05617_ _05617_/A _05634_/Y vssd1 vssd1 vccd1 vccd1 _13737_/Z sky130_fd_sc_hd__ebufn_2
X_09385_ _09385_/A _09414_/Y vssd1 vssd1 vccd1 vccd1 _13865_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_169_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06597_ _06597_/A _06614_/Y vssd1 vssd1 vccd1 vccd1 _13877_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_178_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08336_ _08360_/CLK line[28] vssd1 vssd1 vccd1 vccd1 _08337_/A sky130_fd_sc_hd__dfxtp_1
X_05548_ _05560_/CLK line[19] vssd1 vssd1 vccd1 vccd1 _05549_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_177_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08267_ _08267_/A _08294_/Y vssd1 vssd1 vccd1 vccd1 _13867_/Z sky130_fd_sc_hd__ebufn_2
X_05479_ _05479_/A _05494_/Y vssd1 vssd1 vccd1 vccd1 _13879_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_20_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07218_ _07240_/CLK line[29] vssd1 vssd1 vccd1 vccd1 _07219_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_125_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08198_ _08220_/CLK line[93] vssd1 vssd1 vccd1 vccd1 _08199_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_180_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05011__D line[44] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07149_ _07149_/A _07174_/Y vssd1 vssd1 vccd1 vccd1 _13869_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10852__D line[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10160_ _10180_/CLK line[94] vssd1 vssd1 vccd1 vccd1 _10161_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_121_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10091_ _10091_/A _10114_/Y vssd1 vssd1 vccd1 vccd1 _13731_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_126_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XOVHB\[10\].VALID\[8\].FF OVHB\[10\].V/CLK A[15] vssd1 vssd1 vccd1 vccd1 OVHB\[10\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_47_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12779__D line[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11683__D line[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[11\].VALID\[2\].FF_D A[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06777__D line[69] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13850_ _13850_/A _13859_/Y vssd1 vssd1 vccd1 vccd1 _13850_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09153__D line[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12801_ _12805_/CLK line[7] vssd1 vssd1 vccd1 vccd1 _12802_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_90_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13781_ _13785_/CLK line[71] vssd1 vssd1 vccd1 vccd1 _13782_/A sky130_fd_sc_hd__dfxtp_1
X_10993_ _10993_/A _11024_/Y vssd1 vssd1 vccd1 vccd1 _13793_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_203_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12732_ _12732_/A _12739_/Y vssd1 vssd1 vccd1 vccd1 _13852_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_35_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12663_ _12665_/CLK line[72] vssd1 vssd1 vccd1 vccd1 _12664_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XDATA\[11\].CLKBUF\[1\] clk vssd1 vssd1 vccd1 vccd1 _05562_/CLK sky130_fd_sc_hd__clkbuf_4
XPHY_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11614_ _11614_/A _11619_/Y vssd1 vssd1 vccd1 vccd1 _13854_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12594_ _12594_/A _12599_/Y vssd1 vssd1 vccd1 vccd1 _13714_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07401__D line[98] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12019__D line[33] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11545_ _11545_/CLK line[73] vssd1 vssd1 vccd1 vccd1 _11546_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11476_ _11476_/A _11479_/Y vssd1 vssd1 vccd1 vccd1 _13716_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11858__D line[88] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10427_ _10427_/CLK _10428_/X vssd1 vssd1 vccd1 vccd1 _10425_/CLK sky130_fd_sc_hd__dlclkp_1
X_13215_ _13225_/CLK line[68] vssd1 vssd1 vccd1 vccd1 _13216_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09328__D line[83] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10358_ _13923_/X wr vssd1 vssd1 vccd1 vccd1 _10358_/X sky130_fd_sc_hd__and2_1
X_13146_ _13146_/A _13159_/Y vssd1 vssd1 vccd1 vccd1 _13706_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[2\].VALID\[9\].FF_D A[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13077_ _13085_/CLK line[5] vssd1 vssd1 vccd1 vccd1 _13078_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[10\].VALID\[10\].FF_D A[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10289_ _13923_/X vssd1 vssd1 vccd1 vccd1 _10289_/Y sky130_fd_sc_hd__inv_2
X_12028_ _12028_/A _12039_/Y vssd1 vssd1 vccd1 vccd1 _13708_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_111_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11593__D line[109] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06687__D line[42] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05591__D line[39] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13979_ _13982_/A _13982_/B _13982_/C _13982_/D vssd1 vssd1 vccd1 vccd1 _13979_/X
+ sky130_fd_sc_hd__and4bb_4
X_06520_ _06540_/CLK line[94] vssd1 vssd1 vccd1 vccd1 _06521_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_34_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06451_ _06451_/A _06474_/Y vssd1 vssd1 vccd1 vccd1 _13731_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_21_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05402_ _05420_/CLK line[95] vssd1 vssd1 vccd1 vccd1 _05403_/A sky130_fd_sc_hd__dfxtp_1
X_09170_ _09200_/CLK line[16] vssd1 vssd1 vccd1 vccd1 _09171_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__04935__D line[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[0\].VALID\[6\].TOBUF OVHB\[0\].VALID\[6\].FF/Q OVHB\[0\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04923_/A2 sky130_fd_sc_hd__ebufn_2
X_06382_ _06400_/CLK line[31] vssd1 vssd1 vccd1 vccd1 _06383_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_147_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08121_ _08121_/A _08154_/Y vssd1 vssd1 vccd1 vccd1 _13721_/Z sky130_fd_sc_hd__ebufn_2
X_05333_ _05333_/A _05354_/Y vssd1 vssd1 vccd1 vccd1 _13733_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[25\].VALID\[9\].TOBUF OVHB\[25\].VALID\[9\].FF/Q OVHB\[25\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04914_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_186_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08052_ _08080_/CLK line[26] vssd1 vssd1 vccd1 vccd1 _08053_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_107_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05264_ _05280_/CLK line[17] vssd1 vssd1 vccd1 vccd1 _05265_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11768__D line[61] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07003_ _07003_/A _07034_/Y vssd1 vssd1 vccd1 vccd1 _13723_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_143_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05195_ _05195_/A _05214_/Y vssd1 vssd1 vccd1 vccd1 _13875_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05766__D line[119] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08142__D line[53] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[24\].VALID\[2\].FF_D A[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08954_ _08954_/A _08959_/Y vssd1 vssd1 vccd1 vccd1 _13714_/Z sky130_fd_sc_hd__ebufn_2
X_07905_ _07905_/CLK line[73] vssd1 vssd1 vccd1 vccd1 _07906_/A sky130_fd_sc_hd__dfxtp_1
X_08885_ _08885_/CLK line[9] vssd1 vssd1 vccd1 vccd1 _08886_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_56_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07836_ _07836_/A _07839_/Y vssd1 vssd1 vccd1 vccd1 _13716_/Z sky130_fd_sc_hd__ebufn_2
X_04979_ _04979_/A _05004_/Y vssd1 vssd1 vccd1 vccd1 _13659_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_37_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07767_ _07767_/CLK _07768_/X vssd1 vssd1 vccd1 vccd1 _07765_/CLK sky130_fd_sc_hd__dlclkp_1
XOVHB\[2\].VOBUF OVHB\[2\].V/Q OVHB\[2\].INV/Y vssd1 vssd1 vccd1 vccd1 _04912_/B1
+ sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[17\].VALID\[6\].FF_D A[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11008__D line[83] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09506_ _09506_/A _09519_/Y vssd1 vssd1 vccd1 vccd1 _13706_/Z sky130_fd_sc_hd__ebufn_2
X_06718_ _13905_/X wr vssd1 vssd1 vccd1 vccd1 _06718_/X sky130_fd_sc_hd__and2_1
XFILLER_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07698_ _13911_/X wr vssd1 vssd1 vccd1 vccd1 _07698_/X sky130_fd_sc_hd__and2_1
XANTENNA__09701__D line[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09437_ _09445_/CLK line[5] vssd1 vssd1 vccd1 vccd1 _09438_/A sky130_fd_sc_hd__dfxtp_1
X_06649_ _13905_/X vssd1 vssd1 vccd1 vccd1 _06649_/Y sky130_fd_sc_hd__inv_2
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13223__D line[72] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08317__D line[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09368_ _09368_/A _09379_/Y vssd1 vssd1 vccd1 vccd1 _13848_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_178_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08319_ _08325_/CLK line[6] vssd1 vssd1 vccd1 vccd1 _08320_/A sky130_fd_sc_hd__dfxtp_1
X_09299_ _09305_/CLK line[70] vssd1 vssd1 vccd1 vccd1 _09300_/A sky130_fd_sc_hd__dfxtp_1
X_11330_ _11330_/A _11339_/Y vssd1 vssd1 vccd1 vccd1 _13850_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_115_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[2\].V_RESET_B rst_n vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10582__D line[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11261_ _11265_/CLK line[71] vssd1 vssd1 vccd1 vccd1 _11262_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_180_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05676__D line[92] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13000_ _13000_/A _13019_/Y vssd1 vssd1 vccd1 vccd1 _13840_/Z sky130_fd_sc_hd__ebufn_2
X_10212_ _10212_/A _10219_/Y vssd1 vssd1 vccd1 vccd1 _13852_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08052__D line[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11192_ _11192_/A _11199_/Y vssd1 vssd1 vccd1 vccd1 _13712_/Z sky130_fd_sc_hd__ebufn_2
X_10143_ _10145_/CLK line[72] vssd1 vssd1 vccd1 vccd1 _10144_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07891__D line[66] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[31\].VALID\[8\].TOBUF OVHB\[31\].VALID\[8\].FF/Q OVHB\[31\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04931_/B2 sky130_fd_sc_hd__ebufn_2
X_10074_ _10074_/A _10079_/Y vssd1 vssd1 vccd1 vccd1 _13714_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[3\].VALID\[1\].FF OVHB\[3\].V/CLK A[8] vssd1 vssd1 vccd1 vccd1 OVHB\[3\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XOVHB\[9\].VALID\[1\].TOBUF OVHB\[9\].VALID\[1\].FF/Q OVHB\[9\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04926_/B2 sky130_fd_sc_hd__ebufn_2
X_13902_ _13905_/A _13905_/B _13905_/C _13905_/D vssd1 vssd1 vccd1 vccd1 _13902_/X
+ sky130_fd_sc_hd__and4bb_4
XFILLER_101_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06300__D line[112] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13833_ _13855_/CLK line[109] vssd1 vssd1 vccd1 vccd1 _13834_/A sky130_fd_sc_hd__dfxtp_1
X_13764_ _13764_/A _13789_/Y vssd1 vssd1 vccd1 vccd1 _13764_/Z sky130_fd_sc_hd__ebufn_2
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10976_ _10976_/A _10989_/Y vssd1 vssd1 vccd1 vccd1 _13776_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10757__D line[111] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12715_ _12735_/CLK line[110] vssd1 vssd1 vccd1 vccd1 _12716_/A sky130_fd_sc_hd__dfxtp_1
X_13695_ _13715_/CLK line[46] vssd1 vssd1 vccd1 vccd1 _13696_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13133__D line[45] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08227__D line[106] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05213__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12646_ _12646_/A _12669_/Y vssd1 vssd1 vccd1 vccd1 _13766_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07131__D line[103] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[15\].VALID\[14\].FF_D A[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12972__D line[85] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12577_ _12595_/CLK line[47] vssd1 vssd1 vccd1 vccd1 _12578_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11528_ _11528_/A _11549_/Y vssd1 vssd1 vccd1 vccd1 _13768_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_184_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11459_ _11475_/CLK line[33] vssd1 vssd1 vccd1 vccd1 _11460_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_194_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09058__D line[88] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13158__A _13938_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13129_ _13155_/CLK line[43] vssd1 vssd1 vccd1 vccd1 _13130_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_140_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_OVHB\[25\].VALID\[13\].FF_D A[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05951_ _05951_/A _05984_/Y vssd1 vssd1 vccd1 vccd1 _13791_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_78_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13308__D line[125] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_DATA\[14\].CLKBUF\[1\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08670_ _08670_/A _08679_/Y vssd1 vssd1 vccd1 vccd1 _13710_/Z sky130_fd_sc_hd__ebufn_2
X_05882_ _05910_/CLK line[58] vssd1 vssd1 vccd1 vccd1 _05883_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07306__D line[55] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07621_ _07625_/CLK line[71] vssd1 vssd1 vccd1 vccd1 _07622_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_26_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07552_ _07552_/A _07559_/Y vssd1 vssd1 vccd1 vccd1 _13712_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_34_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[1\].VALID\[3\].FF OVHB\[1\].V/CLK A[10] vssd1 vssd1 vccd1 vccd1 OVHB\[1\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_06503_ _06505_/CLK line[72] vssd1 vssd1 vccd1 vccd1 _06504_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[18\].VALID\[14\].TOBUF OVHB\[18\].VALID\[14\].FF/Q OVHB\[18\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/B2 sky130_fd_sc_hd__ebufn_2
X_07483_ _07485_/CLK line[8] vssd1 vssd1 vccd1 vccd1 _07484_/A sky130_fd_sc_hd__dfxtp_1
XMUX.SEL0BUF\[2\] A[0] vssd1 vssd1 vccd1 vccd1 MUX.SEL0BUF\[2\]/X sky130_fd_sc_hd__clkbuf_2
XFILLER_210_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06434_ _06434_/A _06439_/Y vssd1 vssd1 vccd1 vccd1 _13714_/Z sky130_fd_sc_hd__ebufn_2
X_09222_ _09222_/A _09239_/Y vssd1 vssd1 vccd1 vccd1 _13702_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_139_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07041__D line[76] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09153_ _09165_/CLK line[3] vssd1 vssd1 vccd1 vccd1 _09154_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12882__D line[58] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06365_ _06365_/CLK line[9] vssd1 vssd1 vccd1 vccd1 _06366_/A sky130_fd_sc_hd__dfxtp_1
X_08104_ _08104_/A _08119_/Y vssd1 vssd1 vccd1 vccd1 _13704_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06880__D line[116] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05316_ _05316_/A _05319_/Y vssd1 vssd1 vccd1 vccd1 _13716_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[7\].CLKBUF\[1\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MUX.M\[3\].MUX\[4\]_A1 _13727_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09084_ _09084_/A _09099_/Y vssd1 vssd1 vccd1 vccd1 _13844_/Z sky130_fd_sc_hd__ebufn_2
X_06296_ _06296_/A _06299_/Y vssd1 vssd1 vccd1 vccd1 _13856_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11498__D line[51] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08035_ _08045_/CLK line[4] vssd1 vssd1 vccd1 vccd1 _08036_/A sky130_fd_sc_hd__dfxtp_1
X_05247_ _05247_/CLK _05248_/X vssd1 vssd1 vccd1 vccd1 _05245_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_162_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05178_ _13931_/Y wr vssd1 vssd1 vccd1 vccd1 _05178_/X sky130_fd_sc_hd__and2_1
X_09986_ _09986_/A _10009_/Y vssd1 vssd1 vccd1 vccd1 _13626_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_67_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08937_ _08955_/CLK line[47] vssd1 vssd1 vccd1 vccd1 _08938_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_29_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XOVHB\[11\].VALID\[13\].TOBUF OVHB\[11\].VALID\[13\].FF/Q OVHB\[11\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04916_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_85_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12122__D line[95] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[17\].VALID\[10\].FF_D A[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08868_ _08868_/A _08889_/Y vssd1 vssd1 vccd1 vccd1 _13628_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07216__D line[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06120__D line[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07819_ _07835_/CLK line[33] vssd1 vssd1 vccd1 vccd1 _07820_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11961__D line[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_MUX.M\[1\].MUX\[0\]_A2 _13784_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08799_ _08815_/CLK line[97] vssd1 vssd1 vccd1 vccd1 _08800_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[9\].CGAND _13899_/X wr vssd1 vssd1 vccd1 vccd1 OVHB\[9\].CGAND/X sky130_fd_sc_hd__and2_4
X_10830_ _10830_/A _10849_/Y vssd1 vssd1 vccd1 vccd1 _13630_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09431__D line[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10761_ _10775_/CLK line[98] vssd1 vssd1 vccd1 vccd1 _10762_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_13_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12500_ _12500_/A _12529_/Y vssd1 vssd1 vccd1 vccd1 _13620_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_12_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10692_ _10692_/A _10709_/Y vssd1 vssd1 vccd1 vccd1 _13772_/Z sky130_fd_sc_hd__ebufn_2
X_13480_ _13480_/A _13509_/Y vssd1 vssd1 vccd1 vccd1 _13760_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_197_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13888__D line[120] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12431_ _12455_/CLK line[108] vssd1 vssd1 vccd1 vccd1 _12432_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_185_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XOVHB\[7\].VALID\[6\].TOBUF OVHB\[7\].VALID\[6\].FF/Q OVHB\[7\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04923_/A2 sky130_fd_sc_hd__ebufn_2
XANTENNA__06790__D line[80] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12362_ _12362_/A _12389_/Y vssd1 vssd1 vccd1 vccd1 _13762_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[30\].INV _13970_/X vssd1 vssd1 vccd1 vccd1 OVHB\[30\].INV/Y sky130_fd_sc_hd__inv_2
XFILLER_138_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11313_ _11335_/CLK line[109] vssd1 vssd1 vccd1 vccd1 _11314_/A sky130_fd_sc_hd__dfxtp_1
X_12293_ _12315_/CLK line[45] vssd1 vssd1 vccd1 vccd1 _12294_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_153_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11244_ _11244_/A _11269_/Y vssd1 vssd1 vccd1 vccd1 _13764_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05984__A _13902_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11175_ _11195_/CLK line[46] vssd1 vssd1 vccd1 vccd1 _11176_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09606__D line[82] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10126_ _10126_/A _10149_/Y vssd1 vssd1 vccd1 vccd1 _13766_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_48_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10057_ _10075_/CLK line[47] vssd1 vssd1 vccd1 vccd1 _10058_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09903__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06030__D line[126] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11871__D line[108] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06965__D line[32] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13816_ _13820_/CLK line[87] vssd1 vssd1 vccd1 vccd1 _13817_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[2\].CLKBUF\[5\] clk vssd1 vssd1 vccd1 vccd1 _11302_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_44_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10487__D line[101] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13747_ _13747_/A _13754_/Y vssd1 vssd1 vccd1 vccd1 _13747_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_43_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10959_ _10985_/CLK line[75] vssd1 vssd1 vccd1 vccd1 _10960_/A sky130_fd_sc_hd__dfxtp_1
X_13678_ _13680_/CLK line[24] vssd1 vssd1 vccd1 vccd1 _13679_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_31_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13798__D line[93] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05878__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12629_ _12629_/A _12634_/Y vssd1 vssd1 vccd1 vccd1 _13749_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07796__D line[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06150_ _06150_/A _06159_/Y vssd1 vssd1 vccd1 vccd1 _13710_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_156_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05101_ _05105_/CLK line[71] vssd1 vssd1 vccd1 vccd1 _05102_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_208_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06081_ _06085_/CLK line[7] vssd1 vssd1 vccd1 vccd1 _06082_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[31\].VALID\[13\].TOBUF OVHB\[31\].VALID\[13\].FF/Q OVHB\[31\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04916_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__11111__D line[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05032_ _05032_/A _05039_/Y vssd1 vssd1 vccd1 vccd1 _13712_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06205__D line[78] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[20\].VALID\[5\].FF_D A[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10950__D line[57] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09840_ _09840_/A _09869_/Y vssd1 vssd1 vccd1 vccd1 _13760_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08420__D line[52] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09771_ _09795_/CLK line[44] vssd1 vssd1 vccd1 vccd1 _09772_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[14\].VALID\[1\].TOBUF OVHB\[14\].VALID\[1\].FF/Q OVHB\[14\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04926_/B2 sky130_fd_sc_hd__ebufn_2
X_06983_ _06995_/CLK line[35] vssd1 vssd1 vccd1 vccd1 _06984_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_85_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13038__D line[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08722_ _08722_/A _08749_/Y vssd1 vssd1 vccd1 vccd1 _13762_/Z sky130_fd_sc_hd__ebufn_2
X_05934_ _05934_/A _05949_/Y vssd1 vssd1 vccd1 vccd1 _13774_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[13\].VALID\[9\].FF_D A[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XOVHB\[24\].VALID\[13\].FF OVHB\[24\].V/CLK A[20] vssd1 vssd1 vccd1 vccd1 OVHB\[24\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_05865_ _05875_/CLK line[36] vssd1 vssd1 vccd1 vccd1 _05866_/A sky130_fd_sc_hd__dfxtp_1
X_08653_ _08675_/CLK line[45] vssd1 vssd1 vccd1 vccd1 _08654_/A sky130_fd_sc_hd__dfxtp_1
X_07604_ _07604_/A _07629_/Y vssd1 vssd1 vccd1 vccd1 _13764_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08584_ _08584_/A _08609_/Y vssd1 vssd1 vccd1 vccd1 _13624_/Z sky130_fd_sc_hd__ebufn_2
X_05796_ _05796_/A _05809_/Y vssd1 vssd1 vccd1 vccd1 _13636_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10397__D line[74] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07535_ _07555_/CLK line[46] vssd1 vssd1 vccd1 vccd1 _07536_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[12\].CLKBUF\[3\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07466_ _07466_/A _07489_/Y vssd1 vssd1 vccd1 vccd1 _13626_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[26\].VALID\[0\].FF OVHB\[26\].V/CLK A[7] vssd1 vssd1 vccd1 vccd1 OVHB\[26\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_167_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06417_ _06435_/CLK line[47] vssd1 vssd1 vccd1 vccd1 _06418_/A sky130_fd_sc_hd__dfxtp_1
X_09205_ _09235_/CLK line[32] vssd1 vssd1 vccd1 vccd1 _09206_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[1\].CLKBUF\[2\] clk vssd1 vssd1 vccd1 vccd1 _08117_/CLK sky130_fd_sc_hd__clkbuf_4
X_07397_ _07415_/CLK line[111] vssd1 vssd1 vccd1 vccd1 _07398_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13501__D line[71] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09136_ _09136_/A _09169_/Y vssd1 vssd1 vccd1 vccd1 _13616_/Z sky130_fd_sc_hd__ebufn_2
X_06348_ _06348_/A _06369_/Y vssd1 vssd1 vccd1 vccd1 _13628_/Z sky130_fd_sc_hd__ebufn_2
X_09067_ _09095_/CLK line[106] vssd1 vssd1 vccd1 vccd1 _09068_/A sky130_fd_sc_hd__dfxtp_1
X_06279_ _06295_/CLK line[97] vssd1 vssd1 vccd1 vccd1 _06280_/A sky130_fd_sc_hd__dfxtp_1
X_08018_ _08018_/A _08049_/Y vssd1 vssd1 vccd1 vccd1 _13618_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_78_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10860__D line[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_DATA\[5\].CLKBUF\[3\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05954__D line[91] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08330__D line[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09969_ _09969_/A _09974_/Y vssd1 vssd1 vccd1 vccd1 _13889_/Z sky130_fd_sc_hd__ebufn_2
X_12980_ _12980_/CLK line[89] vssd1 vssd1 vccd1 vccd1 _12981_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_92_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_DATA\[31\].CLKBUF\[5\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDATA\[31\].CLKBUF\[0\] clk vssd1 vssd1 vccd1 vccd1 _11687_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__07524__A _13911_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11931_ _11931_/A _11934_/Y vssd1 vssd1 vccd1 vccd1 _13891_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12787__D line[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_OVHB\[1\].VALID\[0\].FF_D A[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07243__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06785__D line[73] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11862_ _11862_/CLK _11863_/X vssd1 vssd1 vccd1 vccd1 _11860_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__09161__D line[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XDATA\[21\].CLKBUF\[6\] clk vssd1 vssd1 vccd1 vccd1 _08817_/CLK sky130_fd_sc_hd__clkbuf_4
X_13601_ _13601_/A _13614_/Y vssd1 vssd1 vccd1 vccd1 _13881_/Z sky130_fd_sc_hd__ebufn_2
X_10813_ _13924_/X wr vssd1 vssd1 vccd1 vccd1 _10813_/X sky130_fd_sc_hd__and2_1
XFILLER_198_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11793_ _13927_/X wr vssd1 vssd1 vccd1 vccd1 _11793_/X sky130_fd_sc_hd__and2_1
XFILLER_13_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XOVHB\[20\].VALID\[0\].TOBUF OVHB\[20\].VALID\[0\].FF/Q OVHB\[20\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04924_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_13_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10100__D line[52] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MUX.M\[0\].MUX\[1\]_A0 _13630_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13532_ _13540_/CLK line[85] vssd1 vssd1 vccd1 vccd1 _13533_/A sky130_fd_sc_hd__dfxtp_1
X_10744_ _13924_/X vssd1 vssd1 vccd1 vccd1 _10744_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13463_ _13463_/A _13474_/Y vssd1 vssd1 vccd1 vccd1 _13743_/Z sky130_fd_sc_hd__ebufn_2
X_10675_ _10705_/CLK line[64] vssd1 vssd1 vccd1 vccd1 _10676_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13411__D line[44] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12414_ _12420_/CLK line[86] vssd1 vssd1 vccd1 vccd1 _12415_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08505__D line[96] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13394_ _13400_/CLK line[22] vssd1 vssd1 vccd1 vccd1 _13395_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_154_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12345_ _12345_/A _12354_/Y vssd1 vssd1 vccd1 vccd1 _13745_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12027__D line[37] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[24\].VALID\[2\].FF OVHB\[24\].V/CLK A[9] vssd1 vssd1 vccd1 vccd1 OVHB\[24\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_154_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12276_ _12280_/CLK line[23] vssd1 vssd1 vccd1 vccd1 _12277_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_99_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11227_ _11227_/A _11234_/Y vssd1 vssd1 vccd1 vccd1 _13747_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_141_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07418__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09336__D line[87] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_OVHB\[26\].VALID\[9\].FF_D A[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11158_ _11160_/CLK line[24] vssd1 vssd1 vccd1 vccd1 _11159_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_67_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10109_ _10109_/A _10114_/Y vssd1 vssd1 vccd1 vccd1 _13749_/Z sky130_fd_sc_hd__ebufn_2
X_11089_ _11089_/A _11094_/Y vssd1 vssd1 vccd1 vccd1 _13889_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_83_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05650_ _05650_/A _05669_/Y vssd1 vssd1 vccd1 vccd1 _13770_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06695__D line[46] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09071__D line[108] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05581_ _05595_/CLK line[34] vssd1 vssd1 vccd1 vccd1 _05582_/A sky130_fd_sc_hd__dfxtp_1
X_07320_ _07320_/A _07349_/Y vssd1 vssd1 vccd1 vccd1 _13760_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10010__D line[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XDATA\[20\].CLKBUF\[3\] clk vssd1 vssd1 vccd1 vccd1 _08432_/CLK sky130_fd_sc_hd__clkbuf_4
X_07251_ _07275_/CLK line[44] vssd1 vssd1 vccd1 vccd1 _07252_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_31_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[12\].VALID\[6\].TOBUF OVHB\[12\].VALID\[6\].FF/Q OVHB\[12\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04923_/A2 sky130_fd_sc_hd__ebufn_2
X_06202_ _06202_/A _06229_/Y vssd1 vssd1 vccd1 vccd1 _13762_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__04943__D line[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07182_ _07182_/A _07209_/Y vssd1 vssd1 vccd1 vccd1 _13622_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_145_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06133_ _06155_/CLK line[45] vssd1 vssd1 vccd1 vccd1 _06134_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_144_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XOVHB\[5\].VALID\[10\].TOBUF OVHB\[5\].VALID\[10\].FF/Q OVHB\[5\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04932_/B2 sky130_fd_sc_hd__ebufn_2
X_06064_ _06064_/A _06089_/Y vssd1 vssd1 vccd1 vccd1 _13624_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_172_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11776__D line[50] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05015_ _05035_/CLK line[46] vssd1 vssd1 vccd1 vccd1 _05016_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_160_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09246__D line[60] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08150__D line[57] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09823_ _09823_/A _09834_/Y vssd1 vssd1 vccd1 vccd1 _13743_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_100_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09754_ _09760_/CLK line[22] vssd1 vssd1 vccd1 vccd1 _09755_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__04968__A _13931_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06966_ _06966_/A _06999_/Y vssd1 vssd1 vccd1 vccd1 _13686_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[22\].VALID\[4\].FF OVHB\[22\].V/CLK A[11] vssd1 vssd1 vccd1 vccd1 OVHB\[22\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_08705_ _08705_/A _08714_/Y vssd1 vssd1 vccd1 vccd1 _13745_/Z sky130_fd_sc_hd__ebufn_2
X_05917_ _05945_/CLK line[74] vssd1 vssd1 vccd1 vccd1 _05918_/A sky130_fd_sc_hd__dfxtp_1
X_09685_ _09685_/A _09694_/Y vssd1 vssd1 vccd1 vccd1 _13885_/Z sky130_fd_sc_hd__ebufn_2
X_06897_ _06925_/CLK line[10] vssd1 vssd1 vccd1 vccd1 _06898_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12400__D line[94] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08636_ _08640_/CLK line[23] vssd1 vssd1 vccd1 vccd1 _08637_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_54_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05848_ _05848_/A _05879_/Y vssd1 vssd1 vccd1 vccd1 _13688_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[0\].INV _13975_/Y vssd1 vssd1 vccd1 vccd1 OVHB\[0\].INV/Y sky130_fd_sc_hd__inv_2
XPHY_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08567_ _08567_/A _08574_/Y vssd1 vssd1 vccd1 vccd1 _13887_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05779_ _05805_/CLK line[11] vssd1 vssd1 vccd1 vccd1 _05780_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11016__D line[87] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[7\].VALID\[4\].FF_D A[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07518_ _07520_/CLK line[24] vssd1 vssd1 vccd1 vccd1 _07519_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08498_ _08500_/CLK line[88] vssd1 vssd1 vccd1 vccd1 _08499_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07449_ _07449_/A _07454_/Y vssd1 vssd1 vccd1 vccd1 _13889_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[6\].CG_CLK clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08325__D line[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10460_ _10460_/CLK line[89] vssd1 vssd1 vccd1 vccd1 _10461_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[10\].CLKBUF\[5\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09119_ _09119_/A _09134_/Y vssd1 vssd1 vccd1 vccd1 _13879_/Z sky130_fd_sc_hd__ebufn_2
X_10391_ _10391_/A _10394_/Y vssd1 vssd1 vccd1 vccd1 _13751_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_89_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12130_ _12140_/CLK line[84] vssd1 vssd1 vccd1 vccd1 _12131_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10590__D line[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12061_ _12061_/A _12074_/Y vssd1 vssd1 vccd1 vccd1 _13741_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[20\].VALID\[11\].FF OVHB\[20\].V/CLK A[18] vssd1 vssd1 vccd1 vccd1 OVHB\[20\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__05684__D line[81] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08060__D line[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05039__A _13931_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11012_ _11020_/CLK line[85] vssd1 vssd1 vccd1 vccd1 _11013_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_49_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08995__D line[64] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12963_ _12963_/A _12984_/Y vssd1 vssd1 vccd1 vccd1 _13803_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_92_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_DATA\[3\].CLKBUF\[5\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11914_ _11930_/CLK line[113] vssd1 vssd1 vccd1 vccd1 _11915_/A sky130_fd_sc_hd__dfxtp_1
X_12894_ _12910_/CLK line[49] vssd1 vssd1 vccd1 vccd1 _12895_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_72_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11845_ _11845_/A _11864_/Y vssd1 vssd1 vccd1 vccd1 _13805_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[20\].VALID\[6\].FF OVHB\[20\].V/CLK A[13] vssd1 vssd1 vccd1 vccd1 OVHB\[20\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_159_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11776_ _11790_/CLK line[50] vssd1 vssd1 vccd1 vccd1 _11777_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_201_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10765__D line[100] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13515_ _13515_/A _13544_/Y vssd1 vssd1 vccd1 vccd1 _13795_/Z sky130_fd_sc_hd__ebufn_2
X_10727_ _10727_/A _10744_/Y vssd1 vssd1 vccd1 vccd1 _13807_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_41_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05859__D line[33] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13141__D line[34] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[10\].VALID\[13\].FF OVHB\[10\].V/CLK A[20] vssd1 vssd1 vccd1 vccd1 OVHB\[10\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_201_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13446_ _13470_/CLK line[60] vssd1 vssd1 vccd1 vccd1 _13447_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08235__D line[110] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10658_ _10670_/CLK line[51] vssd1 vssd1 vccd1 vccd1 _10659_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_70_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12980__D line[89] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13377_ _13377_/A _13404_/Y vssd1 vssd1 vccd1 vccd1 _13657_/Z sky130_fd_sc_hd__ebufn_2
X_10589_ _10589_/A _10604_/Y vssd1 vssd1 vccd1 vccd1 _13669_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_142_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12328_ _12350_/CLK line[61] vssd1 vssd1 vccd1 vccd1 _12329_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_115_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06333__A _13903_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12259_ _12259_/A _12284_/Y vssd1 vssd1 vccd1 vccd1 _13659_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[28\].VALID\[12\].TOBUF OVHB\[28\].VALID\[12\].FF/Q OVHB\[28\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04929_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_96_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10005__D line[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06820_ _06820_/CLK line[89] vssd1 vssd1 vccd1 vccd1 _06821_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_95_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06751_ _06751_/A _06754_/Y vssd1 vssd1 vccd1 vccd1 _13751_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13316__D line[114] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05702_ _05702_/CLK _05703_/X vssd1 vssd1 vccd1 vccd1 _05700_/CLK sky130_fd_sc_hd__dlclkp_1
X_09470_ _09480_/CLK line[20] vssd1 vssd1 vccd1 vccd1 _09471_/A sky130_fd_sc_hd__dfxtp_1
X_06682_ _06682_/CLK _06683_/X vssd1 vssd1 vccd1 vccd1 _06680_/CLK sky130_fd_sc_hd__dlclkp_1
X_08421_ _08421_/A _08434_/Y vssd1 vssd1 vccd1 vccd1 _13741_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[19\].VALID\[7\].FF OVHB\[19\].V/CLK A[14] vssd1 vssd1 vccd1 vccd1 OVHB\[19\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13613__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05633_ _13901_/X wr vssd1 vssd1 vccd1 vccd1 _05633_/X sky130_fd_sc_hd__and2_1
X_08352_ _08360_/CLK line[21] vssd1 vssd1 vccd1 vccd1 _08353_/A sky130_fd_sc_hd__dfxtp_1
X_05564_ _13901_/X vssd1 vssd1 vccd1 vccd1 _05564_/Y sky130_fd_sc_hd__inv_2
XANTENNA__06508__A _13904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07303_ _07303_/A _07314_/Y vssd1 vssd1 vccd1 vccd1 _13743_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_32_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10675__D line[64] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05495_ _05525_/CLK line[0] vssd1 vssd1 vccd1 vccd1 _05496_/A sky130_fd_sc_hd__dfxtp_1
X_08283_ _08283_/A _08294_/Y vssd1 vssd1 vccd1 vccd1 _13883_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[27\].VALID\[0\].TOBUF OVHB\[27\].VALID\[0\].FF/Q OVHB\[27\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04924_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_177_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07234_ _07240_/CLK line[22] vssd1 vssd1 vccd1 vccd1 _07235_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_158_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XOVHB\[21\].VALID\[11\].TOBUF OVHB\[21\].VALID\[11\].FF/Q OVHB\[21\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04915_/B2 sky130_fd_sc_hd__ebufn_2
X_07165_ _07165_/A _07174_/Y vssd1 vssd1 vccd1 vccd1 _13885_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12890__D line[62] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07984__D line[123] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06116_ _06120_/CLK line[23] vssd1 vssd1 vccd1 vccd1 _06117_/A sky130_fd_sc_hd__dfxtp_1
X_07096_ _07100_/CLK line[87] vssd1 vssd1 vccd1 vccd1 _07097_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[1\].CGAND_A _13932_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06047_ _06047_/A _06054_/Y vssd1 vssd1 vccd1 vccd1 _13887_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09554__A _13920_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MUX.M\[2\].MUX\[2\]_A2 _13807_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09806_ _09830_/CLK line[60] vssd1 vssd1 vccd1 vccd1 _09807_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09273__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05009__D line[43] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07998_ _08010_/CLK line[115] vssd1 vssd1 vccd1 vccd1 _07999_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_87_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09737_ _09737_/A _09764_/Y vssd1 vssd1 vccd1 vccd1 _13657_/Z sky130_fd_sc_hd__ebufn_2
X_06949_ _06949_/A _06964_/Y vssd1 vssd1 vccd1 vccd1 _13669_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12130__D line[84] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09668_ _09690_/CLK line[125] vssd1 vssd1 vccd1 vccd1 _09669_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07224__D line[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08619_ _08619_/A _08644_/Y vssd1 vssd1 vccd1 vccd1 _13659_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09599_ _09599_/A _09624_/Y vssd1 vssd1 vccd1 vccd1 _13799_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11630_ _11650_/CLK line[126] vssd1 vssd1 vccd1 vccd1 _11631_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11561_ _11561_/A _11584_/Y vssd1 vssd1 vccd1 vccd1 _13801_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13300_ _13330_/CLK line[112] vssd1 vssd1 vccd1 vccd1 _13301_/A sky130_fd_sc_hd__dfxtp_1
X_10512_ _10530_/CLK line[127] vssd1 vssd1 vccd1 vccd1 _10513_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09729__A _13921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11492_ _11510_/CLK line[63] vssd1 vssd1 vccd1 vccd1 _11493_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[17\].VALID\[9\].FF OVHB\[17\].V/CLK A[16] vssd1 vssd1 vccd1 vccd1 OVHB\[17\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13231_ _13231_/A _13264_/Y vssd1 vssd1 vccd1 vccd1 _13791_/Z sky130_fd_sc_hd__ebufn_2
X_10443_ _10443_/A _10464_/Y vssd1 vssd1 vccd1 vccd1 _13803_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09448__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XOVHB\[19\].VALID\[6\].TOBUF OVHB\[19\].VALID\[6\].FF/Q OVHB\[19\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04923_/A2 sky130_fd_sc_hd__ebufn_2
XFILLER_156_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13162_ _13190_/CLK line[58] vssd1 vssd1 vccd1 vccd1 _13163_/A sky130_fd_sc_hd__dfxtp_1
X_10374_ _10390_/CLK line[49] vssd1 vssd1 vccd1 vccd1 _10375_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_163_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12113_ _12113_/A _12144_/Y vssd1 vssd1 vccd1 vccd1 _13793_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12305__D line[36] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13093_ _13093_/A _13124_/Y vssd1 vssd1 vccd1 vccd1 _13653_/Z sky130_fd_sc_hd__ebufn_2
X_12044_ _12070_/CLK line[59] vssd1 vssd1 vccd1 vccd1 _12045_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_77_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09614__D line[86] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_OVHB\[2\].VALID\[13\].FF_D A[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12040__D line[48] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12946_ _12946_/A _12949_/Y vssd1 vssd1 vccd1 vccd1 _13786_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_206_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12877_ _12877_/CLK _12878_/X vssd1 vssd1 vccd1 vccd1 _12875_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__11234__A _13933_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06973__D line[45] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11828_ _13927_/X wr vssd1 vssd1 vccd1 vccd1 _11828_/X sky130_fd_sc_hd__and2_1
XFILLER_187_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[12\].VALID\[0\].FF_D A[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10495__D line[105] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11759_ _13927_/X vssd1 vssd1 vccd1 vccd1 _11759_/Y sky130_fd_sc_hd__inv_2
XANTENNA_DATA\[1\].CLKBUF\[7\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05589__D line[38] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05280_ _05280_/CLK line[25] vssd1 vssd1 vccd1 vccd1 _05281_/A sky130_fd_sc_hd__dfxtp_1
X_13429_ _13435_/CLK line[38] vssd1 vssd1 vccd1 vccd1 _13430_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12215__D line[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08970_ _08990_/CLK line[62] vssd1 vssd1 vccd1 vccd1 _08971_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06998__A _13909_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[29\].VALID\[13\].FF OVHB\[29\].V/CLK A[20] vssd1 vssd1 vccd1 vccd1 OVHB\[29\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06213__D line[67] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07921_ _07921_/A _07944_/Y vssd1 vssd1 vccd1 vccd1 _13801_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[0\].VALID\[2\].TOBUF OVHB\[0\].VALID\[2\].FF/Q OVHB\[0\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04930_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_96_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11409__A _13926_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07852_ _07870_/CLK line[63] vssd1 vssd1 vccd1 vccd1 _07853_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_84_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09524__D line[59] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[25\].VALID\[5\].TOBUF OVHB\[25\].VALID\[5\].FF/Q OVHB\[25\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04927_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_84_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06803_ _06803_/A _06824_/Y vssd1 vssd1 vccd1 vccd1 _13803_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11128__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07783_ _07783_/A _07804_/Y vssd1 vssd1 vccd1 vccd1 _13663_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_84_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_04995_ _04995_/A _05004_/Y vssd1 vssd1 vccd1 vccd1 _13675_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13046__D line[119] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09522_ _09550_/CLK line[58] vssd1 vssd1 vccd1 vccd1 _09523_/A sky130_fd_sc_hd__dfxtp_1
X_06734_ _06750_/CLK line[49] vssd1 vssd1 vccd1 vccd1 _06735_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[31\].CG clk OVHB\[31\].CGAND/X vssd1 vssd1 vccd1 vccd1 OVHB\[31\].V/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA_OVHB\[3\].VALID\[7\].FF_D A[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09453_ _09453_/A _09484_/Y vssd1 vssd1 vccd1 vccd1 _13653_/Z sky130_fd_sc_hd__ebufn_2
X_06665_ _06665_/A _06684_/Y vssd1 vssd1 vccd1 vccd1 _13665_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_36_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08404_ _08430_/CLK line[59] vssd1 vssd1 vccd1 vccd1 _08405_/A sky130_fd_sc_hd__dfxtp_1
XPHY_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05616_ _05630_/CLK line[50] vssd1 vssd1 vccd1 vccd1 _05617_/A sky130_fd_sc_hd__dfxtp_1
X_09384_ _09410_/CLK line[123] vssd1 vssd1 vccd1 vccd1 _09385_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_101_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06596_ _06610_/CLK line[114] vssd1 vssd1 vccd1 vccd1 _06597_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_178_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08335_ _08335_/A _08364_/Y vssd1 vssd1 vccd1 vccd1 _13655_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_51_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XOVHB\[3\].CG clk OVHB\[3\].CGAND/X vssd1 vssd1 vccd1 vccd1 OVHB\[3\].V/CLK sky130_fd_sc_hd__dlclkp_1
X_05547_ _05547_/A _05564_/Y vssd1 vssd1 vccd1 vccd1 _13667_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05499__D line[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05478_ _05490_/CLK line[115] vssd1 vssd1 vccd1 vccd1 _05479_/A sky130_fd_sc_hd__dfxtp_1
X_08266_ _08290_/CLK line[124] vssd1 vssd1 vccd1 vccd1 _08267_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_20_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[1\].V_RESET_B rst_n vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07217_ _07217_/A _07244_/Y vssd1 vssd1 vccd1 vccd1 _13657_/Z sky130_fd_sc_hd__ebufn_2
X_08197_ _08197_/A _08224_/Y vssd1 vssd1 vccd1 vccd1 _13797_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07069__A _13909_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07148_ _07170_/CLK line[125] vssd1 vssd1 vccd1 vccd1 _07149_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08603__D line[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07079_ _07079_/A _07104_/Y vssd1 vssd1 vccd1 vccd1 _13799_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_10_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12703__A _13936_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10090_ _10110_/CLK line[62] vssd1 vssd1 vccd1 vccd1 _10091_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_102_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05962__D line[95] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MUX.M\[1\].MUX\[3\]_A0 _13620_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12800_ _12800_/A _12809_/Y vssd1 vssd1 vccd1 vccd1 _13640_/Z sky130_fd_sc_hd__ebufn_2
X_13780_ _13780_/A _13789_/Y vssd1 vssd1 vccd1 vccd1 _13780_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_142_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10992_ _11020_/CLK line[90] vssd1 vssd1 vccd1 vccd1 _10993_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_16_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12731_ _12735_/CLK line[103] vssd1 vssd1 vccd1 vccd1 _12732_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12795__D line[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[25\].VALID\[0\].FF_D A[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07889__D line[65] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12662_ _12662_/A _12669_/Y vssd1 vssd1 vccd1 vccd1 _13782_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11613_ _11615_/CLK line[104] vssd1 vssd1 vccd1 vccd1 _11614_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_42_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[31\].VALID\[4\].TOBUF OVHB\[31\].VALID\[4\].FF/Q OVHB\[31\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04925_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_168_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12593_ _12595_/CLK line[40] vssd1 vssd1 vccd1 vccd1 _12594_/A sky130_fd_sc_hd__dfxtp_1
XPHY_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11204__D line[59] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11544_ _11544_/A _11549_/Y vssd1 vssd1 vccd1 vccd1 _13784_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08363__A _13913_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05202__D line[117] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[18\].VALID\[4\].FF_D A[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11475_ _11475_/CLK line[41] vssd1 vssd1 vccd1 vccd1 _11476_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_137_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13214_ _13214_/A _13229_/Y vssd1 vssd1 vccd1 vccd1 _13774_/Z sky130_fd_sc_hd__ebufn_2
X_10426_ _10426_/A _10429_/Y vssd1 vssd1 vccd1 vccd1 _13786_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08513__D line[109] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[22\].CLKBUF\[1\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12035__D line[41] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13145_ _13155_/CLK line[36] vssd1 vssd1 vccd1 vccd1 _13146_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_98_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10357_ _10357_/CLK _10358_/X vssd1 vssd1 vccd1 vccd1 _10355_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__07129__D line[102] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13076_ _13076_/A _13089_/Y vssd1 vssd1 vccd1 vccd1 _13636_/Z sky130_fd_sc_hd__ebufn_2
X_10288_ _13923_/X wr vssd1 vssd1 vccd1 vccd1 _10288_/X sky130_fd_sc_hd__and2_1
X_12027_ _12035_/CLK line[37] vssd1 vssd1 vccd1 vccd1 _12028_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_38_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13978_ _13982_/C _13982_/B _13982_/A _13982_/D vssd1 vssd1 vccd1 vccd1 _13978_/X
+ sky130_fd_sc_hd__and4b_4
XFILLER_19_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08538__A _13913_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12929_ _12945_/CLK line[65] vssd1 vssd1 vccd1 vccd1 _12930_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_34_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06450_ _06470_/CLK line[62] vssd1 vssd1 vccd1 vccd1 _06451_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_22_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XOVHB\[1\].VALID\[13\].FF OVHB\[1\].V/CLK A[20] vssd1 vssd1 vccd1 vccd1 OVHB\[1\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_05401_ _05401_/A _05424_/Y vssd1 vssd1 vccd1 vccd1 _13801_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11899__A _13927_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06381_ _06381_/A _06404_/Y vssd1 vssd1 vccd1 vccd1 _13661_/Z sky130_fd_sc_hd__ebufn_2
X_05332_ _05350_/CLK line[63] vssd1 vssd1 vccd1 vccd1 _05333_/A sky130_fd_sc_hd__dfxtp_1
X_08120_ _08150_/CLK line[48] vssd1 vssd1 vccd1 vccd1 _08121_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05112__D line[90] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08051_ _08051_/A _08084_/Y vssd1 vssd1 vccd1 vccd1 _13651_/Z sky130_fd_sc_hd__ebufn_2
X_05263_ _05263_/A _05284_/Y vssd1 vssd1 vccd1 vccd1 _13663_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_119_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07002_ _07030_/CLK line[58] vssd1 vssd1 vccd1 vccd1 _07003_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__04951__D line[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05194_ _05210_/CLK line[113] vssd1 vssd1 vccd1 vccd1 _05195_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_127_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[18\].VALID\[10\].TOBUF OVHB\[18\].VALID\[10\].FF/Q OVHB\[18\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04932_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__07039__D line[75] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08953_ _08955_/CLK line[40] vssd1 vssd1 vccd1 vccd1 _08954_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11784__D line[54] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07904_ _07904_/A _07909_/Y vssd1 vssd1 vccd1 vccd1 _13784_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[8\].VALID\[4\].FF OVHB\[8\].V/CLK A[11] vssd1 vssd1 vccd1 vccd1 OVHB\[8\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06878__D line[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10043__A _13922_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08884_ _08884_/A _08889_/Y vssd1 vssd1 vccd1 vccd1 _13644_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09254__D line[49] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07835_ _07835_/CLK line[41] vssd1 vssd1 vccd1 vccd1 _07836_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_56_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07766_ _07766_/A _07769_/Y vssd1 vssd1 vccd1 vccd1 _13646_/Z sky130_fd_sc_hd__ebufn_2
X_04978_ _05000_/CLK line[29] vssd1 vssd1 vccd1 vccd1 _04979_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_37_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09505_ _09515_/CLK line[36] vssd1 vssd1 vccd1 vccd1 _09506_/A sky130_fd_sc_hd__dfxtp_1
X_06717_ _06717_/CLK _06718_/X vssd1 vssd1 vccd1 vccd1 _06715_/CLK sky130_fd_sc_hd__dlclkp_1
X_07697_ _07697_/CLK _07698_/X vssd1 vssd1 vccd1 vccd1 _07695_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_197_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_OVHB\[9\].VALID\[13\].FF_D A[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09436_ _09436_/A _09449_/Y vssd1 vssd1 vccd1 vccd1 _13636_/Z sky130_fd_sc_hd__ebufn_2
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06648_ _13905_/X wr vssd1 vssd1 vccd1 vccd1 _06648_/X sky130_fd_sc_hd__and2_1
XFILLER_169_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07502__D line[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09367_ _09375_/CLK line[101] vssd1 vssd1 vccd1 vccd1 _09368_/A sky130_fd_sc_hd__dfxtp_1
X_06579_ _13904_/X vssd1 vssd1 vccd1 vccd1 _06579_/Y sky130_fd_sc_hd__inv_2
XFILLER_184_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08318_ _08318_/A _08329_/Y vssd1 vssd1 vccd1 vccd1 _13638_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06118__D line[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09298_ _09298_/A _09309_/Y vssd1 vssd1 vccd1 vccd1 _13778_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[25\].VALID\[11\].FF OVHB\[25\].V/CLK A[18] vssd1 vssd1 vccd1 vccd1 OVHB\[25\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11959__D line[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08249_ _08255_/CLK line[102] vssd1 vssd1 vccd1 vccd1 _08250_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10218__A _13922_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09429__D line[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11260_ _11260_/A _11269_/Y vssd1 vssd1 vccd1 vccd1 _13780_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[5\].CGAND _13936_/X wr vssd1 vssd1 vccd1 vccd1 OVHB\[5\].CGAND/X sky130_fd_sc_hd__and2_4
XFILLER_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10211_ _10215_/CLK line[103] vssd1 vssd1 vccd1 vccd1 _10212_/A sky130_fd_sc_hd__dfxtp_1
X_11191_ _11195_/CLK line[39] vssd1 vssd1 vccd1 vccd1 _11192_/A sky130_fd_sc_hd__dfxtp_1
X_10142_ _10142_/A _10149_/Y vssd1 vssd1 vccd1 vccd1 _13782_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_133_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11694__D line[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10073_ _10075_/CLK line[40] vssd1 vssd1 vccd1 vccd1 _10074_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_121_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05692__D line[85] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13901_ _13905_/C _13905_/B _13905_/A _13905_/D vssd1 vssd1 vccd1 vccd1 _13901_/X
+ sky130_fd_sc_hd__and4b_4
XOVHB\[7\].VALID\[2\].TOBUF OVHB\[7\].VALID\[2\].FF/Q OVHB\[7\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04930_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__13264__A _13938_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13832_ _13832_/A _13859_/Y vssd1 vssd1 vccd1 vccd1 _13832_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_35_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13763_ _13785_/CLK line[77] vssd1 vssd1 vccd1 vccd1 _13764_/A sky130_fd_sc_hd__dfxtp_1
X_10975_ _10985_/CLK line[68] vssd1 vssd1 vccd1 vccd1 _10976_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[15\].VALID\[13\].FF OVHB\[15\].V/CLK A[20] vssd1 vssd1 vccd1 vccd1 OVHB\[15\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XOVHB\[6\].VALID\[6\].FF OVHB\[6\].V/CLK A[13] vssd1 vssd1 vccd1 vccd1 OVHB\[6\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12714_ _12714_/A _12739_/Y vssd1 vssd1 vccd1 vccd1 _13834_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_16_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13694_ _13694_/A _13719_/Y vssd1 vssd1 vccd1 vccd1 _13694_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_71_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12645_ _12665_/CLK line[78] vssd1 vssd1 vccd1 vccd1 _12646_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_30_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06028__D line[125] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12576_ _12576_/A _12599_/Y vssd1 vssd1 vccd1 vccd1 _13696_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11869__D line[107] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10773__D line[104] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11527_ _11545_/CLK line[79] vssd1 vssd1 vccd1 vccd1 _11528_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_172_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05867__D line[37] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08243__D line[99] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11458_ _11458_/A _11479_/Y vssd1 vssd1 vccd1 vccd1 _13698_/Z sky130_fd_sc_hd__ebufn_2
X_10409_ _10425_/CLK line[65] vssd1 vssd1 vccd1 vccd1 _10410_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13439__A _13898_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11389_ _11405_/CLK line[1] vssd1 vssd1 vccd1 vccd1 _11390_/A sky130_fd_sc_hd__dfxtp_1
X_13128_ _13128_/A _13159_/Y vssd1 vssd1 vccd1 vccd1 _13688_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13158__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13059_ _13085_/CLK line[11] vssd1 vssd1 vccd1 vccd1 _13060_/A sky130_fd_sc_hd__dfxtp_1
X_05950_ _05980_/CLK line[80] vssd1 vssd1 vccd1 vccd1 _05951_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_DATA\[20\].CLKBUF\[3\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05881_ _05881_/A _05914_/Y vssd1 vssd1 vccd1 vccd1 _13721_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_39_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11109__D line[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07620_ _07620_/A _07629_/Y vssd1 vssd1 vccd1 vccd1 _13780_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_93_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09802__D line[58] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07551_ _07555_/CLK line[39] vssd1 vssd1 vccd1 vccd1 _07552_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10948__D line[56] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13324__D line[118] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06502_ _06502_/A _06509_/Y vssd1 vssd1 vccd1 vccd1 _13782_/Z sky130_fd_sc_hd__ebufn_2
X_07482_ _07482_/A _07489_/Y vssd1 vssd1 vccd1 vccd1 _13642_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08418__D line[51] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09221_ _09235_/CLK line[34] vssd1 vssd1 vccd1 vccd1 _09222_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_210_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06433_ _06435_/CLK line[40] vssd1 vssd1 vccd1 vccd1 _06434_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_210_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09152_ _09152_/A _09169_/Y vssd1 vssd1 vccd1 vccd1 _13632_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09099__A _13915_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06364_ _06364_/A _06369_/Y vssd1 vssd1 vccd1 vccd1 _13644_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_159_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08103_ _08115_/CLK line[35] vssd1 vssd1 vccd1 vccd1 _08104_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_147_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[4\].VALID\[8\].FF OVHB\[4\].V/CLK A[15] vssd1 vssd1 vccd1 vccd1 OVHB\[4\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_05315_ _05315_/CLK line[41] vssd1 vssd1 vccd1 vccd1 _05316_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10683__D line[77] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09083_ _09095_/CLK line[99] vssd1 vssd1 vccd1 vccd1 _09084_/A sky130_fd_sc_hd__dfxtp_1
X_06295_ _06295_/CLK line[105] vssd1 vssd1 vccd1 vccd1 _06296_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.M\[3\].MUX\[4\]_A2 _13797_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05777__D line[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08034_ _08034_/A _08049_/Y vssd1 vssd1 vccd1 vccd1 _13634_/Z sky130_fd_sc_hd__ebufn_2
X_05246_ _05246_/A _05249_/Y vssd1 vssd1 vccd1 vccd1 _13646_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_162_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05177_ _05177_/CLK _05178_/X vssd1 vssd1 vccd1 vccd1 _05175_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__07992__D line[127] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09035__TE_B _09064_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09985_ _10005_/CLK line[14] vssd1 vssd1 vccd1 vccd1 _09986_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_67_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08936_ _08936_/A _08959_/Y vssd1 vssd1 vccd1 vccd1 _13696_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_130_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08867_ _08885_/CLK line[15] vssd1 vssd1 vccd1 vccd1 _08868_/A sky130_fd_sc_hd__dfxtp_1
X_07818_ _07818_/A _07839_/Y vssd1 vssd1 vccd1 vccd1 _13698_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[21\].VALID\[3\].FF_D A[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05017__D line[47] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08798_ _08798_/A _08819_/Y vssd1 vssd1 vccd1 vccd1 _13838_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_44_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MUX.M\[1\].MUX\[0\]_A3 _13854_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10858__D line[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07749_ _07765_/CLK line[1] vssd1 vssd1 vccd1 vccd1 _07750_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_25_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13234__D line[91] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10760_ _10760_/A _10779_/Y vssd1 vssd1 vccd1 vccd1 _13840_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_16_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07232__D line[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09419_ _09445_/CLK line[11] vssd1 vssd1 vccd1 vccd1 _09420_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_200_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10691_ _10705_/CLK line[66] vssd1 vssd1 vccd1 vccd1 _10692_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[14\].VALID\[7\].FF_D A[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12430_ _12430_/A _12459_/Y vssd1 vssd1 vccd1 vccd1 _13830_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_32_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12361_ _12385_/CLK line[76] vssd1 vssd1 vccd1 vccd1 _12362_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_165_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09159__D line[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[5\].VALID\[7\].TOBUF OVHB\[5\].VALID\[7\].FF/Q OVHB\[5\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/A2 sky130_fd_sc_hd__ebufn_2
XFILLER_138_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11312_ _11312_/A _11339_/Y vssd1 vssd1 vccd1 vccd1 _13832_/Z sky130_fd_sc_hd__ebufn_2
X_12292_ _12292_/A _12319_/Y vssd1 vssd1 vccd1 vccd1 _13692_/Z sky130_fd_sc_hd__ebufn_2
X_11243_ _11265_/CLK line[77] vssd1 vssd1 vccd1 vccd1 _11244_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_180_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11174_ _11174_/A _11199_/Y vssd1 vssd1 vccd1 vccd1 _13694_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13409__D line[43] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12313__D line[40] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10125_ _10145_/CLK line[78] vssd1 vssd1 vccd1 vccd1 _10126_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_DATA\[19\].CLKBUF\[4\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07407__D line[101] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[11\].VALID\[11\].FF_D A[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10056_ _10056_/A _10079_/Y vssd1 vssd1 vccd1 vccd1 _13696_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_87_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13815_ _13815_/A _13824_/Y vssd1 vssd1 vccd1 vccd1 _13815_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_189_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13746_ _13750_/CLK line[55] vssd1 vssd1 vccd1 vccd1 _13747_/A sky130_fd_sc_hd__dfxtp_1
X_10958_ _10958_/A _10989_/Y vssd1 vssd1 vccd1 vccd1 _13758_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07142__D line[122] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13677_ _13677_/A _13684_/Y vssd1 vssd1 vccd1 vccd1 _13677_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_188_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10889_ _10915_/CLK line[43] vssd1 vssd1 vccd1 vccd1 _10890_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_31_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06981__D line[34] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12628_ _12630_/CLK line[56] vssd1 vssd1 vccd1 vccd1 _12629_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[21\].VALID\[10\].FF_D A[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11599__D line[97] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12559_ _12559_/A _12564_/Y vssd1 vssd1 vccd1 vccd1 _13679_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_129_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09069__D line[107] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05100_ _05100_/A _05109_/Y vssd1 vssd1 vccd1 vccd1 _13780_/Z sky130_fd_sc_hd__ebufn_2
X_06080_ _06080_/A _06089_/Y vssd1 vssd1 vccd1 vccd1 _13640_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_129_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[13\].VALID\[0\].FF OVHB\[13\].V/CLK A[7] vssd1 vssd1 vccd1 vccd1 OVHB\[13\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_05031_ _05035_/CLK line[39] vssd1 vssd1 vccd1 vccd1 _05032_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[30\].VALID\[4\].FF OVHB\[30\].V/CLK A[11] vssd1 vssd1 vccd1 vccd1 OVHB\[30\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12073__A _13934_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12223__D line[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09770_ _09770_/A _09799_/Y vssd1 vssd1 vccd1 vccd1 _13690_/Z sky130_fd_sc_hd__ebufn_2
X_06982_ _06982_/A _06999_/Y vssd1 vssd1 vccd1 vccd1 _13702_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_113_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[11\].VALID\[11\].FF OVHB\[11\].V/CLK A[18] vssd1 vssd1 vccd1 vccd1 OVHB\[11\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07317__D line[74] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08721_ _08745_/CLK line[76] vssd1 vssd1 vccd1 vccd1 _08722_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06221__D line[71] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XOVHB\[12\].VALID\[2\].TOBUF OVHB\[12\].VALID\[2\].FF/Q OVHB\[12\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04930_/B2 sky130_fd_sc_hd__ebufn_2
X_05933_ _05945_/CLK line[67] vssd1 vssd1 vccd1 vccd1 _05934_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_66_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08652_ _08652_/A _08679_/Y vssd1 vssd1 vccd1 vccd1 _13692_/Z sky130_fd_sc_hd__ebufn_2
X_05864_ _05864_/A _05879_/Y vssd1 vssd1 vccd1 vccd1 _13704_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_93_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09532__D line[63] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07603_ _07625_/CLK line[77] vssd1 vssd1 vccd1 vccd1 _07604_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08583_ _08605_/CLK line[13] vssd1 vssd1 vccd1 vccd1 _08584_/A sky130_fd_sc_hd__dfxtp_1
X_05795_ _05805_/CLK line[4] vssd1 vssd1 vccd1 vccd1 _05796_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_35_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07534_ _07534_/A _07559_/Y vssd1 vssd1 vccd1 vccd1 _13694_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08148__D line[56] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[27\].VALID\[7\].FF_D A[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07465_ _07485_/CLK line[14] vssd1 vssd1 vccd1 vccd1 _07466_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12248__A _13935_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09204_ _13916_/X vssd1 vssd1 vccd1 vccd1 _09204_/Y sky130_fd_sc_hd__inv_2
X_06416_ _06416_/A _06439_/Y vssd1 vssd1 vccd1 vccd1 _13696_/Z sky130_fd_sc_hd__ebufn_2
X_07396_ _07396_/A _07419_/Y vssd1 vssd1 vccd1 vccd1 _13836_/Z sky130_fd_sc_hd__ebufn_2
X_09135_ _09165_/CLK line[0] vssd1 vssd1 vccd1 vccd1 _09136_/A sky130_fd_sc_hd__dfxtp_1
X_06347_ _06365_/CLK line[15] vssd1 vssd1 vccd1 vccd1 _06348_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_136_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09066_ _09066_/A _09099_/Y vssd1 vssd1 vccd1 vccd1 _13826_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[29\].VALID\[5\].FF OVHB\[29\].V/CLK A[12] vssd1 vssd1 vccd1 vccd1 OVHB\[29\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_06278_ _06278_/A _06299_/Y vssd1 vssd1 vccd1 vccd1 _13838_/Z sky130_fd_sc_hd__ebufn_2
X_08017_ _08045_/CLK line[10] vssd1 vssd1 vccd1 vccd1 _08018_/A sky130_fd_sc_hd__dfxtp_1
X_05229_ _05245_/CLK line[1] vssd1 vssd1 vccd1 vccd1 _05230_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MUX.M\[2\].MUX\[5\]_A0 _13673_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09707__D line[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09968_ _09970_/CLK line[120] vssd1 vssd1 vccd1 vccd1 _09969_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[11\].VALID\[2\].FF OVHB\[11\].V/CLK A[9] vssd1 vssd1 vccd1 vccd1 OVHB\[11\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06131__D line[44] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08919_ _08919_/A _08924_/Y vssd1 vssd1 vccd1 vccd1 _13679_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_94_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09899_ _09899_/A _09904_/Y vssd1 vssd1 vccd1 vccd1 _13819_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11972__D line[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11930_ _11930_/CLK line[121] vssd1 vssd1 vccd1 vccd1 _11931_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_206_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05970__D line[84] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10588__D line[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11861_ _11861_/A _11864_/Y vssd1 vssd1 vccd1 vccd1 _13821_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_205_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13600_ _13610_/CLK line[116] vssd1 vssd1 vccd1 vccd1 _13601_/A sky130_fd_sc_hd__dfxtp_1
X_10812_ _10812_/CLK _10813_/X vssd1 vssd1 vccd1 vccd1 _10810_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__08058__D line[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11792_ _11792_/CLK _11793_/X vssd1 vssd1 vccd1 vccd1 _11790_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA_MUX.M\[0\].MUX\[1\]_A1 _13700_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13531_ _13531_/A _13544_/Y vssd1 vssd1 vccd1 vccd1 _13811_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_186_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10743_ _13924_/X wr vssd1 vssd1 vccd1 vccd1 _10743_/X sky130_fd_sc_hd__and2_1
XFILLER_13_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07897__D line[69] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DECH.DEC0.AND1_B A_h[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13462_ _13470_/CLK line[53] vssd1 vssd1 vccd1 vccd1 _13463_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_186_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10674_ _13924_/X vssd1 vssd1 vccd1 vccd1 _10674_/Y sky130_fd_sc_hd__inv_2
X_12413_ _12413_/A _12424_/Y vssd1 vssd1 vccd1 vccd1 _13813_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_127_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13393_ _13393_/A _13404_/Y vssd1 vssd1 vccd1 vccd1 _13673_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_154_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11212__D line[63] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12344_ _12350_/CLK line[54] vssd1 vssd1 vccd1 vccd1 _12345_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06306__D line[124] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05210__D line[121] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[8\].VALID\[12\].TOBUF OVHB\[8\].VALID\[12\].FF/Q OVHB\[8\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04929_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_175_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[8\].VALID\[2\].FF_D A[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12275_ _12275_/A _12284_/Y vssd1 vssd1 vccd1 vccd1 _13675_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_107_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11226_ _11230_/CLK line[55] vssd1 vssd1 vccd1 vccd1 _11227_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08521__D line[98] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13139__D line[33] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11157_ _11157_/A _11164_/Y vssd1 vssd1 vccd1 vccd1 _13677_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_110_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[27\].VALID\[7\].FF OVHB\[27\].V/CLK A[14] vssd1 vssd1 vccd1 vccd1 OVHB\[27\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_68_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10108_ _10110_/CLK line[56] vssd1 vssd1 vccd1 vccd1 _10109_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12978__D line[88] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11088_ _11090_/CLK line[120] vssd1 vssd1 vccd1 vccd1 _11089_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_208_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[26\].VALID\[14\].FF_D A[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10039_ _10039_/A _10044_/Y vssd1 vssd1 vccd1 vccd1 _13679_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[6\].VALID\[13\].FF OVHB\[6\].V/CLK A[20] vssd1 vssd1 vccd1 vccd1 OVHB\[6\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_208_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05880__D line[48] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[17\].CLKBUF\[6\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05580_ _05580_/A _05599_/Y vssd1 vssd1 vccd1 vccd1 _13700_/Z sky130_fd_sc_hd__ebufn_2
X_13729_ _13729_/A _13754_/Y vssd1 vssd1 vccd1 vccd1 _13729_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13602__D line[117] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[1\].VALID\[11\].TOBUF OVHB\[1\].VALID\[11\].FF/Q OVHB\[1\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04915_/B2 sky130_fd_sc_hd__ebufn_2
X_07250_ _07250_/A _07279_/Y vssd1 vssd1 vccd1 vccd1 _13690_/Z sky130_fd_sc_hd__ebufn_2
X_06201_ _06225_/CLK line[76] vssd1 vssd1 vccd1 vccd1 _06202_/A sky130_fd_sc_hd__dfxtp_1
X_07181_ _07205_/CLK line[12] vssd1 vssd1 vccd1 vccd1 _07182_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[10\].VALID\[7\].TOBUF OVHB\[10\].VALID\[7\].FF/Q OVHB\[10\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/A2 sky130_fd_sc_hd__ebufn_2
X_06132_ _06132_/A _06159_/Y vssd1 vssd1 vccd1 vccd1 _13692_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05120__D line[94] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDATA\[19\].CLKBUF\[1\] clk vssd1 vssd1 vccd1 vccd1 _07802_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_133_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10961__D line[76] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06063_ _06085_/CLK line[13] vssd1 vssd1 vccd1 vccd1 _06064_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_144_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05014_ _05014_/A _05039_/Y vssd1 vssd1 vccd1 vccd1 _13694_/Z sky130_fd_sc_hd__ebufn_2
X_09822_ _09830_/CLK line[53] vssd1 vssd1 vccd1 vccd1 _09823_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_59_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07047__D line[79] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09753_ _09753_/A _09764_/Y vssd1 vssd1 vccd1 vccd1 _13673_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12888__D line[61] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06965_ _06995_/CLK line[32] vssd1 vssd1 vccd1 vccd1 _06966_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_74_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__04968__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08704_ _08710_/CLK line[54] vssd1 vssd1 vccd1 vccd1 _08705_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06886__D line[119] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05916_ _05916_/A _05949_/Y vssd1 vssd1 vccd1 vccd1 _13756_/Z sky130_fd_sc_hd__ebufn_2
X_09684_ _09690_/CLK line[118] vssd1 vssd1 vccd1 vccd1 _09685_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_67_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06896_ _06896_/A _06929_/Y vssd1 vssd1 vccd1 vccd1 _13616_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09262__D line[53] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[18\].VALID\[11\].FF_D A[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08635_ _08635_/A _08644_/Y vssd1 vssd1 vccd1 vccd1 _13675_/Z sky130_fd_sc_hd__ebufn_2
X_05847_ _05875_/CLK line[42] vssd1 vssd1 vccd1 vccd1 _05848_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10201__D line[98] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[25\].VALID\[9\].FF OVHB\[25\].V/CLK A[16] vssd1 vssd1 vccd1 vccd1 OVHB\[25\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08566_ _08570_/CLK line[119] vssd1 vssd1 vccd1 vccd1 _08567_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05778_ _05778_/A _05809_/Y vssd1 vssd1 vccd1 vccd1 _13618_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07517_ _07517_/A _07524_/Y vssd1 vssd1 vccd1 vccd1 _13677_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08497_ _08497_/A _08504_/Y vssd1 vssd1 vccd1 vccd1 _13817_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13512__D line[90] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07448_ _07450_/CLK line[120] vssd1 vssd1 vccd1 vccd1 _07449_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_196_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07510__D line[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12128__D line[83] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07379_ _07379_/A _07384_/Y vssd1 vssd1 vccd1 vccd1 _13819_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_108_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09118_ _09130_/CLK line[115] vssd1 vssd1 vccd1 vccd1 _09119_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_89_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[28\].VALID\[10\].FF_D A[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10390_ _10390_/CLK line[57] vssd1 vssd1 vccd1 vccd1 _10391_/A sky130_fd_sc_hd__dfxtp_1
X_09049_ _09049_/A _09064_/Y vssd1 vssd1 vccd1 vccd1 _13809_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_124_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09437__D line[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12060_ _12070_/CLK line[52] vssd1 vssd1 vccd1 vccd1 _12061_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_104_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11011_ _11011_/A _11024_/Y vssd1 vssd1 vccd1 vccd1 _13811_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_89_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12962_ _12980_/CLK line[95] vssd1 vssd1 vccd1 vccd1 _12963_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06796__D line[92] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09172__D line[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11913_ _11913_/A _11934_/Y vssd1 vssd1 vccd1 vccd1 _13873_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_18_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[19\].VALID\[2\].TOBUF OVHB\[19\].VALID\[2\].FF/Q OVHB\[19\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04930_/B2 sky130_fd_sc_hd__ebufn_2
X_12893_ _12893_/A _12914_/Y vssd1 vssd1 vccd1 vccd1 _13733_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11844_ _11860_/CLK line[81] vssd1 vssd1 vccd1 vccd1 _11845_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_61_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09900__D line[89] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11775_ _11775_/A _11794_/Y vssd1 vssd1 vccd1 vccd1 _13735_/Z sky130_fd_sc_hd__ebufn_2
X_10726_ _10740_/CLK line[82] vssd1 vssd1 vccd1 vccd1 _10727_/A sky130_fd_sc_hd__dfxtp_1
X_13514_ _13540_/CLK line[91] vssd1 vssd1 vccd1 vccd1 _13515_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07420__D line[112] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13445_ _13445_/A _13474_/Y vssd1 vssd1 vccd1 vccd1 _13725_/Z sky130_fd_sc_hd__ebufn_2
X_10657_ _10657_/A _10674_/Y vssd1 vssd1 vccd1 vccd1 _13737_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[24\].VALID\[13\].TOBUF OVHB\[24\].VALID\[13\].FF/Q OVHB\[24\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04916_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__06036__D line[114] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13376_ _13400_/CLK line[28] vssd1 vssd1 vccd1 vccd1 _13377_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_127_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10588_ _10600_/CLK line[19] vssd1 vssd1 vccd1 vccd1 _10589_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06614__A _13904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11877__D line[111] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12327_ _12327_/A _12354_/Y vssd1 vssd1 vccd1 vccd1 _13727_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_142_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09347__D line[106] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05875__D line[41] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06333__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08251__D line[103] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12258_ _12280_/CLK line[29] vssd1 vssd1 vccd1 vccd1 _12259_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_130_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[30\].VALID\[6\].FF_D A[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11209_ _11209_/A _11234_/Y vssd1 vssd1 vccd1 vccd1 _13729_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_96_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12189_ _12189_/A _12214_/Y vssd1 vssd1 vccd1 vccd1 _13869_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_122_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12501__D line[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06750_ _06750_/CLK line[57] vssd1 vssd1 vccd1 vccd1 _06751_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_49_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05701_ _05701_/A _05704_/Y vssd1 vssd1 vccd1 vccd1 _13821_/Z sky130_fd_sc_hd__ebufn_2
X_06681_ _06681_/A _06684_/Y vssd1 vssd1 vccd1 vccd1 _13681_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_63_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11117__D line[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08420_ _08430_/CLK line[52] vssd1 vssd1 vccd1 vccd1 _08421_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_24_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05632_ _05632_/CLK _05633_/X vssd1 vssd1 vccd1 vccd1 _05630_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_91_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09810__D line[62] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08351_ _08351_/A _08364_/Y vssd1 vssd1 vccd1 vccd1 _13671_/Z sky130_fd_sc_hd__ebufn_2
X_05563_ _13901_/X wr vssd1 vssd1 vccd1 vccd1 _05563_/X sky130_fd_sc_hd__and2_1
X_07302_ _07310_/CLK line[53] vssd1 vssd1 vccd1 vccd1 _07303_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06508__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08426__D line[55] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08282_ _08290_/CLK line[117] vssd1 vssd1 vccd1 vccd1 _08283_/A sky130_fd_sc_hd__dfxtp_1
X_05494_ _13900_/X vssd1 vssd1 vccd1 vccd1 _05494_/Y sky130_fd_sc_hd__inv_2
XFILLER_149_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07233_ _07233_/A _07244_/Y vssd1 vssd1 vccd1 vccd1 _13673_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[0\].V_RESET_B rst_n vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[25\].VALID\[1\].TOBUF OVHB\[25\].VALID\[1\].FF/Q OVHB\[25\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04926_/B2 sky130_fd_sc_hd__ebufn_2
X_07164_ _07170_/CLK line[118] vssd1 vssd1 vccd1 vccd1 _07165_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.SEL1BUF\[2\]_A A[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06115_ _06115_/A _06124_/Y vssd1 vssd1 vccd1 vccd1 _13675_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10691__D line[66] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07095_ _07095_/A _07104_/Y vssd1 vssd1 vccd1 vccd1 _13815_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[26\].CG_CLK clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05785__D line[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08161__D line[76] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[1\].CGAND_B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[20\].CGAND_A _13913_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06046_ _06050_/CLK line[119] vssd1 vssd1 vccd1 vccd1 _06047_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[2\].VALID\[11\].FF OVHB\[2\].V/CLK A[18] vssd1 vssd1 vccd1 vccd1 OVHB\[2\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_99_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MUX.M\[2\].MUX\[2\]_A3 _13877_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[5\].CGAND_A _13936_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09805_ _09805_/A _09834_/Y vssd1 vssd1 vccd1 vccd1 _13725_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__04919__B1 A_h[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07997_ _07997_/A _08014_/Y vssd1 vssd1 vccd1 vccd1 _13877_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_75_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06948_ _06960_/CLK line[19] vssd1 vssd1 vccd1 vccd1 _06949_/A sky130_fd_sc_hd__dfxtp_1
X_09736_ _09760_/CLK line[28] vssd1 vssd1 vccd1 vccd1 _09737_/A sky130_fd_sc_hd__dfxtp_1
X_09667_ _09667_/A _09694_/Y vssd1 vssd1 vccd1 vccd1 _13867_/Z sky130_fd_sc_hd__ebufn_2
X_06879_ _06879_/A _06894_/Y vssd1 vssd1 vccd1 vccd1 _13879_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11027__D line[106] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08618_ _08640_/CLK line[29] vssd1 vssd1 vccd1 vccd1 _08619_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_82_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09598_ _09620_/CLK line[93] vssd1 vssd1 vccd1 vccd1 _09599_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_188_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05025__D line[36] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10866__D line[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08549_ _08549_/A _08574_/Y vssd1 vssd1 vccd1 vccd1 _13869_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13242__D line[95] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11560_ _11580_/CLK line[94] vssd1 vssd1 vccd1 vccd1 _11561_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08336__D line[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07240__D line[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_DATA\[30\].CLKBUF\[1\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10511_ _10511_/A _10534_/Y vssd1 vssd1 vccd1 vccd1 _13871_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11491_ _11491_/A _11514_/Y vssd1 vssd1 vccd1 vccd1 _13731_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[4\].VALID\[5\].FF_D A[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13230_ _13260_/CLK line[80] vssd1 vssd1 vccd1 vccd1 _13231_/A sky130_fd_sc_hd__dfxtp_1
X_10442_ _10460_/CLK line[95] vssd1 vssd1 vccd1 vccd1 _10443_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_40_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13161_ _13161_/A _13194_/Y vssd1 vssd1 vccd1 vccd1 _13721_/Z sky130_fd_sc_hd__ebufn_2
X_10373_ _10373_/A _10394_/Y vssd1 vssd1 vccd1 vccd1 _13733_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[17\].VALID\[7\].TOBUF OVHB\[17\].VALID\[7\].FF/Q OVHB\[17\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/A2 sky130_fd_sc_hd__ebufn_2
XFILLER_191_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12112_ _12140_/CLK line[90] vssd1 vssd1 vccd1 vccd1 _12113_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_108_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13092_ _13120_/CLK line[26] vssd1 vssd1 vccd1 vccd1 _13093_/A sky130_fd_sc_hd__dfxtp_1
X_12043_ _12043_/A _12074_/Y vssd1 vssd1 vccd1 vccd1 _13723_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10106__D line[55] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XOVHB\[31\].VALID\[0\].TOBUF OVHB\[31\].VALID\[0\].FF/Q OVHB\[31\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04924_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__13417__D line[47] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07415__D line[105] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12945_ _12945_/CLK line[73] vssd1 vssd1 vccd1 vccd1 _12946_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_61_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12876_ _12876_/A _12879_/Y vssd1 vssd1 vccd1 vccd1 _13716_/Z sky130_fd_sc_hd__ebufn_2
X_11827_ _11827_/CLK _11828_/X vssd1 vssd1 vccd1 vccd1 _11825_/CLK sky130_fd_sc_hd__dlclkp_1
X_11758_ _13927_/X wr vssd1 vssd1 vccd1 vccd1 _11758_/X sky130_fd_sc_hd__and2_1
XANTENNA__07150__D line[126] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10709_ _13924_/X vssd1 vssd1 vccd1 vccd1 _10709_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12991__D line[108] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11689_ _13927_/X vssd1 vssd1 vccd1 vccd1 _11689_/Y sky130_fd_sc_hd__inv_2
XFILLER_146_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13428_ _13428_/A _13439_/Y vssd1 vssd1 vccd1 vccd1 _13708_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_139_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XOVHB\[16\].VALID\[11\].FF OVHB\[16\].V/CLK A[18] vssd1 vssd1 vccd1 vccd1 OVHB\[16\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_13359_ _13365_/CLK line[6] vssd1 vssd1 vccd1 vccd1 _13360_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_182_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09077__D line[111] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06998__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10016__D line[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07920_ _07940_/CLK line[94] vssd1 vssd1 vccd1 vccd1 _07921_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_96_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[19\].VALID\[2\].FF_D A[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07851_ _07851_/A _07874_/Y vssd1 vssd1 vccd1 vccd1 _13731_/Z sky130_fd_sc_hd__ebufn_2
X_06802_ _06820_/CLK line[95] vssd1 vssd1 vccd1 vccd1 _06803_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__04949__D line[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12231__D line[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07782_ _07800_/CLK line[31] vssd1 vssd1 vccd1 vccd1 _07783_/A sky130_fd_sc_hd__dfxtp_1
X_04994_ _05000_/CLK line[22] vssd1 vssd1 vccd1 vccd1 _04995_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07325__D line[78] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[23\].VALID\[6\].TOBUF OVHB\[23\].VALID\[6\].FF/Q OVHB\[23\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04923_/A2 sky130_fd_sc_hd__ebufn_2
X_09521_ _09521_/A _09554_/Y vssd1 vssd1 vccd1 vccd1 _13721_/Z sky130_fd_sc_hd__ebufn_2
X_06733_ _06733_/A _06754_/Y vssd1 vssd1 vccd1 vccd1 _13733_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_37_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09452_ _09480_/CLK line[26] vssd1 vssd1 vccd1 vccd1 _09453_/A sky130_fd_sc_hd__dfxtp_1
X_06664_ _06680_/CLK line[17] vssd1 vssd1 vccd1 vccd1 _06665_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_36_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09540__D line[52] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08403_ _08403_/A _08434_/Y vssd1 vssd1 vccd1 vccd1 _13723_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05423__A _13900_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05615_ _05615_/A _05634_/Y vssd1 vssd1 vccd1 vccd1 _13735_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_169_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09383_ _09383_/A _09414_/Y vssd1 vssd1 vccd1 vccd1 _13863_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_51_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06595_ _06595_/A _06614_/Y vssd1 vssd1 vccd1 vccd1 _13875_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_196_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_DATA\[29\].CLKBUF\[2\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08334_ _08360_/CLK line[27] vssd1 vssd1 vccd1 vccd1 _08335_/A sky130_fd_sc_hd__dfxtp_1
X_05546_ _05560_/CLK line[18] vssd1 vssd1 vccd1 vccd1 _05547_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.M\[3\].MUX\[7\]_A0 _13663_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08265_ _08265_/A _08294_/Y vssd1 vssd1 vccd1 vccd1 _13865_/Z sky130_fd_sc_hd__ebufn_2
X_05477_ _05477_/A _05494_/Y vssd1 vssd1 vccd1 vccd1 _13877_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_137_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07216_ _07240_/CLK line[28] vssd1 vssd1 vccd1 vccd1 _07217_/A sky130_fd_sc_hd__dfxtp_1
X_08196_ _08220_/CLK line[92] vssd1 vssd1 vccd1 vccd1 _08197_/A sky130_fd_sc_hd__dfxtp_1
X_07147_ _07147_/A _07174_/Y vssd1 vssd1 vccd1 vccd1 _13867_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12406__D line[82] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07078_ _07100_/CLK line[93] vssd1 vssd1 vccd1 vccd1 _07079_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_133_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12703__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06029_ _06029_/A _06054_/Y vssd1 vssd1 vccd1 vccd1 _13869_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09715__D line[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_MUX.M\[1\].MUX\[3\]_A1 _13690_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09719_ _09725_/CLK line[6] vssd1 vssd1 vccd1 vccd1 _09720_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_16_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10991_ _10991_/A _11024_/Y vssd1 vssd1 vccd1 vccd1 _13791_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11980__D line[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[1\].CGAND _13932_/X wr vssd1 vssd1 vccd1 vccd1 OVHB\[1\].CGAND/X sky130_fd_sc_hd__and2_4
X_12730_ _12730_/A _12739_/Y vssd1 vssd1 vccd1 vccd1 _13850_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_16_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09450__D line[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10596__D line[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12661_ _12665_/CLK line[71] vssd1 vssd1 vccd1 vccd1 _12662_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11612_ _11612_/A _11619_/Y vssd1 vssd1 vccd1 vccd1 _13852_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08066__D line[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12592_ _12592_/A _12599_/Y vssd1 vssd1 vccd1 vccd1 _13712_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08644__A _13914_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11543_ _11545_/CLK line[72] vssd1 vssd1 vccd1 vccd1 _11544_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_DATA\[2\].CLKBUF\[1\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08363__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11474_ _11474_/A _11479_/Y vssd1 vssd1 vccd1 vccd1 _13714_/Z sky130_fd_sc_hd__ebufn_2
X_13213_ _13225_/CLK line[67] vssd1 vssd1 vccd1 vccd1 _13214_/A sky130_fd_sc_hd__dfxtp_1
X_10425_ _10425_/CLK line[73] vssd1 vssd1 vccd1 vccd1 _10426_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11220__D line[52] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13144_ _13144_/A _13159_/Y vssd1 vssd1 vccd1 vccd1 _13704_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06314__D line[113] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDATA\[9\].CLKBUF\[2\] clk vssd1 vssd1 vccd1 vccd1 _13717_/CLK sky130_fd_sc_hd__clkbuf_4
X_10356_ _10356_/A _10359_/Y vssd1 vssd1 vccd1 vccd1 _13716_/Z sky130_fd_sc_hd__ebufn_2
X_13075_ _13085_/CLK line[4] vssd1 vssd1 vccd1 vccd1 _13076_/A sky130_fd_sc_hd__dfxtp_1
X_10287_ _10287_/CLK _10288_/X vssd1 vssd1 vccd1 vccd1 _10285_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__09625__D line[96] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12026_ _12026_/A _12039_/Y vssd1 vssd1 vccd1 vccd1 _13706_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13147__D line[37] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08819__A _13914_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13977_ _13982_/C _13982_/A _13982_/B _13982_/D vssd1 vssd1 vccd1 vccd1 _13977_/X
+ sky130_fd_sc_hd__and4bb_4
XFILLER_18_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08538__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12928_ _12928_/A _12949_/Y vssd1 vssd1 vccd1 vccd1 _13768_/Z sky130_fd_sc_hd__ebufn_2
X_12859_ _12875_/CLK line[33] vssd1 vssd1 vccd1 vccd1 _12860_/A sky130_fd_sc_hd__dfxtp_1
X_05400_ _05420_/CLK line[94] vssd1 vssd1 vccd1 vccd1 _05401_/A sky130_fd_sc_hd__dfxtp_1
X_06380_ _06400_/CLK line[30] vssd1 vssd1 vccd1 vccd1 _06381_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_33_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05331_ _05331_/A _05354_/Y vssd1 vssd1 vccd1 vccd1 _13731_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_147_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XOVHB\[14\].VALID\[11\].TOBUF OVHB\[14\].VALID\[11\].FF/Q OVHB\[14\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04915_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__13610__D line[121] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XDATA\[29\].CLKBUF\[6\] clk vssd1 vssd1 vccd1 vccd1 _11057_/CLK sky130_fd_sc_hd__clkbuf_4
X_08050_ _08080_/CLK line[16] vssd1 vssd1 vccd1 vccd1 _08051_/A sky130_fd_sc_hd__dfxtp_1
X_05262_ _05280_/CLK line[31] vssd1 vssd1 vccd1 vccd1 _05263_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08704__D line[54] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__04916__A2_N _04916_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07001_ _07001_/A _07034_/Y vssd1 vssd1 vccd1 vccd1 _13721_/Z sky130_fd_sc_hd__ebufn_2
X_05193_ _05193_/A _05214_/Y vssd1 vssd1 vccd1 vccd1 _13873_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11130__D line[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10324__A _13923_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08952_ _08952_/A _08959_/Y vssd1 vssd1 vccd1 vccd1 _13712_/Z sky130_fd_sc_hd__ebufn_2
X_07903_ _07905_/CLK line[72] vssd1 vssd1 vccd1 vccd1 _07904_/A sky130_fd_sc_hd__dfxtp_1
X_08883_ _08885_/CLK line[8] vssd1 vssd1 vccd1 vccd1 _08884_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10043__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13057__D line[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07834_ _07834_/A _07839_/Y vssd1 vssd1 vccd1 vccd1 _13714_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_29_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07055__D line[68] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07765_ _07765_/CLK line[9] vssd1 vssd1 vccd1 vccd1 _07766_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12896__D line[50] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_04977_ _04977_/A _05004_/Y vssd1 vssd1 vccd1 vccd1 _13657_/Z sky130_fd_sc_hd__ebufn_2
X_09504_ _09504_/A _09519_/Y vssd1 vssd1 vccd1 vccd1 _13704_/Z sky130_fd_sc_hd__ebufn_2
X_06716_ _06716_/A _06719_/Y vssd1 vssd1 vccd1 vccd1 _13716_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_24_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07696_ _07696_/A _07699_/Y vssd1 vssd1 vccd1 vccd1 _13856_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09270__D line[57] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09435_ _09445_/CLK line[4] vssd1 vssd1 vccd1 vccd1 _09436_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_24_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06647_ _06647_/CLK _06648_/X vssd1 vssd1 vccd1 vccd1 _06645_/CLK sky130_fd_sc_hd__dlclkp_1
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11305__D line[96] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09366_ _09366_/A _09379_/Y vssd1 vssd1 vccd1 vccd1 _13846_/Z sky130_fd_sc_hd__ebufn_2
X_06578_ _13904_/X wr vssd1 vssd1 vccd1 vccd1 _06578_/X sky130_fd_sc_hd__and2_1
XANTENNA_OVHB\[0\].VALID\[8\].FF_D A[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05303__D line[35] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08317_ _08325_/CLK line[5] vssd1 vssd1 vccd1 vccd1 _08318_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_166_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05529_ _13901_/X vssd1 vssd1 vccd1 vccd1 _05529_/Y sky130_fd_sc_hd__inv_2
XFILLER_166_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09297_ _09305_/CLK line[69] vssd1 vssd1 vccd1 vccd1 _09298_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_138_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13520__D line[94] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08614__D line[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08248_ _08248_/A _08259_/Y vssd1 vssd1 vccd1 vccd1 _13848_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10218__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12136__D line[87] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08179_ _08185_/CLK line[70] vssd1 vssd1 vccd1 vccd1 _08180_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[27\].CLKBUF\[4\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10210_ _10210_/A _10219_/Y vssd1 vssd1 vccd1 vccd1 _13850_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_97_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XDATA\[28\].CLKBUF\[3\] clk vssd1 vssd1 vccd1 vccd1 _10672_/CLK sky130_fd_sc_hd__clkbuf_4
X_11190_ _11190_/A _11199_/Y vssd1 vssd1 vccd1 vccd1 _13710_/Z sky130_fd_sc_hd__ebufn_2
X_10141_ _10145_/CLK line[71] vssd1 vssd1 vccd1 vccd1 _10142_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_79_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09445__D line[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10072_ _10072_/A _10079_/Y vssd1 vssd1 vccd1 vccd1 _13712_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_48_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13900_ _13905_/C _13905_/A _13905_/B _13905_/D vssd1 vssd1 vccd1 vccd1 _13900_/X
+ sky130_fd_sc_hd__and4bb_4
XFILLER_208_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13831_ _13855_/CLK line[108] vssd1 vssd1 vccd1 vccd1 _13832_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[5\].VALID\[3\].TOBUF OVHB\[5\].VALID\[3\].FF/Q OVHB\[5\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04919_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_35_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[3\].VALID\[14\].FF_D A[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10974_ _10974_/A _10989_/Y vssd1 vssd1 vccd1 vccd1 _13774_/Z sky130_fd_sc_hd__ebufn_2
X_13762_ _13762_/A _13789_/Y vssd1 vssd1 vccd1 vccd1 _13762_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09180__D line[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06159__A _13903_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12713_ _12735_/CLK line[109] vssd1 vssd1 vccd1 vccd1 _12714_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_71_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13693_ _13715_/CLK line[45] vssd1 vssd1 vccd1 vccd1 _13694_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_31_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[21\].VALID\[0\].FF OVHB\[21\].V/CLK A[7] vssd1 vssd1 vccd1 vccd1 OVHB\[21\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12644_ _12644_/A _12669_/Y vssd1 vssd1 vccd1 vccd1 _13764_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_176_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12575_ _12595_/CLK line[46] vssd1 vssd1 vccd1 vccd1 _12576_/A sky130_fd_sc_hd__dfxtp_1
XPHY_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[22\].VALID\[1\].FF_D A[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11526_ _11526_/A _11549_/Y vssd1 vssd1 vccd1 vccd1 _13766_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_7_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12046__D line[60] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11457_ _11475_/CLK line[47] vssd1 vssd1 vccd1 vccd1 _11458_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[21\].CG clk OVHB\[21\].CGAND/X vssd1 vssd1 vccd1 vccd1 OVHB\[21\].V/CLK sky130_fd_sc_hd__dlclkp_1
X_10408_ _10408_/A _10429_/Y vssd1 vssd1 vccd1 vccd1 _13768_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06044__D line[118] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11388_ _11388_/A _11409_/Y vssd1 vssd1 vccd1 vccd1 _13628_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11885__D line[100] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[15\].VALID\[5\].FF_D A[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06979__D line[33] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[0\].CLKBUF\[3\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10339_ _10355_/CLK line[33] vssd1 vssd1 vccd1 vccd1 _10340_/A sky130_fd_sc_hd__dfxtp_1
X_13127_ _13155_/CLK line[42] vssd1 vssd1 vccd1 vccd1 _13128_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09355__D line[110] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13058_ _13058_/A _13089_/Y vssd1 vssd1 vccd1 vccd1 _13618_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[27\].CLKBUF\[0\] clk vssd1 vssd1 vccd1 vccd1 _10287_/CLK sky130_fd_sc_hd__clkbuf_4
XMUX.M\[3\].MUX\[1\] _13681_/Z _13751_/Z _13821_/Z _13891_/Z MUX.SEL0BUF\[3\]/X MUX.SEL1BUF\[3\]/X
+ vssd1 vssd1 vccd1 vccd1 Do[25] sky130_fd_sc_hd__mux4_1
X_12009_ _12035_/CLK line[43] vssd1 vssd1 vccd1 vccd1 _12010_/A sky130_fd_sc_hd__dfxtp_1
X_05880_ _05910_/CLK line[48] vssd1 vssd1 vccd1 vccd1 _05881_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07453__A _13910_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XDATA\[17\].CLKBUF\[6\] clk vssd1 vssd1 vccd1 vccd1 _07417_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_66_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07550_ _07550_/A _07559_/Y vssd1 vssd1 vccd1 vccd1 _13710_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07603__D line[77] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06501_ _06505_/CLK line[71] vssd1 vssd1 vccd1 vccd1 _06502_/A sky130_fd_sc_hd__dfxtp_1
X_07481_ _07485_/CLK line[7] vssd1 vssd1 vccd1 vccd1 _07482_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_22_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11125__D line[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09220_ _09220_/A _09239_/Y vssd1 vssd1 vccd1 vccd1 _13700_/Z sky130_fd_sc_hd__ebufn_2
X_06432_ _06432_/A _06439_/Y vssd1 vssd1 vccd1 vccd1 _13712_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06219__D line[70] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09151_ _09165_/CLK line[2] vssd1 vssd1 vccd1 vccd1 _09152_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_148_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06363_ _06365_/CLK line[8] vssd1 vssd1 vccd1 vccd1 _06364_/A sky130_fd_sc_hd__dfxtp_1
X_08102_ _08102_/A _08119_/Y vssd1 vssd1 vccd1 vccd1 _13702_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[7\].VALID\[11\].FF OVHB\[7\].V/CLK A[18] vssd1 vssd1 vccd1 vccd1 OVHB\[7\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_05314_ _05314_/A _05319_/Y vssd1 vssd1 vccd1 vccd1 _13714_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_30_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09082_ _09082_/A _09099_/Y vssd1 vssd1 vccd1 vccd1 _13842_/Z sky130_fd_sc_hd__ebufn_2
X_06294_ _06294_/A _06299_/Y vssd1 vssd1 vccd1 vccd1 _13854_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.M\[3\].MUX\[4\]_A3 _13867_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08033_ _08045_/CLK line[3] vssd1 vssd1 vccd1 vccd1 _08034_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_135_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05245_ _05245_/CLK line[9] vssd1 vssd1 vccd1 vccd1 _05246_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_190_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07628__A _13911_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05176_ _05176_/A _05179_/Y vssd1 vssd1 vccd1 vccd1 _13856_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11795__D line[64] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[5\].VALID\[10\].FF_D A[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09984_ _09984_/A _10009_/Y vssd1 vssd1 vccd1 vccd1 _13624_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05793__D line[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08935_ _08955_/CLK line[46] vssd1 vssd1 vccd1 vccd1 _08936_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10989__A _13925_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08866_ _08866_/A _08889_/Y vssd1 vssd1 vccd1 vccd1 _13626_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_17_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07817_ _07835_/CLK line[47] vssd1 vssd1 vccd1 vccd1 _07818_/A sky130_fd_sc_hd__dfxtp_1
X_08797_ _08815_/CLK line[111] vssd1 vssd1 vccd1 vccd1 _08798_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_44_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07748_ _07748_/A _07769_/Y vssd1 vssd1 vccd1 vccd1 _13628_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_199_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07679_ _07695_/CLK line[97] vssd1 vssd1 vccd1 vccd1 _07680_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[16\].CLKBUF\[3\] clk vssd1 vssd1 vccd1 vccd1 _07032_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__11035__D line[110] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09418_ _09418_/A _09449_/Y vssd1 vssd1 vccd1 vccd1 _13618_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_16_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06129__D line[43] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10690_ _10690_/A _10709_/Y vssd1 vssd1 vccd1 vccd1 _13770_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05033__D line[40] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10874__D line[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMUX.M\[2\].MUX\[3\] _13669_/Z _13739_/Z _13809_/Z _13879_/Z MUX.SEL0BUF\[2\]/X MUX.SEL1BUF\[2\]/X
+ vssd1 vssd1 vccd1 vccd1 Do[19] sky130_fd_sc_hd__mux4_1
X_09349_ _09375_/CLK line[107] vssd1 vssd1 vccd1 vccd1 _09350_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_185_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13250__D line[84] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05968__D line[83] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08344__D line[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12360_ _12360_/A _12389_/Y vssd1 vssd1 vccd1 vccd1 _13760_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_148_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XOVHB\[18\].VALID\[3\].FF OVHB\[18\].V/CLK A[10] vssd1 vssd1 vccd1 vccd1 OVHB\[18\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_11311_ _11335_/CLK line[108] vssd1 vssd1 vccd1 vccd1 _11312_/A sky130_fd_sc_hd__dfxtp_1
X_12291_ _12315_/CLK line[44] vssd1 vssd1 vccd1 vccd1 _12292_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[28\].VALID\[5\].FF_D A[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[3\].VALID\[8\].TOBUF OVHB\[3\].VALID\[8\].FF/Q OVHB\[3\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04931_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_107_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11242_ _11242_/A _11269_/Y vssd1 vssd1 vccd1 vccd1 _13762_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_180_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11173_ _11195_/CLK line[45] vssd1 vssd1 vccd1 vccd1 _11174_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_122_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10124_ _10124_/A _10149_/Y vssd1 vssd1 vccd1 vccd1 _13764_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_67_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_DATA\[25\].CLKBUF\[6\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10055_ _10075_/CLK line[46] vssd1 vssd1 vccd1 vccd1 _10056_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_57_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05208__D line[120] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13425__D line[36] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13814_ _13820_/CLK line[86] vssd1 vssd1 vccd1 vccd1 _13815_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08519__D line[97] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13745_ _13745_/A _13754_/Y vssd1 vssd1 vccd1 vccd1 _13745_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_204_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10957_ _10985_/CLK line[74] vssd1 vssd1 vccd1 vccd1 _10958_/A sky130_fd_sc_hd__dfxtp_1
X_13676_ _13680_/CLK line[23] vssd1 vssd1 vccd1 vccd1 _13677_/A sky130_fd_sc_hd__dfxtp_1
X_10888_ _10888_/A _10919_/Y vssd1 vssd1 vccd1 vccd1 _13688_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10784__D line[123] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12627_ _12627_/A _12634_/Y vssd1 vssd1 vccd1 vccd1 _13747_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_31_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13160__D line[48] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XDATA\[15\].CLKBUF\[0\] clk vssd1 vssd1 vccd1 vccd1 _06647_/CLK sky130_fd_sc_hd__clkbuf_4
XPHY_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12558_ _12560_/CLK line[24] vssd1 vssd1 vccd1 vccd1 _12559_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_8_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11509_ _11509_/A _11514_/Y vssd1 vssd1 vccd1 vccd1 _13749_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_144_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12354__A _13935_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12489_ _12489_/A _12494_/Y vssd1 vssd1 vccd1 vccd1 _13889_/Z sky130_fd_sc_hd__ebufn_2
X_05030_ _05030_/A _05039_/Y vssd1 vssd1 vccd1 vccd1 _13710_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12073__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09085__D line[100] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[16\].VALID\[5\].FF OVHB\[16\].V/CLK A[12] vssd1 vssd1 vccd1 vccd1 OVHB\[16\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_06981_ _06995_/CLK line[34] vssd1 vssd1 vccd1 vccd1 _06982_/A sky130_fd_sc_hd__dfxtp_1
XMUX.M\[1\].MUX\[5\] _13624_/Z _13694_/Z _13764_/Z _13834_/Z MUX.SEL0BUF\[1\]/X MUX.SEL1BUF\[1\]/X
+ vssd1 vssd1 vccd1 vccd1 Do[13] sky130_fd_sc_hd__mux4_1
XANTENNA__10024__D line[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08720_ _08720_/A _08749_/Y vssd1 vssd1 vccd1 vccd1 _13760_/Z sky130_fd_sc_hd__ebufn_2
X_05932_ _05932_/A _05949_/Y vssd1 vssd1 vccd1 vccd1 _13772_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05118__D line[93] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[10\].VALID\[3\].TOBUF OVHB\[10\].VALID\[3\].FF/Q OVHB\[10\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04919_/B2 sky130_fd_sc_hd__ebufn_2
X_08651_ _08675_/CLK line[44] vssd1 vssd1 vccd1 vccd1 _08652_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10959__D line[75] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05863_ _05875_/CLK line[35] vssd1 vssd1 vccd1 vccd1 _05864_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[9\].VALID\[0\].FF_D A[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13335__D line[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07602_ _07602_/A _07629_/Y vssd1 vssd1 vccd1 vccd1 _13762_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_93_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__04957__D line[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08582_ _08582_/A _08609_/Y vssd1 vssd1 vccd1 vccd1 _13622_/Z sky130_fd_sc_hd__ebufn_2
X_05794_ _05794_/A _05809_/Y vssd1 vssd1 vccd1 vccd1 _13634_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07333__D line[67] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07533_ _07555_/CLK line[45] vssd1 vssd1 vccd1 vccd1 _07534_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12529__A _13936_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07464_ _07464_/A _07489_/Y vssd1 vssd1 vccd1 vccd1 _13624_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12248__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09203_ _13916_/X wr vssd1 vssd1 vccd1 vccd1 _09203_/X sky130_fd_sc_hd__and2_1
X_06415_ _06435_/CLK line[46] vssd1 vssd1 vccd1 vccd1 _06416_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_148_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07395_ _07415_/CLK line[110] vssd1 vssd1 vccd1 vccd1 _07396_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_50_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09134_ _13915_/X vssd1 vssd1 vccd1 vccd1 _09134_/Y sky130_fd_sc_hd__inv_2
X_06346_ _06346_/A _06369_/Y vssd1 vssd1 vccd1 vccd1 _13626_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_147_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09065_ _09095_/CLK line[96] vssd1 vssd1 vccd1 vccd1 _09066_/A sky130_fd_sc_hd__dfxtp_1
X_06277_ _06295_/CLK line[111] vssd1 vssd1 vccd1 vccd1 _06278_/A sky130_fd_sc_hd__dfxtp_1
X_08016_ _08016_/A _08049_/Y vssd1 vssd1 vccd1 vccd1 _13616_/Z sky130_fd_sc_hd__ebufn_2
X_05228_ _05228_/A _05249_/Y vssd1 vssd1 vccd1 vccd1 _13628_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_104_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MUX.M\[2\].MUX\[5\]_A1 _13743_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12414__D line[86] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05159_ _05175_/CLK line[97] vssd1 vssd1 vccd1 vccd1 _05160_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_162_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07508__D line[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09967_ _09967_/A _09974_/Y vssd1 vssd1 vccd1 vccd1 _13887_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_103_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08918_ _08920_/CLK line[24] vssd1 vssd1 vccd1 vccd1 _08919_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09898_ _09900_/CLK line[88] vssd1 vssd1 vccd1 vccd1 _09899_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08189__A _13932_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09723__D line[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08849_ _08849_/A _08854_/Y vssd1 vssd1 vccd1 vccd1 _13889_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13823__A _13899_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11860_ _11860_/CLK line[89] vssd1 vssd1 vccd1 vccd1 _11861_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[14\].VALID\[7\].FF OVHB\[14\].V/CLK A[14] vssd1 vssd1 vccd1 vccd1 OVHB\[14\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_168_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10811_ _10811_/A _10814_/Y vssd1 vssd1 vccd1 vccd1 _13891_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_26_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11791_ _11791_/A _11794_/Y vssd1 vssd1 vccd1 vccd1 _13751_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_41_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13530_ _13540_/CLK line[84] vssd1 vssd1 vccd1 vccd1 _13531_/A sky130_fd_sc_hd__dfxtp_1
X_10742_ _10742_/CLK _10743_/X vssd1 vssd1 vccd1 vccd1 _10740_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA_MUX.M\[0\].MUX\[1\]_A2 _13770_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XMUX.M\[0\].MUX\[7\] _13642_/Z _13712_/Z _13782_/Z _13852_/Z MUX.SEL0BUF\[0\]/X MUX.SEL1BUF\[0\]/X
+ vssd1 vssd1 vccd1 vccd1 Do[7] sky130_fd_sc_hd__mux4_1
XOVHB\[4\].VALID\[13\].TOBUF OVHB\[4\].VALID\[13\].FF/Q OVHB\[4\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04916_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_185_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13461_ _13461_/A _13474_/Y vssd1 vssd1 vccd1 vccd1 _13741_/Z sky130_fd_sc_hd__ebufn_2
X_10673_ _13924_/X wr vssd1 vssd1 vccd1 vccd1 _10673_/X sky130_fd_sc_hd__and2_1
XANTENNA__05698__D line[88] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08074__D line[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12412_ _12420_/CLK line[85] vssd1 vssd1 vccd1 vccd1 _12413_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_138_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13392_ _13400_/CLK line[21] vssd1 vssd1 vccd1 vccd1 _13393_/A sky130_fd_sc_hd__dfxtp_1
X_12343_ _12343_/A _12354_/Y vssd1 vssd1 vccd1 vccd1 _13743_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[11\].VALID\[8\].FF_D A[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12274_ _12280_/CLK line[22] vssd1 vssd1 vccd1 vccd1 _12275_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_175_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11225_ _11225_/A _11234_/Y vssd1 vssd1 vccd1 vccd1 _13745_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_153_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12324__D line[59] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09483__A _13920_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11156_ _11160_/CLK line[23] vssd1 vssd1 vccd1 vccd1 _11157_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06322__D line[117] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10107_ _10107_/A _10114_/Y vssd1 vssd1 vccd1 vccd1 _13747_/Z sky130_fd_sc_hd__ebufn_2
X_11087_ _11087_/A _11094_/Y vssd1 vssd1 vccd1 vccd1 _13887_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_0_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09633__D line[109] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10038_ _10040_/CLK line[24] vssd1 vssd1 vccd1 vccd1 _10039_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13155__D line[41] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08249__D line[102] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11989_ _11989_/A _12004_/Y vssd1 vssd1 vccd1 vccd1 _13669_/Z sky130_fd_sc_hd__ebufn_2
X_13728_ _13750_/CLK line[61] vssd1 vssd1 vccd1 vccd1 _13729_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_31_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13659_ _13659_/A _13684_/Y vssd1 vssd1 vccd1 vccd1 _13659_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11403__D line[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06200_ _06200_/A _06229_/Y vssd1 vssd1 vccd1 vccd1 _13760_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[12\].VALID\[9\].FF OVHB\[12\].V/CLK A[16] vssd1 vssd1 vccd1 vccd1 OVHB\[12\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__09658__A _13920_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07180_ _07180_/A _07209_/Y vssd1 vssd1 vccd1 vccd1 _13620_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_157_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06131_ _06155_/CLK line[44] vssd1 vssd1 vccd1 vccd1 _06132_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09049__TE_B _09064_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09808__D line[61] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06062_ _06062_/A _06089_/Y vssd1 vssd1 vccd1 vccd1 _13622_/Z sky130_fd_sc_hd__ebufn_2
X_05013_ _05035_/CLK line[45] vssd1 vssd1 vccd1 vccd1 _05014_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_99_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13908__A A[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09821_ _09821_/A _09834_/Y vssd1 vssd1 vccd1 vccd1 _13741_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06232__D line[90] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09752_ _09760_/CLK line[21] vssd1 vssd1 vccd1 vccd1 _09753_/A sky130_fd_sc_hd__dfxtp_1
X_06964_ _13909_/Y vssd1 vssd1 vccd1 vccd1 _06964_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08703_ _08703_/A _08714_/Y vssd1 vssd1 vccd1 vccd1 _13743_/Z sky130_fd_sc_hd__ebufn_2
X_05915_ _05945_/CLK line[64] vssd1 vssd1 vccd1 vccd1 _05916_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10689__D line[65] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09683_ _09683_/A _09694_/Y vssd1 vssd1 vccd1 vccd1 _13883_/Z sky130_fd_sc_hd__ebufn_2
X_06895_ _06925_/CLK line[0] vssd1 vssd1 vccd1 vccd1 _06896_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13065__D line[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08634_ _08640_/CLK line[22] vssd1 vssd1 vccd1 vccd1 _08635_/A sky130_fd_sc_hd__dfxtp_1
X_05846_ _05846_/A _05879_/Y vssd1 vssd1 vccd1 vccd1 _13686_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08159__D line[75] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07063__D line[72] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[31\].VALID\[4\].FF_D A[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05777_ _05805_/CLK line[10] vssd1 vssd1 vccd1 vccd1 _05778_/A sky130_fd_sc_hd__dfxtp_1
X_08565_ _08565_/A _08574_/Y vssd1 vssd1 vccd1 vccd1 _13885_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07998__D line[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11163__A _13933_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07516_ _07520_/CLK line[23] vssd1 vssd1 vccd1 vccd1 _07517_/A sky130_fd_sc_hd__dfxtp_1
X_08496_ _08500_/CLK line[87] vssd1 vssd1 vccd1 vccd1 _08497_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07447_ _07447_/A _07454_/Y vssd1 vssd1 vccd1 vccd1 _13887_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11313__D line[109] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[30\].VALID\[14\].FF_D A[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06407__D line[42] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[24\].VALID\[8\].FF_D A[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07378_ _07380_/CLK line[88] vssd1 vssd1 vccd1 vccd1 _07379_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_195_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05311__D line[39] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09117_ _09117_/A _09134_/Y vssd1 vssd1 vccd1 vccd1 _13877_/Z sky130_fd_sc_hd__ebufn_2
X_06329_ _06329_/A _06334_/Y vssd1 vssd1 vccd1 vccd1 _13889_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_89_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09048_ _09060_/CLK line[83] vssd1 vssd1 vccd1 vccd1 _09049_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_163_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08622__D line[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07238__D line[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11010_ _11020_/CLK line[84] vssd1 vssd1 vccd1 vccd1 _11011_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_145_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11338__A _13933_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12961_ _12961_/A _12984_/Y vssd1 vssd1 vccd1 vccd1 _13801_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_73_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_OVHB\[12\].VALID\[12\].FF_D A[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11912_ _11930_/CLK line[127] vssd1 vssd1 vccd1 vccd1 _11913_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_45_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12892_ _12910_/CLK line[63] vssd1 vssd1 vccd1 vccd1 _12893_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_205_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XDATA\[7\].CLKBUF\[7\] clk vssd1 vssd1 vccd1 vccd1 _13332_/CLK sky130_fd_sc_hd__clkbuf_4
XOVHB\[17\].VALID\[3\].TOBUF OVHB\[17\].VALID\[3\].FF/Q OVHB\[17\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04919_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_54_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11843_ _11843_/A _11864_/Y vssd1 vssd1 vccd1 vccd1 _13803_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[7\].VALID\[0\].FF OVHB\[7\].V/CLK A[7] vssd1 vssd1 vccd1 vccd1 OVHB\[7\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13703__D line[35] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XOVHB\[20\].VALID\[14\].TOBUF OVHB\[20\].VALID\[14\].FF/Q OVHB\[20\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[18\].CLKBUF\[0\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11774_ _11790_/CLK line[49] vssd1 vssd1 vccd1 vccd1 _11775_/A sky130_fd_sc_hd__dfxtp_1
X_13513_ _13513_/A _13544_/Y vssd1 vssd1 vccd1 vccd1 _13793_/Z sky130_fd_sc_hd__ebufn_2
X_10725_ _10725_/A _10744_/Y vssd1 vssd1 vccd1 vccd1 _13805_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_201_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13444_ _13470_/CLK line[59] vssd1 vssd1 vccd1 vccd1 _13445_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05221__D line[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10656_ _10670_/CLK line[50] vssd1 vssd1 vccd1 vccd1 _10657_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_173_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_OVHB\[22\].VALID\[11\].FF_D A[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10587_ _10587_/A _10604_/Y vssd1 vssd1 vccd1 vccd1 _13667_/Z sky130_fd_sc_hd__ebufn_2
X_13375_ _13375_/A _13404_/Y vssd1 vssd1 vccd1 vccd1 _13655_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_126_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12326_ _12350_/CLK line[60] vssd1 vssd1 vccd1 vccd1 _12327_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_126_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12054__D line[49] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12257_ _12257_/A _12284_/Y vssd1 vssd1 vccd1 vccd1 _13657_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_142_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XOVHB\[26\].V OVHB\[26\].V/CLK TIE/HI rst_n vssd1 vssd1 vccd1 vccd1 OVHB\[26\].V/Q
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07148__D line[125] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11208_ _11230_/CLK line[61] vssd1 vssd1 vccd1 vccd1 _11209_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_141_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12188_ _12210_/CLK line[125] vssd1 vssd1 vccd1 vccd1 _12189_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12989__D line[107] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11893__D line[104] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[5\].VALID\[3\].FF_D A[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11139_ _11139_/A _11164_/Y vssd1 vssd1 vccd1 vccd1 _13659_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06987__D line[37] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09363__D line[99] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05700_ _05700_/CLK line[89] vssd1 vssd1 vccd1 vccd1 _05701_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10302__D line[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06680_ _06680_/CLK line[25] vssd1 vssd1 vccd1 vccd1 _06681_/A sky130_fd_sc_hd__dfxtp_1
X_05631_ _05631_/A _05634_/Y vssd1 vssd1 vccd1 vccd1 _13751_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_91_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08350_ _08360_/CLK line[20] vssd1 vssd1 vccd1 vccd1 _08351_/A sky130_fd_sc_hd__dfxtp_1
X_05562_ _05562_/CLK _05563_/X vssd1 vssd1 vccd1 vccd1 _05560_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_211_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07611__D line[66] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07301_ _07301_/A _07314_/Y vssd1 vssd1 vccd1 vccd1 _13741_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12229__D line[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDATA\[6\].CLKBUF\[4\] clk vssd1 vssd1 vccd1 vccd1 _12947_/CLK sky130_fd_sc_hd__clkbuf_4
X_08281_ _08281_/A _08294_/Y vssd1 vssd1 vccd1 vccd1 _13881_/Z sky130_fd_sc_hd__ebufn_2
X_05493_ _13900_/X wr vssd1 vssd1 vccd1 vccd1 _05493_/X sky130_fd_sc_hd__and2_1
XFILLER_177_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07232_ _07240_/CLK line[21] vssd1 vssd1 vccd1 vccd1 _07233_/A sky130_fd_sc_hd__dfxtp_1
X_07163_ _07163_/A _07174_/Y vssd1 vssd1 vccd1 vccd1 _13883_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[5\].VALID\[2\].FF OVHB\[5\].V/CLK A[9] vssd1 vssd1 vccd1 vccd1 OVHB\[5\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XOVHB\[23\].VALID\[2\].TOBUF OVHB\[23\].VALID\[2\].FF/Q OVHB\[23\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04930_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__09538__D line[51] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06114_ _06120_/CLK line[22] vssd1 vssd1 vccd1 vccd1 _06115_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__04970__D line[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07094_ _07100_/CLK line[86] vssd1 vssd1 vccd1 vccd1 _07095_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_132_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06045_ _06045_/A _06054_/Y vssd1 vssd1 vccd1 vccd1 _13885_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[20\].CGAND_B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XOVHB\[17\].V OVHB\[17\].V/CLK TIE/HI rst_n vssd1 vssd1 vccd1 vccd1 OVHB\[17\].V/Q
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_87_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[5\].CGAND_B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09804_ _09830_/CLK line[59] vssd1 vssd1 vccd1 vccd1 _09805_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[24\].CGAND_A _13920_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06897__D line[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__04919__B2 _04919_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07996_ _08010_/CLK line[114] vssd1 vssd1 vccd1 vccd1 _07997_/A sky130_fd_sc_hd__dfxtp_1
X_09735_ _09735_/A _09764_/Y vssd1 vssd1 vccd1 vccd1 _13655_/Z sky130_fd_sc_hd__ebufn_2
X_06947_ _06947_/A _06964_/Y vssd1 vssd1 vccd1 vccd1 _13667_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_101_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[9\].CGAND_A _13899_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09666_ _09690_/CLK line[124] vssd1 vssd1 vccd1 vccd1 _09667_/A sky130_fd_sc_hd__dfxtp_1
X_06878_ _06890_/CLK line[115] vssd1 vssd1 vccd1 vccd1 _06879_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_43_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08617_ _08617_/A _08644_/Y vssd1 vssd1 vccd1 vccd1 _13657_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05829_ _05829_/A _05844_/Y vssd1 vssd1 vccd1 vccd1 _13669_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09597_ _09597_/A _09624_/Y vssd1 vssd1 vccd1 vccd1 _13797_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_42_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08548_ _08570_/CLK line[125] vssd1 vssd1 vccd1 vccd1 _08549_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08479_ _08479_/A _08504_/Y vssd1 vssd1 vccd1 vccd1 _13799_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_168_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11043__D line[99] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06137__D line[47] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10510_ _10530_/CLK line[126] vssd1 vssd1 vccd1 vccd1 _10511_/A sky130_fd_sc_hd__dfxtp_1
X_11490_ _11510_/CLK line[62] vssd1 vssd1 vccd1 vccd1 _11491_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11978__D line[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10441_ _10441_/A _10464_/Y vssd1 vssd1 vccd1 vccd1 _13801_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_108_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XDATA\[5\].CLKBUF\[1\] clk vssd1 vssd1 vccd1 vccd1 _12562_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__05976__D line[87] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08352__D line[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10372_ _10390_/CLK line[63] vssd1 vssd1 vccd1 vccd1 _10373_/A sky130_fd_sc_hd__dfxtp_1
X_13160_ _13190_/CLK line[48] vssd1 vssd1 vccd1 vccd1 _13161_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_200_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12111_ _12111_/A _12144_/Y vssd1 vssd1 vccd1 vccd1 _13791_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[15\].VALID\[8\].TOBUF OVHB\[15\].VALID\[8\].FF/Q OVHB\[15\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04931_/B2 sky130_fd_sc_hd__ebufn_2
X_13091_ _13091_/A _13124_/Y vssd1 vssd1 vccd1 vccd1 _13651_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_156_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12042_ _12070_/CLK line[58] vssd1 vssd1 vccd1 vccd1 _12043_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[3\].VALID\[4\].FF OVHB\[3\].V/CLK A[11] vssd1 vssd1 vccd1 vccd1 OVHB\[3\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_78_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12602__D line[58] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06600__D line[116] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11218__D line[51] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12944_ _12944_/A _12949_/Y vssd1 vssd1 vccd1 vccd1 _13784_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_46_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09911__D line[108] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12875_ _12875_/CLK line[41] vssd1 vssd1 vccd1 vccd1 _12876_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13433__D line[40] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11826_ _11826_/A _11829_/Y vssd1 vssd1 vccd1 vccd1 _13786_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08527__D line[101] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDATA\[25\].CLKBUF\[5\] clk vssd1 vssd1 vccd1 vccd1 _09902_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_202_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11757_ _11757_/CLK _11758_/X vssd1 vssd1 vccd1 vccd1 _11755_/CLK sky130_fd_sc_hd__dlclkp_1
XPHY_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10708_ _13924_/X wr vssd1 vssd1 vccd1 vccd1 _10708_/X sky130_fd_sc_hd__and2_1
XPHY_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11688_ _13927_/X wr vssd1 vssd1 vccd1 vccd1 _11688_/X sky130_fd_sc_hd__and2_1
XANTENNA__10792__D line[127] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13427_ _13435_/CLK line[37] vssd1 vssd1 vccd1 vccd1 _13428_/A sky130_fd_sc_hd__dfxtp_1
X_10639_ _13924_/X vssd1 vssd1 vccd1 vccd1 _10639_/Y sky130_fd_sc_hd__inv_2
XANTENNA__05886__D line[60] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[16\].CLKBUF\[2\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08262__D line[122] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13358_ _13358_/A _13369_/Y vssd1 vssd1 vccd1 vccd1 _13638_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_115_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12309_ _12315_/CLK line[38] vssd1 vssd1 vccd1 vccd1 _12310_/A sky130_fd_sc_hd__dfxtp_1
X_13289_ _13295_/CLK line[102] vssd1 vssd1 vccd1 vccd1 _13290_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13608__D line[120] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07850_ _07870_/CLK line[62] vssd1 vssd1 vccd1 vccd1 _07851_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09093__D line[104] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06510__D line[80] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06801_ _06801_/A _06824_/Y vssd1 vssd1 vccd1 vccd1 _13801_/Z sky130_fd_sc_hd__ebufn_2
X_04993_ _04993_/A _05004_/Y vssd1 vssd1 vccd1 vccd1 _13673_/Z sky130_fd_sc_hd__ebufn_2
X_07781_ _07781_/A _07804_/Y vssd1 vssd1 vccd1 vccd1 _13661_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10032__D line[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13193__A _13938_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09520_ _09550_/CLK line[48] vssd1 vssd1 vccd1 vccd1 _09521_/A sky130_fd_sc_hd__dfxtp_1
X_06732_ _06750_/CLK line[63] vssd1 vssd1 vccd1 vccd1 _06733_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[21\].VALID\[7\].TOBUF OVHB\[21\].VALID\[7\].FF/Q OVHB\[21\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/A2 sky130_fd_sc_hd__ebufn_2
XANTENNA__05126__D line[82] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[9\].CLKBUF\[2\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05704__A _13901_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[1\].VALID\[6\].FF OVHB\[1\].V/CLK A[13] vssd1 vssd1 vccd1 vccd1 OVHB\[1\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_09451_ _09451_/A _09484_/Y vssd1 vssd1 vccd1 vccd1 _13651_/Z sky130_fd_sc_hd__ebufn_2
X_06663_ _06663_/A _06684_/Y vssd1 vssd1 vccd1 vccd1 _13663_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10967__D line[79] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13343__D line[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[19\].VALID\[12\].FF_D A[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08402_ _08430_/CLK line[58] vssd1 vssd1 vccd1 vccd1 _08403_/A sky130_fd_sc_hd__dfxtp_1
X_05614_ _05630_/CLK line[49] vssd1 vssd1 vccd1 vccd1 _05615_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__04965__D line[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08437__D line[74] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05423__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09382_ _09410_/CLK line[122] vssd1 vssd1 vccd1 vccd1 _09383_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_52_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06594_ _06610_/CLK line[113] vssd1 vssd1 vccd1 vccd1 _06595_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07341__D line[71] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08333_ _08333_/A _08364_/Y vssd1 vssd1 vccd1 vccd1 _13653_/Z sky130_fd_sc_hd__ebufn_2
X_05545_ _05545_/A _05564_/Y vssd1 vssd1 vccd1 vccd1 _13665_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_32_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08264_ _08290_/CLK line[123] vssd1 vssd1 vccd1 vccd1 _08265_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_20_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MUX.M\[3\].MUX\[7\]_A1 _13733_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05476_ _05490_/CLK line[114] vssd1 vssd1 vccd1 vccd1 _05477_/A sky130_fd_sc_hd__dfxtp_1
X_07215_ _07215_/A _07244_/Y vssd1 vssd1 vccd1 vccd1 _13655_/Z sky130_fd_sc_hd__ebufn_2
X_08195_ _08195_/A _08224_/Y vssd1 vssd1 vccd1 vccd1 _13795_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[24\].CLKBUF\[2\] clk vssd1 vssd1 vccd1 vccd1 _09517_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__09268__D line[56] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07146_ _07170_/CLK line[124] vssd1 vssd1 vccd1 vccd1 _07147_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_106_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_OVHB\[29\].VALID\[11\].FF_D A[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13368__A _13898_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07077_ _07077_/A _07104_/Y vssd1 vssd1 vccd1 vccd1 _13797_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10207__D line[101] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06028_ _06050_/CLK line[125] vssd1 vssd1 vccd1 vccd1 _06029_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08900__D line[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13518__D line[93] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07516__D line[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07979_ _13912_/X vssd1 vssd1 vccd1 vccd1 _07979_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MUX.M\[1\].MUX\[3\]_A2 _13760_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09718_ _09718_/A _09729_/Y vssd1 vssd1 vccd1 vccd1 _13638_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_28_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10990_ _11020_/CLK line[80] vssd1 vssd1 vccd1 vccd1 _10991_/A sky130_fd_sc_hd__dfxtp_1
X_09649_ _09655_/CLK line[102] vssd1 vssd1 vccd1 vccd1 _09650_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_55_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12660_ _12660_/A _12669_/Y vssd1 vssd1 vccd1 vccd1 _13780_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07251__D line[44] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11611_ _11615_/CLK line[103] vssd1 vssd1 vccd1 vccd1 _11612_/A sky130_fd_sc_hd__dfxtp_1
XPHY_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12591_ _12595_/CLK line[39] vssd1 vssd1 vccd1 vccd1 _12592_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11542_ _11542_/A _11549_/Y vssd1 vssd1 vccd1 vccd1 _13782_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[17\].VALID\[13\].TOBUF OVHB\[17\].VALID\[13\].FF/Q OVHB\[17\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04916_/B2 sky130_fd_sc_hd__ebufn_2
XPHY_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11473_ _11475_/CLK line[40] vssd1 vssd1 vccd1 vccd1 _11474_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09178__D line[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13212_ _13212_/A _13229_/Y vssd1 vssd1 vccd1 vccd1 _13772_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_109_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10424_ _10424_/A _10429_/Y vssd1 vssd1 vccd1 vccd1 _13784_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_152_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10117__D line[74] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13143_ _13155_/CLK line[35] vssd1 vssd1 vccd1 vccd1 _13144_/A sky130_fd_sc_hd__dfxtp_1
X_10355_ _10355_/CLK line[41] vssd1 vssd1 vccd1 vccd1 _10356_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_3_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_OVHB\[1\].VALID\[6\].FF_D A[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13074_ _13074_/A _13089_/Y vssd1 vssd1 vccd1 vccd1 _13634_/Z sky130_fd_sc_hd__ebufn_2
X_10286_ _10286_/A _10289_/Y vssd1 vssd1 vccd1 vccd1 _13646_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_2_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12332__D line[63] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12025_ _12035_/CLK line[36] vssd1 vssd1 vccd1 vccd1 _12026_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_111_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XDATA\[13\].CLKBUF\[5\] clk vssd1 vssd1 vccd1 vccd1 _06262_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__07426__D line[124] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[28\].VALID\[1\].FF OVHB\[28\].V/CLK A[8] vssd1 vssd1 vccd1 vccd1 OVHB\[28\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06330__D line[121] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13976_ _13982_/C _13982_/B _13982_/A _13982_/D vssd1 vssd1 vccd1 vccd1 _13976_/X
+ sky130_fd_sc_hd__and4bb_4
XFILLER_202_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09641__D line[98] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12927_ _12945_/CLK line[79] vssd1 vssd1 vccd1 vccd1 _12928_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_46_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[10\].VALID\[12\].TOBUF OVHB\[10\].VALID\[12\].FF/Q OVHB\[10\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04929_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_34_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12858_ _12858_/A _12879_/Y vssd1 vssd1 vccd1 vccd1 _13698_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_61_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11809_ _11825_/CLK line[65] vssd1 vssd1 vccd1 vccd1 _11810_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12789_ _12805_/CLK line[1] vssd1 vssd1 vccd1 vccd1 _12790_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_30_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05330_ _05350_/CLK line[62] vssd1 vssd1 vccd1 vccd1 _05331_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_147_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05261_ _05261_/A _05284_/Y vssd1 vssd1 vccd1 vccd1 _13661_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12507__D line[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07000_ _07030_/CLK line[48] vssd1 vssd1 vccd1 vccd1 _07001_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_174_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06505__D line[73] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05192_ _05210_/CLK line[127] vssd1 vssd1 vccd1 vccd1 _05193_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09816__D line[50] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08951_ _08955_/CLK line[39] vssd1 vssd1 vccd1 vccd1 _08952_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[14\].CLKBUF\[4\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07902_ _07902_/A _07909_/Y vssd1 vssd1 vccd1 vccd1 _13782_/Z sky130_fd_sc_hd__ebufn_2
X_08882_ _08882_/A _08889_/Y vssd1 vssd1 vccd1 vccd1 _13642_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_111_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06240__D line[94] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07833_ _07835_/CLK line[40] vssd1 vssd1 vccd1 vccd1 _07834_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_96_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07764_ _07764_/A _07769_/Y vssd1 vssd1 vccd1 vccd1 _13644_/Z sky130_fd_sc_hd__ebufn_2
X_04976_ _05000_/CLK line[28] vssd1 vssd1 vccd1 vccd1 _04977_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_112_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[16\].VALID\[3\].FF_D A[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDATA\[12\].CLKBUF\[2\] clk vssd1 vssd1 vccd1 vccd1 _05877_/CLK sky130_fd_sc_hd__clkbuf_4
X_09503_ _09515_/CLK line[35] vssd1 vssd1 vccd1 vccd1 _09504_/A sky130_fd_sc_hd__dfxtp_1
X_06715_ _06715_/CLK line[41] vssd1 vssd1 vccd1 vccd1 _06716_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10697__D line[69] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13073__D line[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07695_ _07695_/CLK line[105] vssd1 vssd1 vccd1 vccd1 _07696_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_24_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09434_ _09434_/A _09449_/Y vssd1 vssd1 vccd1 vccd1 _13634_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08167__D line[79] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06646_ _06646_/A _06649_/Y vssd1 vssd1 vccd1 vccd1 _13646_/Z sky130_fd_sc_hd__ebufn_2
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XOVHB\[26\].VALID\[3\].FF OVHB\[26\].V/CLK A[10] vssd1 vssd1 vccd1 vccd1 OVHB\[26\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_188_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09365_ _09375_/CLK line[100] vssd1 vssd1 vccd1 vccd1 _09366_/A sky130_fd_sc_hd__dfxtp_1
X_06577_ _06577_/CLK _06578_/X vssd1 vssd1 vccd1 vccd1 _06575_/CLK sky130_fd_sc_hd__dlclkp_1
X_08316_ _08316_/A _08329_/Y vssd1 vssd1 vccd1 vccd1 _13636_/Z sky130_fd_sc_hd__ebufn_2
X_05528_ _13901_/X wr vssd1 vssd1 vccd1 vccd1 _05528_/X sky130_fd_sc_hd__and2_1
XANTENNA_DATA\[7\].CLKBUF\[4\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09296_ _09296_/A _09309_/Y vssd1 vssd1 vccd1 vccd1 _13776_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_20_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05459_ _13900_/X vssd1 vssd1 vccd1 vccd1 _05459_/Y sky130_fd_sc_hd__inv_2
X_08247_ _08255_/CLK line[101] vssd1 vssd1 vccd1 vccd1 _08248_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11321__D line[98] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06415__D line[46] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08178_ _08178_/A _08189_/Y vssd1 vssd1 vccd1 vccd1 _13778_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_192_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07129_ _07135_/CLK line[102] vssd1 vssd1 vccd1 vccd1 _07130_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_97_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[10\].CG_CLK clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10140_ _10140_/A _10149_/Y vssd1 vssd1 vccd1 vccd1 _13780_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08630__D line[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13248__D line[83] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[30\].VALID\[12\].TOBUF OVHB\[30\].VALID\[12\].FF/Q OVHB\[30\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04929_/B2 sky130_fd_sc_hd__ebufn_2
X_10071_ _10075_/CLK line[39] vssd1 vssd1 vccd1 vccd1 _10072_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_87_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13830_ _13830_/A _13859_/Y vssd1 vssd1 vccd1 vccd1 _13830_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_46_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XOVHB\[3\].VALID\[4\].TOBUF OVHB\[3\].VALID\[4\].FF/Q OVHB\[3\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04925_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_56_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13761_ _13785_/CLK line[76] vssd1 vssd1 vccd1 vccd1 _13762_/A sky130_fd_sc_hd__dfxtp_1
X_10973_ _10985_/CLK line[67] vssd1 vssd1 vccd1 vccd1 _10974_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_204_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MUX.M\[0\].MUX\[4\]_A0 _13636_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12712_ _12712_/A _12739_/Y vssd1 vssd1 vccd1 vccd1 _13832_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_16_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XOVHB\[28\].VALID\[7\].TOBUF OVHB\[28\].VALID\[7\].FF/Q OVHB\[28\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/A2 sky130_fd_sc_hd__ebufn_2
X_13692_ _13692_/A _13719_/Y vssd1 vssd1 vccd1 vccd1 _13692_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_204_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12643_ _12665_/CLK line[77] vssd1 vssd1 vccd1 vccd1 _12644_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_102_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13711__D line[39] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08805__D line[100] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12574_ _12574_/A _12599_/Y vssd1 vssd1 vccd1 vccd1 _13694_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_196_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[29\].VOBUF OVHB\[29\].V/Q OVHB\[29\].INV/Y vssd1 vssd1 vccd1 vccd1 _04912_/B1
+ sky130_fd_sc_hd__ebufn_2
XPHY_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11525_ _11545_/CLK line[78] vssd1 vssd1 vccd1 vccd1 _11526_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_184_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XOVHB\[24\].VALID\[5\].FF OVHB\[24\].V/CLK A[12] vssd1 vssd1 vccd1 vccd1 OVHB\[24\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_11456_ _11456_/A _11479_/Y vssd1 vssd1 vccd1 vccd1 _13696_/Z sky130_fd_sc_hd__ebufn_2
X_10407_ _10425_/CLK line[79] vssd1 vssd1 vccd1 vccd1 _10408_/A sky130_fd_sc_hd__dfxtp_1
X_11387_ _11405_/CLK line[15] vssd1 vssd1 vccd1 vccd1 _11388_/A sky130_fd_sc_hd__dfxtp_1
X_13126_ _13126_/A _13159_/Y vssd1 vssd1 vccd1 vccd1 _13686_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_124_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08540__D line[112] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10338_ _10338_/A _10359_/Y vssd1 vssd1 vccd1 vccd1 _13698_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_97_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12062__D line[53] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13057_ _13085_/CLK line[10] vssd1 vssd1 vccd1 vccd1 _13058_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_140_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10269_ _10285_/CLK line[1] vssd1 vssd1 vccd1 vccd1 _10270_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07156__D line[114] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12008_ _12008_/A _12039_/Y vssd1 vssd1 vccd1 vccd1 _13688_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07734__A _13911_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12997__D line[111] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[29\].VALID\[3\].FF_D A[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06995__D line[41] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07453__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09371__D line[103] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13959_ _13960_/A _13960_/B _13960_/C _13960_/D vssd1 vssd1 vccd1 vccd1 _13959_/X
+ sky130_fd_sc_hd__and4b_4
XANTENNA__10310__D line[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06500_ _06500_/A _06509_/Y vssd1 vssd1 vccd1 vccd1 _13780_/Z sky130_fd_sc_hd__ebufn_2
X_07480_ _07480_/A _07489_/Y vssd1 vssd1 vccd1 vccd1 _13640_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_62_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05404__D line[81] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06431_ _06435_/CLK line[39] vssd1 vssd1 vccd1 vccd1 _06432_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_21_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13621__D line[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06362_ _06362_/A _06369_/Y vssd1 vssd1 vccd1 vccd1 _13642_/Z sky130_fd_sc_hd__ebufn_2
X_09150_ _09150_/A _09169_/Y vssd1 vssd1 vccd1 vccd1 _13630_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08715__D line[64] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05313_ _05315_/CLK line[40] vssd1 vssd1 vccd1 vccd1 _05314_/A sky130_fd_sc_hd__dfxtp_1
X_08101_ _08115_/CLK line[34] vssd1 vssd1 vccd1 vccd1 _08102_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12237__D line[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09081_ _09095_/CLK line[98] vssd1 vssd1 vccd1 vccd1 _09082_/A sky130_fd_sc_hd__dfxtp_1
X_06293_ _06295_/CLK line[104] vssd1 vssd1 vccd1 vccd1 _06294_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_174_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08032_ _08032_/A _08049_/Y vssd1 vssd1 vccd1 vccd1 _13632_/Z sky130_fd_sc_hd__ebufn_2
X_05244_ _05244_/A _05249_/Y vssd1 vssd1 vccd1 vccd1 _13644_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07909__A _13912_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05175_ _05175_/CLK line[105] vssd1 vssd1 vccd1 vccd1 _05176_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07628__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09546__D line[55] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09983_ _10005_/CLK line[13] vssd1 vssd1 vccd1 vccd1 _09984_/A sky130_fd_sc_hd__dfxtp_1
X_08934_ _08934_/A _08959_/Y vssd1 vssd1 vccd1 vccd1 _13694_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[22\].VALID\[7\].FF OVHB\[22\].V/CLK A[14] vssd1 vssd1 vccd1 vccd1 OVHB\[22\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_130_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08865_ _08885_/CLK line[14] vssd1 vssd1 vccd1 vccd1 _08866_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[30\].VALID\[12\].FF OVHB\[30\].V/CLK A[19] vssd1 vssd1 vccd1 vccd1 OVHB\[30\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_111_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12700__D line[89] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07816_ _07816_/A _07839_/Y vssd1 vssd1 vccd1 vccd1 _13696_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_123_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09281__D line[76] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08796_ _08796_/A _08819_/Y vssd1 vssd1 vccd1 vccd1 _13836_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_38_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07747_ _07765_/CLK line[15] vssd1 vssd1 vccd1 vccd1 _07748_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_84_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_DATA\[12\].CLKBUF\[6\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_04959_ _04965_/CLK line[6] vssd1 vssd1 vccd1 vccd1 _04960_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10220__D line[112] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07678_ _07678_/A _07699_/Y vssd1 vssd1 vccd1 vccd1 _13838_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_16_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09417_ _09445_/CLK line[10] vssd1 vssd1 vccd1 vccd1 _09418_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DECH.DEC0.AND1_A_N A_h[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06629_ _06645_/CLK line[1] vssd1 vssd1 vccd1 vccd1 _06630_/A sky130_fd_sc_hd__dfxtp_1
X_09348_ _09348_/A _09379_/Y vssd1 vssd1 vccd1 vccd1 _13828_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[30\].VOBUF OVHB\[30\].V/Q OVHB\[30\].INV/Y vssd1 vssd1 vccd1 vccd1 _04912_/B1
+ sky130_fd_sc_hd__ebufn_2
XANTENNA__12147__D line[106] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09279_ _09305_/CLK line[75] vssd1 vssd1 vccd1 vccd1 _09280_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11051__D line[103] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11310_ _11310_/A _11339_/Y vssd1 vssd1 vccd1 vccd1 _13830_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_32_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06145__D line[36] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12290_ _12290_/A _12319_/Y vssd1 vssd1 vccd1 vccd1 _13690_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_113_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11986__D line[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11241_ _11265_/CLK line[76] vssd1 vssd1 vccd1 vccd1 _11242_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[20\].VALID\[14\].FF OVHB\[20\].V/CLK A[21] vssd1 vssd1 vccd1 vccd1 OVHB\[20\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XOVHB\[1\].VALID\[9\].TOBUF OVHB\[1\].VALID\[9\].FF/Q OVHB\[1\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04914_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[5\].CLKBUF\[6\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09456__D line[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08360__D line[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11172_ _11172_/A _11199_/Y vssd1 vssd1 vccd1 vccd1 _13692_/Z sky130_fd_sc_hd__ebufn_2
X_10123_ _10145_/CLK line[77] vssd1 vssd1 vccd1 vccd1 _10124_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_164_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10054_ _10054_/A _10079_/Y vssd1 vssd1 vccd1 vccd1 _13694_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12610__D line[62] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07704__D line[123] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05074__A _13931_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__04915__A2_N _04915_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13813_ _13813_/A _13824_/Y vssd1 vssd1 vccd1 vccd1 _13813_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11226__D line[55] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XOVHB\[20\].VALID\[9\].FF OVHB\[20\].V/CLK A[16] vssd1 vssd1 vccd1 vccd1 OVHB\[20\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_113_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13744_ _13750_/CLK line[54] vssd1 vssd1 vccd1 vccd1 _13745_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_73_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10956_ _10956_/A _10989_/Y vssd1 vssd1 vccd1 vccd1 _13756_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_188_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13675_ _13675_/A _13684_/Y vssd1 vssd1 vccd1 vccd1 _13675_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_43_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10887_ _10915_/CLK line[42] vssd1 vssd1 vccd1 vccd1 _10888_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_31_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12626_ _12630_/CLK line[55] vssd1 vssd1 vccd1 vccd1 _12627_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08535__D line[105] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12557_ _12557_/A _12564_/Y vssd1 vssd1 vccd1 vccd1 _13677_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06055__D line[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11508_ _11510_/CLK line[56] vssd1 vssd1 vccd1 vccd1 _11509_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_172_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12488_ _12490_/CLK line[120] vssd1 vssd1 vccd1 vccd1 _12489_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_172_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11439_ _11439_/A _11444_/Y vssd1 vssd1 vccd1 vccd1 _13679_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05894__D line[49] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05249__A _13900_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08270__D line[126] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13109_ _13109_/A _13124_/Y vssd1 vssd1 vccd1 vccd1 _13669_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_86_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06980_ _06980_/A _06999_/Y vssd1 vssd1 vccd1 vccd1 _13700_/Z sky130_fd_sc_hd__ebufn_2
X_05931_ _05945_/CLK line[66] vssd1 vssd1 vccd1 vccd1 _05932_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[12\].VALID\[6\].FF_D A[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08650_ _08650_/A _08679_/Y vssd1 vssd1 vccd1 vccd1 _13690_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_39_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05862_ _05862_/A _05879_/Y vssd1 vssd1 vccd1 vccd1 _13702_/Z sky130_fd_sc_hd__ebufn_2
X_07601_ _07625_/CLK line[76] vssd1 vssd1 vccd1 vccd1 _07602_/A sky130_fd_sc_hd__dfxtp_1
X_08581_ _08605_/CLK line[12] vssd1 vssd1 vccd1 vccd1 _08582_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11136__D line[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05793_ _05805_/CLK line[3] vssd1 vssd1 vccd1 vccd1 _05794_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_54_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10040__D line[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07532_ _07532_/A _07559_/Y vssd1 vssd1 vccd1 vccd1 _13692_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05134__D line[86] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10975__D line[68] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07463_ _07485_/CLK line[13] vssd1 vssd1 vccd1 vccd1 _07464_/A sky130_fd_sc_hd__dfxtp_1
XMUX.SEL0BUF\[0\] A[0] vssd1 vssd1 vccd1 vccd1 MUX.SEL0BUF\[0\]/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__13351__D line[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09202_ _09202_/CLK _09203_/X vssd1 vssd1 vccd1 vccd1 _09200_/CLK sky130_fd_sc_hd__dlclkp_1
X_06414_ _06414_/A _06439_/Y vssd1 vssd1 vccd1 vccd1 _13694_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_50_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08445__D line[78] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07394_ _07394_/A _07419_/Y vssd1 vssd1 vccd1 vccd1 _13834_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_210_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09133_ _13915_/X wr vssd1 vssd1 vccd1 vccd1 _09133_/X sky130_fd_sc_hd__and2_1
X_06345_ _06365_/CLK line[14] vssd1 vssd1 vccd1 vccd1 _06346_/A sky130_fd_sc_hd__dfxtp_1
X_09064_ _13915_/X vssd1 vssd1 vccd1 vccd1 _09064_/Y sky130_fd_sc_hd__inv_2
X_06276_ _06276_/A _06299_/Y vssd1 vssd1 vccd1 vccd1 _13836_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06543__A _13904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08015_ _08045_/CLK line[0] vssd1 vssd1 vccd1 vccd1 _08016_/A sky130_fd_sc_hd__dfxtp_1
X_05227_ _05245_/CLK line[15] vssd1 vssd1 vccd1 vccd1 _05228_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_190_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MUX.M\[2\].MUX\[5\]_A2 _13813_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05158_ _05158_/A _05179_/Y vssd1 vssd1 vccd1 vccd1 _13838_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_89_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10215__D line[105] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09966_ _09970_/CLK line[119] vssd1 vssd1 vccd1 vccd1 _09967_/A sky130_fd_sc_hd__dfxtp_1
X_05089_ _05105_/CLK line[65] vssd1 vssd1 vccd1 vccd1 _05090_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05309__D line[38] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08917_ _08917_/A _08924_/Y vssd1 vssd1 vccd1 vccd1 _13677_/Z sky130_fd_sc_hd__ebufn_2
X_09897_ _09897_/A _09904_/Y vssd1 vssd1 vccd1 vccd1 _13817_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_69_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13526__D line[82] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XDATA\[3\].CLKBUF\[6\] clk vssd1 vssd1 vccd1 vccd1 _12177_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA_DATA\[26\].CLKBUF\[0\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08848_ _08850_/CLK line[120] vssd1 vssd1 vccd1 vccd1 _08849_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[27\].VALID\[11\].TOBUF OVHB\[27\].VALID\[11\].FF/Q OVHB\[27\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04915_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_84_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[0\].VALID\[14\].TOBUF OVHB\[0\].VALID\[14\].FF/Q OVHB\[0\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_72_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13823__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08779_ _08779_/A _08784_/Y vssd1 vssd1 vccd1 vccd1 _13819_/Z sky130_fd_sc_hd__ebufn_2
X_10810_ _10810_/CLK line[121] vssd1 vssd1 vccd1 vccd1 _10811_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[11\].CG clk OVHB\[11\].CGAND/X vssd1 vssd1 vccd1 vccd1 OVHB\[11\].V/CLK sky130_fd_sc_hd__dlclkp_1
X_11790_ _11790_/CLK line[57] vssd1 vssd1 vccd1 vccd1 _11791_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_25_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05044__D line[59] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06718__A _13905_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10741_ _10741_/A _10744_/Y vssd1 vssd1 vccd1 vccd1 _13821_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10885__D line[32] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MUX.M\[0\].MUX\[1\]_A3 _13840_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13460_ _13470_/CLK line[52] vssd1 vssd1 vccd1 vccd1 _13461_/A sky130_fd_sc_hd__dfxtp_1
X_10672_ _10672_/CLK _10673_/X vssd1 vssd1 vccd1 vccd1 _10670_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_201_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12411_ _12411_/A _12424_/Y vssd1 vssd1 vccd1 vccd1 _13811_/Z sky130_fd_sc_hd__ebufn_2
X_13391_ _13391_/A _13404_/Y vssd1 vssd1 vccd1 vccd1 _13671_/Z sky130_fd_sc_hd__ebufn_2
X_12342_ _12350_/CLK line[53] vssd1 vssd1 vccd1 vccd1 _12343_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_127_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12273_ _12273_/A _12284_/Y vssd1 vssd1 vccd1 vccd1 _13673_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_175_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09186__D line[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09764__A _13921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11224_ _11230_/CLK line[54] vssd1 vssd1 vccd1 vccd1 _11225_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[20\].VALID\[10\].TOBUF OVHB\[20\].VALID\[10\].FF/Q OVHB\[20\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04932_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_150_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10125__D line[78] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11155_ _11155_/A _11164_/Y vssd1 vssd1 vccd1 vccd1 _13675_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09483__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[25\].VALID\[6\].FF_D A[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05219__D line[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10106_ _10110_/CLK line[55] vssd1 vssd1 vccd1 vccd1 _10107_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_122_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11086_ _11090_/CLK line[119] vssd1 vssd1 vccd1 vccd1 _11087_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_76_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12340__D line[52] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10037_ _10037_/A _10044_/Y vssd1 vssd1 vccd1 vccd1 _13677_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_75_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07434__D line[113] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11988_ _12000_/CLK line[19] vssd1 vssd1 vccd1 vccd1 _11989_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[2\].CLKBUF\[3\] clk vssd1 vssd1 vccd1 vccd1 _11232_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_189_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13727_ _13727_/A _13754_/Y vssd1 vssd1 vccd1 vccd1 _13727_/Z sky130_fd_sc_hd__ebufn_2
X_10939_ _10939_/A _10954_/Y vssd1 vssd1 vccd1 vccd1 _13739_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_210_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13658_ _13680_/CLK line[29] vssd1 vssd1 vccd1 vccd1 _13659_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09939__A _13921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12609_ _12609_/A _12634_/Y vssd1 vssd1 vccd1 vccd1 _13729_/Z sky130_fd_sc_hd__ebufn_2
XPHY_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09658__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13589_ _13589_/A _13614_/Y vssd1 vssd1 vccd1 vccd1 _13869_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_185_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06130_ _06130_/A _06159_/Y vssd1 vssd1 vccd1 vccd1 _13690_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_117_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06061_ _06085_/CLK line[12] vssd1 vssd1 vccd1 vccd1 _06062_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12515__D line[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07609__D line[65] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05012_ _05012_/A _05039_/Y vssd1 vssd1 vccd1 vccd1 _13692_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_125_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09820_ _09830_/CLK line[52] vssd1 vssd1 vccd1 vccd1 _09821_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[8\].VALID\[9\].TOBUF OVHB\[8\].VALID\[9\].FF/Q OVHB\[8\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04914_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[6\].VALID\[11\].FF_D A[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09824__D line[54] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09751_ _09751_/A _09764_/Y vssd1 vssd1 vccd1 vccd1 _13671_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_140_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06963_ _13909_/Y wr vssd1 vssd1 vccd1 vccd1 _06963_/X sky130_fd_sc_hd__and2_1
XANTENNA__12250__D line[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08702_ _08710_/CLK line[53] vssd1 vssd1 vccd1 vccd1 _08703_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[22\].CLKBUF\[7\] clk vssd1 vssd1 vccd1 vccd1 _09132_/CLK sky130_fd_sc_hd__clkbuf_4
X_05914_ _13902_/X vssd1 vssd1 vccd1 vccd1 _05914_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09682_ _09690_/CLK line[117] vssd1 vssd1 vccd1 vccd1 _09683_/A sky130_fd_sc_hd__dfxtp_1
X_06894_ _13905_/X vssd1 vssd1 vccd1 vccd1 _06894_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08633_ _08633_/A _08644_/Y vssd1 vssd1 vccd1 vccd1 _13673_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_54_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05845_ _05875_/CLK line[32] vssd1 vssd1 vccd1 vccd1 _05846_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_199_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11444__A _13926_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08564_ _08570_/CLK line[118] vssd1 vssd1 vccd1 vccd1 _08565_/A sky130_fd_sc_hd__dfxtp_1
X_05776_ _05776_/A _05809_/Y vssd1 vssd1 vccd1 vccd1 _13616_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_120_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11163__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07515_ _07515_/A _07524_/Y vssd1 vssd1 vccd1 vccd1 _13675_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_81_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[6\].VALID\[1\].FF_D A[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13081__D line[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08495_ _08495_/A _08504_/Y vssd1 vssd1 vccd1 vccd1 _13815_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[6\].CG clk OVHB\[6\].CGAND/X vssd1 vssd1 vccd1 vccd1 OVHB\[6\].V/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__05799__D line[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08175__D line[68] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07446_ _07450_/CLK line[119] vssd1 vssd1 vccd1 vccd1 _07447_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_210_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XDATA\[1\].CLKBUF\[0\] clk vssd1 vssd1 vccd1 vccd1 _08047_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_210_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07377_ _07377_/A _07384_/Y vssd1 vssd1 vccd1 vccd1 _13817_/Z sky130_fd_sc_hd__ebufn_2
X_09116_ _09130_/CLK line[114] vssd1 vssd1 vccd1 vccd1 _09117_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_136_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06328_ _06330_/CLK line[120] vssd1 vssd1 vccd1 vccd1 _06329_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__04932__A1_N A_h[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09047_ _09047_/A _09064_/Y vssd1 vssd1 vccd1 vccd1 _13807_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12425__D line[96] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06259_ _06259_/A _06264_/Y vssd1 vssd1 vccd1 vccd1 _13819_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06423__D line[35] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11619__A _13926_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09734__D line[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09949_ _09949_/A _09974_/Y vssd1 vssd1 vccd1 vccd1 _13869_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.M\[1\].MUX\[6\]_A0 _13626_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11338__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13256__D line[87] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12960_ _12980_/CLK line[94] vssd1 vssd1 vccd1 vccd1 _12961_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_180_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11911_ _11911_/A _11934_/Y vssd1 vssd1 vccd1 vccd1 _13871_/Z sky130_fd_sc_hd__ebufn_2
X_12891_ _12891_/A _12914_/Y vssd1 vssd1 vccd1 vccd1 _13731_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_73_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11842_ _11860_/CLK line[95] vssd1 vssd1 vccd1 vccd1 _11843_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[21\].CLKBUF\[4\] clk vssd1 vssd1 vccd1 vccd1 _08747_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_54_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XOVHB\[15\].VALID\[4\].TOBUF OVHB\[15\].VALID\[4\].FF/Q OVHB\[15\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04925_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_54_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11773_ _11773_/A _11794_/Y vssd1 vssd1 vccd1 vccd1 _13733_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[24\].CLKBUF\[2\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11504__D line[54] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13512_ _13540_/CLK line[90] vssd1 vssd1 vccd1 vccd1 _13513_/A sky130_fd_sc_hd__dfxtp_1
X_10724_ _10740_/CLK line[81] vssd1 vssd1 vccd1 vccd1 _10725_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08085__D line[32] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13443_ _13443_/A _13474_/Y vssd1 vssd1 vccd1 vccd1 _13723_/Z sky130_fd_sc_hd__ebufn_2
X_10655_ _10655_/A _10674_/Y vssd1 vssd1 vccd1 vccd1 _13735_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09909__D line[107] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07279__A _13910_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13374_ _13400_/CLK line[27] vssd1 vssd1 vccd1 vccd1 _13375_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08813__D line[104] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10586_ _10600_/CLK line[18] vssd1 vssd1 vccd1 vccd1 _10587_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_186_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12325_ _12325_/A _12354_/Y vssd1 vssd1 vccd1 vccd1 _13725_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_5_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12913__A _13937_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12256_ _12280_/CLK line[28] vssd1 vssd1 vccd1 vccd1 _12257_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_123_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11207_ _11207_/A _11234_/Y vssd1 vssd1 vccd1 vccd1 _13727_/Z sky130_fd_sc_hd__ebufn_2
X_12187_ _12187_/A _12214_/Y vssd1 vssd1 vccd1 vccd1 _13867_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_205_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11138_ _11160_/CLK line[29] vssd1 vssd1 vccd1 vccd1 _11139_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_95_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13166__D line[60] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12070__D line[57] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11069_ _11069_/A _11094_/Y vssd1 vssd1 vccd1 vccd1 _13869_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07164__D line[118] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05630_ _05630_/CLK line[57] vssd1 vssd1 vccd1 vccd1 _05631_/A sky130_fd_sc_hd__dfxtp_1
X_05561_ _05561_/A _05564_/Y vssd1 vssd1 vccd1 vccd1 _13681_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11414__D line[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07300_ _07310_/CLK line[52] vssd1 vssd1 vccd1 vccd1 _07301_/A sky130_fd_sc_hd__dfxtp_1
X_05492_ _05492_/CLK _05493_/X vssd1 vssd1 vccd1 vccd1 _05490_/CLK sky130_fd_sc_hd__dlclkp_1
X_08280_ _08290_/CLK line[116] vssd1 vssd1 vccd1 vccd1 _08281_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08573__A _13913_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05412__D line[85] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDATA\[20\].CLKBUF\[1\] clk vssd1 vssd1 vccd1 vccd1 _08362_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_177_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07231_ _07231_/A _07244_/Y vssd1 vssd1 vccd1 vccd1 _13671_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_20_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07162_ _07170_/CLK line[117] vssd1 vssd1 vccd1 vccd1 _07163_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08723__D line[77] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDATA\[10\].CLKBUF\[7\] clk vssd1 vssd1 vccd1 vccd1 _05492_/CLK sky130_fd_sc_hd__clkbuf_4
XOVHB\[21\].VALID\[3\].TOBUF OVHB\[21\].VALID\[3\].FF/Q OVHB\[21\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04919_/B2 sky130_fd_sc_hd__ebufn_2
X_06113_ _06113_/A _06124_/Y vssd1 vssd1 vccd1 vccd1 _13673_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13919__A A[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07093_ _07093_/A _07104_/Y vssd1 vssd1 vccd1 vccd1 _13813_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12245__D line[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07339__D line[70] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06044_ _06050_/CLK line[118] vssd1 vssd1 vccd1 vccd1 _06045_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_114_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[8\].VALID\[7\].FF OVHB\[8\].V/CLK A[14] vssd1 vssd1 vccd1 vccd1 OVHB\[8\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_115_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09803_ _09803_/A _09834_/Y vssd1 vssd1 vccd1 vccd1 _13723_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[24\].CGAND_B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07995_ _07995_/A _08014_/Y vssd1 vssd1 vccd1 vccd1 _13875_/Z sky130_fd_sc_hd__ebufn_2
X_09734_ _09760_/CLK line[27] vssd1 vssd1 vccd1 vccd1 _09735_/A sky130_fd_sc_hd__dfxtp_1
X_06946_ _06960_/CLK line[18] vssd1 vssd1 vccd1 vccd1 _06947_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07074__D line[91] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08748__A _13914_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09665_ _09665_/A _09694_/Y vssd1 vssd1 vccd1 vccd1 _13865_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[9\].CGAND_B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06877_ _06877_/A _06894_/Y vssd1 vssd1 vccd1 vccd1 _13877_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[28\].CGAND_A _13924_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13804__D line[81] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08616_ _08640_/CLK line[28] vssd1 vssd1 vccd1 vccd1 _08617_/A sky130_fd_sc_hd__dfxtp_1
X_05828_ _05840_/CLK line[19] vssd1 vssd1 vccd1 vccd1 _05829_/A sky130_fd_sc_hd__dfxtp_1
X_09596_ _09620_/CLK line[92] vssd1 vssd1 vccd1 vccd1 _09597_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_131_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08547_ _08547_/A _08574_/Y vssd1 vssd1 vccd1 vccd1 _13867_/Z sky130_fd_sc_hd__ebufn_2
X_05759_ _05759_/A _05774_/Y vssd1 vssd1 vccd1 vccd1 _13879_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_152_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08478_ _08500_/CLK line[93] vssd1 vssd1 vccd1 vccd1 _08479_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05322__D line[58] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XOVHB\[25\].VALID\[14\].FF OVHB\[25\].V/CLK A[21] vssd1 vssd1 vccd1 vccd1 OVHB\[25\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07429_ _07429_/A _07454_/Y vssd1 vssd1 vccd1 vccd1 _13869_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_210_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10440_ _10460_/CLK line[94] vssd1 vssd1 vccd1 vccd1 _10441_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12155__D line[110] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10371_ _10371_/A _10394_/Y vssd1 vssd1 vccd1 vccd1 _13731_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07249__D line[43] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12110_ _12140_/CLK line[80] vssd1 vssd1 vccd1 vccd1 _12111_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_40_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06153__D line[40] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[21\].VALID\[9\].FF_D A[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13090_ _13120_/CLK line[16] vssd1 vssd1 vccd1 vccd1 _13091_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11994__D line[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XOVHB\[13\].VALID\[9\].TOBUF OVHB\[13\].VALID\[9\].FF/Q OVHB\[13\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04914_/B2 sky130_fd_sc_hd__ebufn_2
X_12041_ _12041_/A _12074_/Y vssd1 vssd1 vccd1 vccd1 _13721_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10253__A _13922_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09464__D line[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09033__TE_B _09064_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10403__D line[77] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12943_ _12945_/CLK line[72] vssd1 vssd1 vccd1 vccd1 _12944_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[6\].VALID\[9\].FF OVHB\[6\].V/CLK A[16] vssd1 vssd1 vccd1 vccd1 OVHB\[6\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_34_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12874_ _12874_/A _12879_/Y vssd1 vssd1 vccd1 vccd1 _13714_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07712__D line[127] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11825_ _11825_/CLK line[73] vssd1 vssd1 vccd1 vccd1 _11826_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06328__D line[120] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11756_ _11756_/A _11759_/Y vssd1 vssd1 vccd1 vccd1 _13716_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10707_ _10707_/CLK _10708_/X vssd1 vssd1 vccd1 vccd1 _10705_/CLK sky130_fd_sc_hd__dlclkp_1
XPHY_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11687_ _11687_/CLK _11688_/X vssd1 vssd1 vccd1 vccd1 _11685_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__10428__A _13923_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09639__D line[97] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13426_ _13426_/A _13439_/Y vssd1 vssd1 vccd1 vccd1 _13706_/Z sky130_fd_sc_hd__ebufn_2
X_10638_ _13924_/X wr vssd1 vssd1 vccd1 vccd1 _10638_/X sky130_fd_sc_hd__and2_1
XFILLER_10_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_DATA\[22\].CLKBUF\[4\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13357_ _13365_/CLK line[5] vssd1 vssd1 vccd1 vccd1 _13358_/A sky130_fd_sc_hd__dfxtp_1
X_10569_ _13924_/X vssd1 vssd1 vccd1 vccd1 _10569_/Y sky130_fd_sc_hd__inv_2
XANTENNA__06063__D line[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12308_ _12308_/A _12319_/Y vssd1 vssd1 vccd1 vccd1 _13708_/Z sky130_fd_sc_hd__ebufn_2
X_13288_ _13288_/A _13299_/Y vssd1 vssd1 vccd1 vccd1 _13848_/Z sky130_fd_sc_hd__ebufn_2
X_12239_ _12245_/CLK line[6] vssd1 vssd1 vccd1 vccd1 _12240_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13474__A _13898_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06800_ _06820_/CLK line[94] vssd1 vssd1 vccd1 vccd1 _06801_/A sky130_fd_sc_hd__dfxtp_1
X_07780_ _07800_/CLK line[30] vssd1 vssd1 vccd1 vccd1 _07781_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_68_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_04992_ _05000_/CLK line[21] vssd1 vssd1 vccd1 vccd1 _04993_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_83_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13193__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06731_ _06731_/A _06754_/Y vssd1 vssd1 vccd1 vccd1 _13731_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[2\].VALID\[4\].FF_D A[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09450_ _09480_/CLK line[16] vssd1 vssd1 vccd1 vccd1 _09451_/A sky130_fd_sc_hd__dfxtp_1
X_06662_ _06680_/CLK line[31] vssd1 vssd1 vccd1 vccd1 _06663_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06088__A _13903_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08401_ _08401_/A _08434_/Y vssd1 vssd1 vccd1 vccd1 _13721_/Z sky130_fd_sc_hd__ebufn_2
X_05613_ _05613_/A _05634_/Y vssd1 vssd1 vccd1 vccd1 _13733_/Z sky130_fd_sc_hd__ebufn_2
X_09381_ _09381_/A _09414_/Y vssd1 vssd1 vccd1 vccd1 _13861_/Z sky130_fd_sc_hd__ebufn_2
X_06593_ _06593_/A _06614_/Y vssd1 vssd1 vccd1 vccd1 _13873_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_196_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11144__D line[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08332_ _08360_/CLK line[26] vssd1 vssd1 vccd1 vccd1 _08333_/A sky130_fd_sc_hd__dfxtp_1
X_05544_ _05560_/CLK line[17] vssd1 vssd1 vccd1 vccd1 _05545_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06238__D line[93] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10983__D line[72] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08263_ _08263_/A _08294_/Y vssd1 vssd1 vccd1 vccd1 _13863_/Z sky130_fd_sc_hd__ebufn_2
X_05475_ _05475_/A _05494_/Y vssd1 vssd1 vccd1 vccd1 _13875_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.M\[3\].MUX\[7\]_A2 _13803_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07214_ _07240_/CLK line[27] vssd1 vssd1 vccd1 vccd1 _07215_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08453__D line[67] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08194_ _08220_/CLK line[91] vssd1 vssd1 vccd1 vccd1 _08195_/A sky130_fd_sc_hd__dfxtp_1
X_07145_ _07145_/A _07174_/Y vssd1 vssd1 vccd1 vccd1 _13865_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13649__A _13899_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07076_ _07100_/CLK line[92] vssd1 vssd1 vccd1 vccd1 _07077_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13368__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06027_ _06027_/A _06054_/Y vssd1 vssd1 vccd1 vccd1 _13867_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06701__D line[34] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11319__D line[97] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07978_ _13912_/X wr vssd1 vssd1 vccd1 vccd1 _07978_/X sky130_fd_sc_hd__and2_1
XANTENNA_MUX.M\[1\].MUX\[3\]_A3 _13830_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09717_ _09725_/CLK line[5] vssd1 vssd1 vccd1 vccd1 _09718_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_101_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06929_ _13909_/Y vssd1 vssd1 vccd1 vccd1 _06929_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13534__D line[86] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09648_ _09648_/A _09659_/Y vssd1 vssd1 vccd1 vccd1 _13848_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08628__D line[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[13\].VALID\[13\].FF_D A[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[13\].VALID\[14\].TOBUF OVHB\[13\].VALID\[14\].FF/Q OVHB\[13\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/B2 sky130_fd_sc_hd__ebufn_2
XOVHB\[15\].VALID\[1\].FF OVHB\[15\].V/CLK A[8] vssd1 vssd1 vccd1 vccd1 OVHB\[15\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_42_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09579_ _09585_/CLK line[70] vssd1 vssd1 vccd1 vccd1 _09580_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11610_ _11610_/A _11619_/Y vssd1 vssd1 vccd1 vccd1 _13850_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_42_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12590_ _12590_/A _12599_/Y vssd1 vssd1 vccd1 vccd1 _13710_/Z sky130_fd_sc_hd__ebufn_2
XPHY_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05052__D line[63] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10893__D line[45] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11541_ _11545_/CLK line[71] vssd1 vssd1 vccd1 vccd1 _11542_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XOVHB\[31\].VALID\[10\].FF OVHB\[31\].V/CLK A[17] vssd1 vssd1 vccd1 vccd1 OVHB\[31\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05987__D line[106] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[17\].VALID\[1\].FF_D A[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11472_ _11472_/A _11479_/Y vssd1 vssd1 vccd1 vccd1 _13712_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13211_ _13225_/CLK line[66] vssd1 vssd1 vccd1 vccd1 _13212_/A sky130_fd_sc_hd__dfxtp_1
X_10423_ _10425_/CLK line[72] vssd1 vssd1 vccd1 vccd1 _10424_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[3\].VALID\[0\].TOBUF OVHB\[3\].VALID\[0\].FF/Q OVHB\[3\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04924_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[23\].VALID\[12\].FF_D A[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13142_ _13142_/A _13159_/Y vssd1 vssd1 vccd1 vccd1 _13702_/Z sky130_fd_sc_hd__ebufn_2
X_10354_ _10354_/A _10359_/Y vssd1 vssd1 vccd1 vccd1 _13714_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[28\].VALID\[3\].TOBUF OVHB\[28\].VALID\[3\].FF/Q OVHB\[28\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04919_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__13709__D line[38] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13073_ _13085_/CLK line[3] vssd1 vssd1 vccd1 vccd1 _13074_/A sky130_fd_sc_hd__dfxtp_1
X_10285_ _10285_/CLK line[9] vssd1 vssd1 vccd1 vccd1 _10286_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09194__D line[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12024_ _12024_/A _12039_/Y vssd1 vssd1 vccd1 vccd1 _13704_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10133__D line[67] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[25\].VOBUF OVHB\[25\].V/Q OVHB\[25\].INV/Y vssd1 vssd1 vccd1 vccd1 _04912_/B1
+ sky130_fd_sc_hd__ebufn_2
XFILLER_93_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05227__D line[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13975_ _13982_/A _13982_/B _13982_/C _13982_/D vssd1 vssd1 vccd1 vccd1 _13975_/Y
+ sky130_fd_sc_hd__nor4b_4
XANTENNA__13444__D line[59] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[21\].VALID\[12\].FF OVHB\[21\].V/CLK A[19] vssd1 vssd1 vccd1 vccd1 OVHB\[21\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_202_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12926_ _12926_/A _12949_/Y vssd1 vssd1 vccd1 vccd1 _13766_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_202_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07442__D line[117] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12857_ _12875_/CLK line[47] vssd1 vssd1 vccd1 vccd1 _12858_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_61_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[8\].VALID\[8\].FF_D A[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11808_ _11808_/A _11829_/Y vssd1 vssd1 vccd1 vccd1 _13768_/Z sky130_fd_sc_hd__ebufn_2
X_12788_ _12788_/A _12809_/Y vssd1 vssd1 vccd1 vccd1 _13628_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11739_ _11755_/CLK line[33] vssd1 vssd1 vccd1 vccd1 _11740_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09369__D line[102] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05260_ _05280_/CLK line[30] vssd1 vssd1 vccd1 vccd1 _05261_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[13\].VALID\[3\].FF OVHB\[13\].V/CLK A[10] vssd1 vssd1 vccd1 vccd1 OVHB\[13\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10308__D line[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13409_ _13435_/CLK line[43] vssd1 vssd1 vccd1 vccd1 _13410_/A sky130_fd_sc_hd__dfxtp_1
X_05191_ _05191_/A _05214_/Y vssd1 vssd1 vccd1 vccd1 _13871_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[30\].VALID\[7\].FF OVHB\[30\].V/CLK A[14] vssd1 vssd1 vccd1 vccd1 OVHB\[30\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_155_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13619__D line[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12523__D line[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08950_ _08950_/A _08959_/Y vssd1 vssd1 vccd1 vccd1 _13710_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[11\].VALID\[14\].FF OVHB\[11\].V/CLK A[21] vssd1 vssd1 vccd1 vccd1 OVHB\[11\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07617__D line[69] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07901_ _07905_/CLK line[71] vssd1 vssd1 vccd1 vccd1 _07902_/A sky130_fd_sc_hd__dfxtp_1
X_08881_ _08885_/CLK line[7] vssd1 vssd1 vccd1 vccd1 _08882_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[20\].CLKBUF\[6\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07832_ _07832_/A _07839_/Y vssd1 vssd1 vccd1 vccd1 _13712_/Z sky130_fd_sc_hd__ebufn_2
X_07763_ _07765_/CLK line[8] vssd1 vssd1 vccd1 vccd1 _07764_/A sky130_fd_sc_hd__dfxtp_1
X_04975_ _04975_/A _05004_/Y vssd1 vssd1 vccd1 vccd1 _13655_/Z sky130_fd_sc_hd__ebufn_2
X_09502_ _09502_/A _09519_/Y vssd1 vssd1 vccd1 vccd1 _13702_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__04976__D line[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06714_ _06714_/A _06719_/Y vssd1 vssd1 vccd1 vccd1 _13714_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07694_ _07694_/A _07699_/Y vssd1 vssd1 vccd1 vccd1 _13854_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07352__D line[90] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09433_ _09445_/CLK line[3] vssd1 vssd1 vccd1 vccd1 _09434_/A sky130_fd_sc_hd__dfxtp_1
X_06645_ _06645_/CLK line[9] vssd1 vssd1 vccd1 vccd1 _06646_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_64_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09364_ _09364_/A _09379_/Y vssd1 vssd1 vccd1 vccd1 _13844_/Z sky130_fd_sc_hd__ebufn_2
X_06576_ _06576_/A _06579_/Y vssd1 vssd1 vccd1 vccd1 _13856_/Z sky130_fd_sc_hd__ebufn_2
X_08315_ _08325_/CLK line[4] vssd1 vssd1 vccd1 vccd1 _08316_/A sky130_fd_sc_hd__dfxtp_1
X_05527_ _05527_/CLK _05528_/X vssd1 vssd1 vccd1 vccd1 _05525_/CLK sky130_fd_sc_hd__dlclkp_1
X_09295_ _09305_/CLK line[68] vssd1 vssd1 vccd1 vccd1 _09296_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_32_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09279__D line[75] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08183__D line[72] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08246_ _08246_/A _08259_/Y vssd1 vssd1 vccd1 vccd1 _13846_/Z sky130_fd_sc_hd__ebufn_2
X_05458_ _13900_/X wr vssd1 vssd1 vccd1 vccd1 _05458_/X sky130_fd_sc_hd__and2_1
XOVHB\[29\].VALID\[8\].FF OVHB\[29\].V/CLK A[15] vssd1 vssd1 vccd1 vccd1 OVHB\[29\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__05600__D line[48] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08177_ _08185_/CLK line[69] vssd1 vssd1 vccd1 vccd1 _08178_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_180_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12283__A _13935_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05389_ _13900_/X vssd1 vssd1 vccd1 vccd1 _05389_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07128_ _07128_/A _07139_/Y vssd1 vssd1 vccd1 vccd1 _13848_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_134_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12433__D line[109] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07059_ _07065_/CLK line[70] vssd1 vssd1 vccd1 vccd1 _07060_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07527__D line[42] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[11\].VALID\[5\].FF OVHB\[11\].V/CLK A[12] vssd1 vssd1 vccd1 vccd1 OVHB\[11\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06431__D line[39] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10070_ _10070_/A _10079_/Y vssd1 vssd1 vccd1 vccd1 _13710_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11049__D line[102] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09742__D line[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08358__D line[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13760_ _13760_/A _13789_/Y vssd1 vssd1 vccd1 vccd1 _13760_/Z sky130_fd_sc_hd__ebufn_2
X_10972_ _10972_/A _10989_/Y vssd1 vssd1 vccd1 vccd1 _13772_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_46_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XOVHB\[1\].VALID\[5\].TOBUF OVHB\[1\].VALID\[5\].FF/Q OVHB\[1\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04927_/B2 sky130_fd_sc_hd__ebufn_2
X_12711_ _12735_/CLK line[108] vssd1 vssd1 vccd1 vccd1 _12712_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.M\[0\].MUX\[4\]_A1 _13706_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13691_ _13715_/CLK line[44] vssd1 vssd1 vccd1 vccd1 _13692_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_43_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12458__A _13935_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[26\].VALID\[8\].TOBUF OVHB\[26\].VALID\[8\].FF/Q OVHB\[26\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04931_/B2 sky130_fd_sc_hd__ebufn_2
XPHY_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12642_ _12642_/A _12669_/Y vssd1 vssd1 vccd1 vccd1 _13762_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_31_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12608__D line[61] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12573_ _12595_/CLK line[45] vssd1 vssd1 vccd1 vccd1 _12574_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11524_ _11524_/A _11549_/Y vssd1 vssd1 vccd1 vccd1 _13764_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08093__D line[45] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06606__D line[119] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11455_ _11475_/CLK line[46] vssd1 vssd1 vccd1 vccd1 _11456_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_172_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09917__D line[111] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10406_ _10406_/A _10429_/Y vssd1 vssd1 vccd1 vccd1 _13766_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_125_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11386_ _11386_/A _11409_/Y vssd1 vssd1 vccd1 vccd1 _13626_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_152_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13125_ _13155_/CLK line[32] vssd1 vssd1 vccd1 vccd1 _13126_/A sky130_fd_sc_hd__dfxtp_1
X_10337_ _10355_/CLK line[47] vssd1 vssd1 vccd1 vccd1 _10338_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_112_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_DATA\[19\].CLKBUF\[7\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06341__D line[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13056_ _13056_/A _13089_/Y vssd1 vssd1 vccd1 vccd1 _13616_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_140_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10268_ _10268_/A _10289_/Y vssd1 vssd1 vccd1 vccd1 _13628_/Z sky130_fd_sc_hd__ebufn_2
X_12007_ _12035_/CLK line[42] vssd1 vssd1 vccd1 vccd1 _12008_/A sky130_fd_sc_hd__dfxtp_1
X_10199_ _10215_/CLK line[97] vssd1 vssd1 vccd1 vccd1 _10200_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10798__D line[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13174__D line[49] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08268__D line[125] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13958_ _13960_/B _13960_/A _13960_/C _13960_/D vssd1 vssd1 vccd1 vccd1 _13958_/X
+ sky130_fd_sc_hd__and4b_4
X_12909_ _12909_/A _12914_/Y vssd1 vssd1 vccd1 vccd1 _13749_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_34_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13889_ _13889_/A _13894_/Y vssd1 vssd1 vccd1 vccd1 _13889_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[30\].CLKBUF\[6\] clk vssd1 vssd1 vccd1 vccd1 _11617_/CLK sky130_fd_sc_hd__clkbuf_4
X_06430_ _06430_/A _06439_/Y vssd1 vssd1 vccd1 vccd1 _13710_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_21_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06361_ _06365_/CLK line[7] vssd1 vssd1 vccd1 vccd1 _06362_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11422__D line[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08100_ _08100_/A _08119_/Y vssd1 vssd1 vccd1 vccd1 _13700_/Z sky130_fd_sc_hd__ebufn_2
X_05312_ _05312_/A _05319_/Y vssd1 vssd1 vccd1 vccd1 _13712_/Z sky130_fd_sc_hd__ebufn_2
X_09080_ _09080_/A _09099_/Y vssd1 vssd1 vccd1 vccd1 _13840_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06516__D line[92] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06292_ _06292_/A _06299_/Y vssd1 vssd1 vccd1 vccd1 _13852_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05420__D line[89] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08031_ _08045_/CLK line[2] vssd1 vssd1 vccd1 vccd1 _08032_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_163_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10038__D line[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05243_ _05245_/CLK line[8] vssd1 vssd1 vccd1 vccd1 _05244_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_128_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08731__D line[66] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05174_ _05174_/A _05179_/Y vssd1 vssd1 vccd1 vccd1 _13854_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13349__D line[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09982_ _09982_/A _10009_/Y vssd1 vssd1 vccd1 vccd1 _13622_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_89_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08933_ _08955_/CLK line[45] vssd1 vssd1 vccd1 vccd1 _08934_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[7\].VALID\[11\].TOBUF OVHB\[7\].VALID\[11\].FF/Q OVHB\[7\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04915_/B2 sky130_fd_sc_hd__ebufn_2
X_08864_ _08864_/A _08889_/Y vssd1 vssd1 vccd1 vccd1 _13624_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_96_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07815_ _07835_/CLK line[46] vssd1 vssd1 vccd1 vccd1 _07816_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_57_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_OVHB\[20\].VALID\[0\].FF_D A[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08795_ _08815_/CLK line[110] vssd1 vssd1 vccd1 vccd1 _08796_/A sky130_fd_sc_hd__dfxtp_1
X_07746_ _07746_/A _07769_/Y vssd1 vssd1 vccd1 vccd1 _13626_/Z sky130_fd_sc_hd__ebufn_2
X_04958_ _04958_/A _04969_/Y vssd1 vssd1 vccd1 vccd1 _13638_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07082__D line[95] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07677_ _07695_/CLK line[111] vssd1 vssd1 vccd1 vccd1 _07678_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_25_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13812__D line[85] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09416_ _09416_/A _09449_/Y vssd1 vssd1 vccd1 vccd1 _13616_/Z sky130_fd_sc_hd__ebufn_2
X_06628_ _06628_/A _06649_/Y vssd1 vssd1 vccd1 vccd1 _13628_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_25_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08906__D line[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[13\].VALID\[4\].FF_D A[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09347_ _09375_/CLK line[106] vssd1 vssd1 vccd1 vccd1 _09348_/A sky130_fd_sc_hd__dfxtp_1
X_06559_ _06575_/CLK line[97] vssd1 vssd1 vccd1 vccd1 _06560_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_139_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09278_ _09278_/A _09309_/Y vssd1 vssd1 vccd1 vccd1 _13758_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05330__D line[62] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08229_ _08255_/CLK line[107] vssd1 vssd1 vccd1 vccd1 _08230_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[9\].CG_CLK clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[0\].VALID\[10\].TOBUF OVHB\[0\].VALID\[10\].FF/Q OVHB\[0\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04932_/B2 sky130_fd_sc_hd__ebufn_2
X_11240_ _11240_/A _11269_/Y vssd1 vssd1 vccd1 vccd1 _13760_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_106_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12163__D line[99] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11171_ _11195_/CLK line[44] vssd1 vssd1 vccd1 vccd1 _11172_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07257__D line[47] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10122_ _10122_/A _10149_/Y vssd1 vssd1 vccd1 vccd1 _13762_/Z sky130_fd_sc_hd__ebufn_2
X_10053_ _10075_/CLK line[45] vssd1 vssd1 vccd1 vccd1 _10054_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09472__D line[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10411__D line[66] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13812_ _13820_/CLK line[85] vssd1 vssd1 vccd1 vccd1 _13813_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_180_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05505__D line[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13743_ _13743_/A _13754_/Y vssd1 vssd1 vccd1 vccd1 _13743_/Z sky130_fd_sc_hd__ebufn_2
X_10955_ _10985_/CLK line[64] vssd1 vssd1 vccd1 vccd1 _10956_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13722__D line[58] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13674_ _13680_/CLK line[22] vssd1 vssd1 vccd1 vccd1 _13675_/A sky130_fd_sc_hd__dfxtp_1
X_10886_ _10886_/A _10919_/Y vssd1 vssd1 vccd1 vccd1 _13686_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07720__D line[116] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12338__D line[51] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12625_ _12625_/A _12634_/Y vssd1 vssd1 vccd1 vccd1 _13745_/Z sky130_fd_sc_hd__ebufn_2
XPHY_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12556_ _12560_/CLK line[23] vssd1 vssd1 vccd1 vccd1 _12557_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11507_ _11507_/A _11514_/Y vssd1 vssd1 vccd1 vccd1 _13747_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12487_ _12487_/A _12494_/Y vssd1 vssd1 vccd1 vccd1 _13887_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09647__D line[101] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11438_ _11440_/CLK line[24] vssd1 vssd1 vccd1 vccd1 _11439_/A sky130_fd_sc_hd__dfxtp_1
X_11369_ _11369_/A _11374_/Y vssd1 vssd1 vccd1 vccd1 _13889_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_98_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06071__D line[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13108_ _13120_/CLK line[19] vssd1 vssd1 vccd1 vccd1 _13109_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12801__D line[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05930_ _05930_/A _05949_/Y vssd1 vssd1 vccd1 vccd1 _13770_/Z sky130_fd_sc_hd__ebufn_2
X_13039_ _13039_/A _13054_/Y vssd1 vssd1 vccd1 vccd1 _13879_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09382__D line[122] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05861_ _05875_/CLK line[34] vssd1 vssd1 vccd1 vccd1 _05862_/A sky130_fd_sc_hd__dfxtp_1
X_07600_ _07600_/A _07629_/Y vssd1 vssd1 vccd1 vccd1 _13760_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_208_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08580_ _08580_/A _08609_/Y vssd1 vssd1 vccd1 vccd1 _13620_/Z sky130_fd_sc_hd__ebufn_2
X_05792_ _05792_/A _05809_/Y vssd1 vssd1 vccd1 vccd1 _13632_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_66_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07531_ _07555_/CLK line[44] vssd1 vssd1 vccd1 vccd1 _07532_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[2\].VALID\[0\].FF OVHB\[2\].V/CLK A[7] vssd1 vssd1 vccd1 vccd1 OVHB\[2\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[26\].VALID\[4\].FF_D A[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[13\].CLKBUF\[0\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07462_ _07462_/A _07489_/Y vssd1 vssd1 vccd1 vccd1 _13622_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07630__D line[80] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09201_ _09201_/A _09204_/Y vssd1 vssd1 vccd1 vccd1 _13681_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_179_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06413_ _06435_/CLK line[45] vssd1 vssd1 vccd1 vccd1 _06414_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[8\].VALID\[5\].TOBUF OVHB\[8\].VALID\[5\].FF/Q OVHB\[8\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04927_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_210_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07393_ _07415_/CLK line[109] vssd1 vssd1 vccd1 vccd1 _07394_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11152__D line[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09132_ _09132_/CLK _09133_/X vssd1 vssd1 vccd1 vccd1 _09130_/CLK sky130_fd_sc_hd__dlclkp_1
X_06344_ _06344_/A _06369_/Y vssd1 vssd1 vccd1 vccd1 _13624_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06246__D line[82] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06824__A _13905_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[19\].VALID\[8\].FF_D A[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09063_ _13915_/X wr vssd1 vssd1 vccd1 vccd1 _09063_/X sky130_fd_sc_hd__and2_1
XFILLER_136_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06275_ _06295_/CLK line[110] vssd1 vssd1 vccd1 vccd1 _06276_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09557__D line[74] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06543__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08014_ _13912_/X vssd1 vssd1 vccd1 vccd1 _08014_/Y sky130_fd_sc_hd__inv_2
X_05226_ _05226_/A _05249_/Y vssd1 vssd1 vccd1 vccd1 _13626_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08461__D line[71] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[2\].VALID\[14\].FF OVHB\[2\].V/CLK A[21] vssd1 vssd1 vccd1 vccd1 OVHB\[2\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13079__D line[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MUX.M\[2\].MUX\[5\]_A3 _13883_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05157_ _05175_/CLK line[111] vssd1 vssd1 vccd1 vccd1 _05158_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[23\].VALID\[12\].TOBUF OVHB\[23\].VALID\[12\].FF/Q OVHB\[23\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04929_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_131_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_DATA\[6\].CLKBUF\[0\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09965_ _09965_/A _09974_/Y vssd1 vssd1 vccd1 vccd1 _13885_/Z sky130_fd_sc_hd__ebufn_2
X_05088_ _05088_/A _05109_/Y vssd1 vssd1 vccd1 vccd1 _13768_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12711__D line[108] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08916_ _08920_/CLK line[23] vssd1 vssd1 vccd1 vccd1 _08917_/A sky130_fd_sc_hd__dfxtp_1
X_09896_ _09900_/CLK line[87] vssd1 vssd1 vccd1 vccd1 _09897_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07805__D line[32] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08847_ _08847_/A _08854_/Y vssd1 vssd1 vccd1 vccd1 _13887_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11327__D line[101] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08778_ _08780_/CLK line[88] vssd1 vssd1 vccd1 vccd1 _08779_/A sky130_fd_sc_hd__dfxtp_1
X_07729_ _07729_/A _07734_/Y vssd1 vssd1 vccd1 vccd1 _13889_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06718__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10740_ _10740_/CLK line[89] vssd1 vssd1 vccd1 vccd1 _10741_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_41_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08636__D line[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10671_ _10671_/A _10674_/Y vssd1 vssd1 vccd1 vccd1 _13751_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11062__D line[122] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12410_ _12420_/CLK line[84] vssd1 vssd1 vccd1 vccd1 _12411_/A sky130_fd_sc_hd__dfxtp_1
X_13390_ _13400_/CLK line[20] vssd1 vssd1 vccd1 vccd1 _13391_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05060__D line[52] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[0\].VALID\[2\].FF OVHB\[0\].V/CLK A[9] vssd1 vssd1 vccd1 vccd1 OVHB\[0\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_12341_ _12341_/A _12354_/Y vssd1 vssd1 vccd1 vccd1 _13741_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_138_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05995__D line[110] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08371__D line[44] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12272_ _12280_/CLK line[21] vssd1 vssd1 vccd1 vccd1 _12273_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_4_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11223_ _11223_/A _11234_/Y vssd1 vssd1 vccd1 vccd1 _13743_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[15\].VALID\[0\].TOBUF OVHB\[15\].VALID\[0\].FF/Q OVHB\[15\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04924_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11154_ _11160_/CLK line[22] vssd1 vssd1 vccd1 vccd1 _11155_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_68_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XOVHB\[26\].VALID\[12\].FF OVHB\[26\].V/CLK A[19] vssd1 vssd1 vccd1 vccd1 OVHB\[26\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_122_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10105_ _10105_/A _10114_/Y vssd1 vssd1 vccd1 vccd1 _13745_/Z sky130_fd_sc_hd__ebufn_2
X_11085_ _11085_/A _11094_/Y vssd1 vssd1 vccd1 vccd1 _13885_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_0_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10036_ _10040_/CLK line[23] vssd1 vssd1 vccd1 vccd1 _10037_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_48_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11237__D line[74] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10141__D line[71] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05235__D line[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11987_ _11987_/A _12004_/Y vssd1 vssd1 vccd1 vccd1 _13667_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13452__D line[63] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13726_ _13750_/CLK line[60] vssd1 vssd1 vccd1 vccd1 _13727_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08546__D line[124] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10938_ _10950_/CLK line[51] vssd1 vssd1 vccd1 vccd1 _10939_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07450__D line[121] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12068__D line[56] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10869_ _10869_/A _10884_/Y vssd1 vssd1 vccd1 vccd1 _13669_/Z sky130_fd_sc_hd__ebufn_2
X_13657_ _13657_/A _13684_/Y vssd1 vssd1 vccd1 vccd1 _13657_/Z sky130_fd_sc_hd__ebufn_2
X_12608_ _12630_/CLK line[61] vssd1 vssd1 vccd1 vccd1 _12609_/A sky130_fd_sc_hd__dfxtp_1
XPHY_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13588_ _13610_/CLK line[125] vssd1 vssd1 vccd1 vccd1 _13589_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[16\].VALID\[14\].FF OVHB\[16\].V/CLK A[21] vssd1 vssd1 vccd1 vccd1 OVHB\[16\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_12539_ _12539_/A _12564_/Y vssd1 vssd1 vccd1 vccd1 _13659_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11700__D line[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06060_ _06060_/A _06089_/Y vssd1 vssd1 vccd1 vccd1 _13620_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_144_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05011_ _05035_/CLK line[44] vssd1 vssd1 vccd1 vccd1 _05012_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10316__D line[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13627__D line[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09750_ _09760_/CLK line[20] vssd1 vssd1 vccd1 vccd1 _09751_/A sky130_fd_sc_hd__dfxtp_1
X_06962_ _06962_/CLK _06963_/X vssd1 vssd1 vccd1 vccd1 _06960_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__07625__D line[73] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08701_ _08701_/A _08714_/Y vssd1 vssd1 vccd1 vccd1 _13741_/Z sky130_fd_sc_hd__ebufn_2
X_05913_ _13902_/X wr vssd1 vssd1 vccd1 vccd1 _05913_/X sky130_fd_sc_hd__and2_1
X_09681_ _09681_/A _09694_/Y vssd1 vssd1 vccd1 vccd1 _13881_/Z sky130_fd_sc_hd__ebufn_2
X_06893_ _13905_/X wr vssd1 vssd1 vccd1 vccd1 _06893_/X sky130_fd_sc_hd__and2_1
XFILLER_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08632_ _08640_/CLK line[21] vssd1 vssd1 vccd1 vccd1 _08633_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_54_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10051__D line[44] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05844_ _13902_/X vssd1 vssd1 vccd1 vccd1 _05844_/Y sky130_fd_sc_hd__inv_2
XANTENNA__05145__D line[96] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08563_ _08563_/A _08574_/Y vssd1 vssd1 vccd1 vccd1 _13883_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05775_ _05805_/CLK line[0] vssd1 vssd1 vccd1 vccd1 _05776_/A sky130_fd_sc_hd__dfxtp_1
X_07514_ _07520_/CLK line[22] vssd1 vssd1 vccd1 vccd1 _07515_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13940__A A_h[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__04984__D line[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08494_ _08500_/CLK line[86] vssd1 vssd1 vccd1 vccd1 _08495_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_211_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07360__D line[94] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07445_ _07445_/A _07454_/Y vssd1 vssd1 vccd1 vccd1 _13885_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_50_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07376_ _07380_/CLK line[87] vssd1 vssd1 vccd1 vccd1 _07377_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_13_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09115_ _09115_/A _09134_/Y vssd1 vssd1 vccd1 vccd1 _13875_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[11\].CLKBUF\[2\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06327_ _06327_/A _06334_/Y vssd1 vssd1 vccd1 vccd1 _13887_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09287__D line[79] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09046_ _09060_/CLK line[82] vssd1 vssd1 vccd1 vccd1 _09047_/A sky130_fd_sc_hd__dfxtp_1
X_06258_ _06260_/CLK line[88] vssd1 vssd1 vccd1 vccd1 _06259_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_190_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10226__D line[124] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05209_ _05209_/A _05214_/Y vssd1 vssd1 vccd1 vccd1 _13889_/Z sky130_fd_sc_hd__ebufn_2
X_06189_ _06189_/A _06194_/Y vssd1 vssd1 vccd1 vccd1 _13749_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_1_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[0\].VALID\[12\].FF_D A[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12441__D line[98] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__04929__A2_N _04929_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09948_ _09970_/CLK line[125] vssd1 vssd1 vccd1 vccd1 _09949_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.M\[1\].MUX\[6\]_A1 _13696_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07535__D line[46] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09879_ _09879_/A _09904_/Y vssd1 vssd1 vccd1 vccd1 _13799_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_38_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11910_ _11930_/CLK line[126] vssd1 vssd1 vccd1 vccd1 _11911_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_38_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_DATA\[4\].CLKBUF\[2\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12890_ _12910_/CLK line[62] vssd1 vssd1 vccd1 vccd1 _12891_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09750__D line[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05633__A _13901_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11841_ _11841_/A _11864_/Y vssd1 vssd1 vccd1 vccd1 _13801_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_33_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11772_ _11790_/CLK line[63] vssd1 vssd1 vccd1 vccd1 _11773_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[13\].VALID\[5\].TOBUF OVHB\[13\].VALID\[5\].FF/Q OVHB\[13\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04927_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_202_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_DATA\[30\].CLKBUF\[4\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10723_ _10723_/A _10744_/Y vssd1 vssd1 vccd1 vccd1 _13803_/Z sky130_fd_sc_hd__ebufn_2
X_13511_ _13511_/A _13544_/Y vssd1 vssd1 vccd1 vccd1 _13791_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_159_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13442_ _13470_/CLK line[58] vssd1 vssd1 vccd1 vccd1 _13443_/A sky130_fd_sc_hd__dfxtp_1
X_10654_ _10670_/CLK line[49] vssd1 vssd1 vccd1 vccd1 _10655_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_70_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13373_ _13373_/A _13404_/Y vssd1 vssd1 vccd1 vccd1 _13653_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12616__D line[50] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10585_ _10585_/A _10604_/Y vssd1 vssd1 vccd1 vccd1 _13665_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_139_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12324_ _12350_/CLK line[59] vssd1 vssd1 vccd1 vccd1 _12325_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12913__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12255_ _12255_/A _12284_/Y vssd1 vssd1 vccd1 vccd1 _13655_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_79_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09925__D line[100] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11206_ _11230_/CLK line[60] vssd1 vssd1 vccd1 vccd1 _11207_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05808__A _13902_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12186_ _12210_/CLK line[124] vssd1 vssd1 vccd1 vccd1 _12187_/A sky130_fd_sc_hd__dfxtp_1
X_11137_ _11137_/A _11164_/Y vssd1 vssd1 vccd1 vccd1 _13657_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_205_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11068_ _11090_/CLK line[125] vssd1 vssd1 vccd1 vccd1 _11069_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_48_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10019_ _10019_/A _10044_/Y vssd1 vssd1 vccd1 vccd1 _13659_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[22\].VALID\[7\].FF_D A[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09660__D line[112] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13182__D line[53] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05560_ _05560_/CLK line[25] vssd1 vssd1 vccd1 vccd1 _05561_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08276__D line[114] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08854__A _13914_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13709_ _13715_/CLK line[38] vssd1 vssd1 vccd1 vccd1 _13710_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_177_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05491_ _05491_/A _05494_/Y vssd1 vssd1 vccd1 vccd1 _13891_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08573__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07230_ _07240_/CLK line[20] vssd1 vssd1 vccd1 vccd1 _07231_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_149_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07161_ _07161_/A _07174_/Y vssd1 vssd1 vccd1 vccd1 _13881_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_164_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XOVHB\[22\].VALID\[10\].FF OVHB\[22\].V/CLK A[17] vssd1 vssd1 vccd1 vccd1 OVHB\[22\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11430__D line[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06112_ _06120_/CLK line[21] vssd1 vssd1 vccd1 vccd1 _06113_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06524__D line[81] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07092_ _07100_/CLK line[85] vssd1 vssd1 vccd1 vccd1 _07093_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_145_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06043_ _06043_/A _06054_/Y vssd1 vssd1 vccd1 vccd1 _13883_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_172_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09835__D line[64] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13357__D line[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09802_ _09830_/CLK line[58] vssd1 vssd1 vccd1 vccd1 _09803_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_115_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07994_ _08010_/CLK line[113] vssd1 vssd1 vccd1 vccd1 _07995_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[23\].VALID\[1\].FF OVHB\[23\].V/CLK A[8] vssd1 vssd1 vccd1 vccd1 OVHB\[23\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_06945_ _06945_/A _06964_/Y vssd1 vssd1 vccd1 vccd1 _13665_/Z sky130_fd_sc_hd__ebufn_2
X_09733_ _09733_/A _09764_/Y vssd1 vssd1 vccd1 vccd1 _13653_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_86_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08748__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09664_ _09690_/CLK line[123] vssd1 vssd1 vccd1 vccd1 _09665_/A sky130_fd_sc_hd__dfxtp_1
X_06876_ _06890_/CLK line[114] vssd1 vssd1 vccd1 vccd1 _06877_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[28\].CGAND_B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08615_ _08615_/A _08644_/Y vssd1 vssd1 vccd1 vccd1 _13655_/Z sky130_fd_sc_hd__ebufn_2
X_05827_ _05827_/A _05844_/Y vssd1 vssd1 vccd1 vccd1 _13667_/Z sky130_fd_sc_hd__ebufn_2
X_09595_ _09595_/A _09624_/Y vssd1 vssd1 vccd1 vccd1 _13795_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13092__D line[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11605__D line[100] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XOVHB\[12\].VALID\[12\].FF OVHB\[12\].V/CLK A[19] vssd1 vssd1 vccd1 vccd1 OVHB\[12\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_DATA\[29\].CLKBUF\[5\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08546_ _08570_/CLK line[124] vssd1 vssd1 vccd1 vccd1 _08547_/A sky130_fd_sc_hd__dfxtp_1
X_05758_ _05770_/CLK line[115] vssd1 vssd1 vccd1 vccd1 _05759_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07090__D line[84] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08477_ _08477_/A _08504_/Y vssd1 vssd1 vccd1 vccd1 _13797_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_23_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05689_ _05689_/A _05704_/Y vssd1 vssd1 vccd1 vccd1 _13809_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13820__D line[89] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07428_ _07450_/CLK line[125] vssd1 vssd1 vccd1 vccd1 _07429_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08914__D line[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[3\].VALID\[2\].FF_D A[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07359_ _07359_/A _07384_/Y vssd1 vssd1 vccd1 vccd1 _13799_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11340__D line[112] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10370_ _10390_/CLK line[62] vssd1 vssd1 vccd1 vccd1 _10371_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_40_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09029_ _13915_/X vssd1 vssd1 vccd1 vccd1 _09029_/Y sky130_fd_sc_hd__inv_2
XOVHB\[13\].VALID\[10\].TOBUF OVHB\[13\].VALID\[10\].FF/Q OVHB\[13\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04932_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_108_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10534__A _13923_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12040_ _12070_/CLK line[48] vssd1 vssd1 vccd1 vccd1 _12041_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_104_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10253__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13267__D line[106] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12171__D line[103] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07265__D line[36] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12942_ _12942_/A _12949_/Y vssd1 vssd1 vccd1 vccd1 _13782_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09480__D line[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12873_ _12875_/CLK line[40] vssd1 vssd1 vccd1 vccd1 _12874_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11515__D line[64] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XOVHB\[21\].VALID\[3\].FF OVHB\[21\].V/CLK A[10] vssd1 vssd1 vccd1 vccd1 OVHB\[21\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_11824_ _11824_/A _11829_/Y vssd1 vssd1 vccd1 vccd1 _13784_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_45_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05513__D line[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11755_ _11755_/CLK line[41] vssd1 vssd1 vccd1 vccd1 _11756_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13730__D line[62] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10709__A _13924_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[2\].CLKBUF\[4\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10706_ _10706_/A _10709_/Y vssd1 vssd1 vccd1 vccd1 _13786_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08824__D line[123] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06194__A _13903_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11686_ _11686_/A _11689_/Y vssd1 vssd1 vccd1 vccd1 _13646_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10428__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[21\].VOBUF OVHB\[21\].V/Q OVHB\[21\].INV/Y vssd1 vssd1 vccd1 vccd1 _04912_/B1
+ sky130_fd_sc_hd__ebufn_2
XPHY_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12346__D line[55] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13425_ _13435_/CLK line[36] vssd1 vssd1 vccd1 vccd1 _13426_/A sky130_fd_sc_hd__dfxtp_1
X_10637_ _10637_/CLK _10638_/X vssd1 vssd1 vccd1 vccd1 _10635_/CLK sky130_fd_sc_hd__dlclkp_1
XOVHB\[24\].CG clk OVHB\[24\].CGAND/X vssd1 vssd1 vccd1 vccd1 OVHB\[24\].V/CLK sky130_fd_sc_hd__dlclkp_1
X_13356_ _13356_/A _13369_/Y vssd1 vssd1 vccd1 vccd1 _13636_/Z sky130_fd_sc_hd__ebufn_2
X_10568_ _13924_/X wr vssd1 vssd1 vccd1 vccd1 _10568_/X sky130_fd_sc_hd__and2_1
XFILLER_127_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12307_ _12315_/CLK line[37] vssd1 vssd1 vccd1 vccd1 _12308_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_155_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10499_ _13923_/X vssd1 vssd1 vccd1 vccd1 _10499_/Y sky130_fd_sc_hd__inv_2
X_13287_ _13295_/CLK line[101] vssd1 vssd1 vccd1 vccd1 _13288_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09655__D line[105] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12238_ _12238_/A _12249_/Y vssd1 vssd1 vccd1 vccd1 _13638_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_107_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12081__D line[76] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12169_ _12175_/CLK line[102] vssd1 vssd1 vccd1 vccd1 _12170_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_68_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07175__D line[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_04991_ _04991_/A _05004_/Y vssd1 vssd1 vccd1 vccd1 _13671_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[7\].VALID\[12\].FF_D A[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06730_ _06750_/CLK line[62] vssd1 vssd1 vccd1 vccd1 _06731_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_37_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09390__D line[126] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06369__A _13904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07903__D line[72] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__04931__A1_N A_h[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06661_ _06661_/A _06684_/Y vssd1 vssd1 vccd1 vccd1 _13661_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06088__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08400_ _08430_/CLK line[48] vssd1 vssd1 vccd1 vccd1 _08401_/A sky130_fd_sc_hd__dfxtp_1
X_05612_ _05630_/CLK line[63] vssd1 vssd1 vccd1 vccd1 _05613_/A sky130_fd_sc_hd__dfxtp_1
X_09380_ _09410_/CLK line[112] vssd1 vssd1 vccd1 vccd1 _09381_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_36_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06592_ _06610_/CLK line[127] vssd1 vssd1 vccd1 vccd1 _06593_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_33_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08331_ _08331_/A _08364_/Y vssd1 vssd1 vccd1 vccd1 _13651_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_51_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05543_ _05543_/A _05564_/Y vssd1 vssd1 vccd1 vccd1 _13663_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[7\].VALID\[14\].FF OVHB\[7\].V/CLK A[21] vssd1 vssd1 vccd1 vccd1 OVHB\[7\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_08262_ _08290_/CLK line[122] vssd1 vssd1 vccd1 vccd1 _08263_/A sky130_fd_sc_hd__dfxtp_1
X_05474_ _05490_/CLK line[113] vssd1 vssd1 vccd1 vccd1 _05475_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.M\[3\].MUX\[7\]_A3 _13873_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07213_ _07213_/A _07244_/Y vssd1 vssd1 vccd1 vccd1 _13653_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12256__D line[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08193_ _08193_/A _08224_/Y vssd1 vssd1 vccd1 vccd1 _13793_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11160__D line[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07144_ _07170_/CLK line[123] vssd1 vssd1 vccd1 vccd1 _07145_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06254__D line[86] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07075_ _07075_/A _07104_/Y vssd1 vssd1 vccd1 vccd1 _13795_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[9\].VALID\[6\].FF_D A[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09565__D line[78] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06026_ _06050_/CLK line[124] vssd1 vssd1 vccd1 vccd1 _06027_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_99_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10504__D line[123] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07663__A _13911_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07977_ _07977_/CLK _07978_/X vssd1 vssd1 vccd1 vccd1 _07975_/CLK sky130_fd_sc_hd__dlclkp_1
X_09716_ _09716_/A _09729_/Y vssd1 vssd1 vccd1 vccd1 _13636_/Z sky130_fd_sc_hd__ebufn_2
X_06928_ _13909_/Y wr vssd1 vssd1 vccd1 vccd1 _06928_/X sky130_fd_sc_hd__and2_1
XFILLER_74_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07813__D line[45] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09647_ _09655_/CLK line[101] vssd1 vssd1 vccd1 vccd1 _09648_/A sky130_fd_sc_hd__dfxtp_1
X_06859_ _13905_/X vssd1 vssd1 vccd1 vccd1 _06859_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11335__D line[105] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06429__D line[38] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09578_ _09578_/A _09589_/Y vssd1 vssd1 vccd1 vccd1 _13778_/Z sky130_fd_sc_hd__ebufn_2
XPHY_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08529_ _08535_/CLK line[102] vssd1 vssd1 vccd1 vccd1 _08530_/A sky130_fd_sc_hd__dfxtp_1
XPHY_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11540_ _11540_/A _11549_/Y vssd1 vssd1 vccd1 vccd1 _13780_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XOVHB\[18\].VALID\[6\].FF OVHB\[18\].V/CLK A[13] vssd1 vssd1 vccd1 vccd1 OVHB\[18\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11471_ _11475_/CLK line[39] vssd1 vssd1 vccd1 vccd1 _11472_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[27\].CLKBUF\[7\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11070__D line[126] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06164__D line[59] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10422_ _10422_/A _10429_/Y vssd1 vssd1 vccd1 vccd1 _13782_/Z sky130_fd_sc_hd__ebufn_2
X_13210_ _13210_/A _13229_/Y vssd1 vssd1 vccd1 vccd1 _13770_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07838__A _13912_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10353_ _10355_/CLK line[40] vssd1 vssd1 vccd1 vccd1 _10354_/A sky130_fd_sc_hd__dfxtp_1
X_13141_ _13155_/CLK line[34] vssd1 vssd1 vccd1 vccd1 _13142_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[1\].VALID\[1\].TOBUF OVHB\[1\].VALID\[1\].FF/Q OVHB\[1\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04926_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_124_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13072_ _13072_/A _13089_/Y vssd1 vssd1 vccd1 vccd1 _13632_/Z sky130_fd_sc_hd__ebufn_2
X_10284_ _10284_/A _10289_/Y vssd1 vssd1 vccd1 vccd1 _13644_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[26\].VALID\[4\].TOBUF OVHB\[26\].VALID\[4\].FF/Q OVHB\[26\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04925_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_183_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12023_ _12035_/CLK line[35] vssd1 vssd1 vccd1 vccd1 _12024_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_3_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13974_ A_h[2] vssd1 vssd1 vccd1 vccd1 _13982_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_206_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12925_ _12945_/CLK line[78] vssd1 vssd1 vccd1 vccd1 _12926_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_34_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11245__D line[78] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06339__D line[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12856_ _12856_/A _12879_/Y vssd1 vssd1 vccd1 vccd1 _13696_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[10\].CGAND_A _13900_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05243__D line[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11807_ _11825_/CLK line[79] vssd1 vssd1 vccd1 vccd1 _11808_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12787_ _12805_/CLK line[15] vssd1 vssd1 vccd1 vccd1 _12788_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13460__D line[52] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08554__D line[113] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11738_ _11738_/A _11759_/Y vssd1 vssd1 vccd1 vccd1 _13698_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_159_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[28\].CGAND _13924_/X wr vssd1 vssd1 vccd1 vccd1 OVHB\[28\].CGAND/X sky130_fd_sc_hd__and2_4
X_11669_ _11685_/CLK line[1] vssd1 vssd1 vccd1 vccd1 _11670_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13408_ _13408_/A _13439_/Y vssd1 vssd1 vccd1 vccd1 _13688_/Z sky130_fd_sc_hd__ebufn_2
X_05190_ _05210_/CLK line[126] vssd1 vssd1 vccd1 vccd1 _05191_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_155_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_DATA\[0\].CLKBUF\[6\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XOVHB\[2\].V OVHB\[2\].V/CLK TIE/HI rst_n vssd1 vssd1 vccd1 vccd1 OVHB\[2\].V/Q sky130_fd_sc_hd__dfrtp_1
X_13339_ _13365_/CLK line[11] vssd1 vssd1 vccd1 vccd1 _13340_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06802__D line[95] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[16\].VALID\[8\].FF OVHB\[16\].V/CLK A[15] vssd1 vssd1 vccd1 vccd1 OVHB\[16\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_69_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07900_ _07900_/A _07909_/Y vssd1 vssd1 vccd1 vccd1 _13780_/Z sky130_fd_sc_hd__ebufn_2
X_08880_ _08880_/A _08889_/Y vssd1 vssd1 vccd1 vccd1 _13640_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_96_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05418__D line[88] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07831_ _07835_/CLK line[39] vssd1 vssd1 vccd1 vccd1 _07832_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_96_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13635__D line[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_04974_ _05000_/CLK line[27] vssd1 vssd1 vccd1 vccd1 _04975_/A sky130_fd_sc_hd__dfxtp_1
X_07762_ _07762_/A _07769_/Y vssd1 vssd1 vccd1 vccd1 _13642_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08729__D line[65] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09501_ _09515_/CLK line[34] vssd1 vssd1 vccd1 vccd1 _09502_/A sky130_fd_sc_hd__dfxtp_1
X_06713_ _06715_/CLK line[40] vssd1 vssd1 vccd1 vccd1 _06714_/A sky130_fd_sc_hd__dfxtp_1
X_07693_ _07695_/CLK line[104] vssd1 vssd1 vccd1 vccd1 _07694_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_37_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09432_ _09432_/A _09449_/Y vssd1 vssd1 vccd1 vccd1 _13632_/Z sky130_fd_sc_hd__ebufn_2
X_06644_ _06644_/A _06649_/Y vssd1 vssd1 vccd1 vccd1 _13644_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05153__D line[109] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09203__A _13916_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10994__D line[91] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09363_ _09375_/CLK line[99] vssd1 vssd1 vccd1 vccd1 _09364_/A sky130_fd_sc_hd__dfxtp_1
X_06575_ _06575_/CLK line[105] vssd1 vssd1 vccd1 vccd1 _06576_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13370__D line[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__04992__D line[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05526_ _05526_/A _05529_/Y vssd1 vssd1 vccd1 vccd1 _13646_/Z sky130_fd_sc_hd__ebufn_2
X_08314_ _08314_/A _08329_/Y vssd1 vssd1 vccd1 vccd1 _13634_/Z sky130_fd_sc_hd__ebufn_2
X_09294_ _09294_/A _09309_/Y vssd1 vssd1 vccd1 vccd1 _13774_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_166_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08245_ _08255_/CLK line[100] vssd1 vssd1 vccd1 vccd1 _08246_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_177_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05457_ _05457_/CLK _05458_/X vssd1 vssd1 vccd1 vccd1 _05455_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__12564__A _13936_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08176_ _08176_/A _08189_/Y vssd1 vssd1 vccd1 vccd1 _13776_/Z sky130_fd_sc_hd__ebufn_2
X_05388_ _13900_/X wr vssd1 vssd1 vccd1 vccd1 _05388_/X sky130_fd_sc_hd__and2_1
XANTENNA__12283__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07127_ _07135_/CLK line[101] vssd1 vssd1 vccd1 vccd1 _07128_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_106_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09047__TE_B _09064_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09295__D line[68] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05178__A _13931_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07058_ _07058_/A _07069_/Y vssd1 vssd1 vccd1 vccd1 _13778_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_161_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06009_ _06015_/CLK line[102] vssd1 vssd1 vccd1 vccd1 _06010_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10234__D line[113] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05328__D line[61] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13545__D line[96] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[3\].VALID\[12\].FF OVHB\[3\].V/CLK A[19] vssd1 vssd1 vccd1 vccd1 OVHB\[3\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07543__D line[35] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10971_ _10985_/CLK line[66] vssd1 vssd1 vccd1 vccd1 _10972_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_90_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12739__A _13936_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12710_ _12710_/A _12739_/Y vssd1 vssd1 vccd1 vccd1 _13830_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_43_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_MUX.M\[0\].MUX\[4\]_A2 _13776_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13690_ _13690_/A _13719_/Y vssd1 vssd1 vccd1 vccd1 _13690_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12458__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12641_ _12665_/CLK line[76] vssd1 vssd1 vccd1 vccd1 _12642_/A sky130_fd_sc_hd__dfxtp_1
XPHY_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[24\].VALID\[9\].TOBUF OVHB\[24\].VALID\[9\].FF/Q OVHB\[24\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04914_/B2 sky130_fd_sc_hd__ebufn_2
XPHY_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12572_ _12572_/A _12599_/Y vssd1 vssd1 vccd1 vccd1 _13692_/Z sky130_fd_sc_hd__ebufn_2
XPHY_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11523_ _11545_/CLK line[77] vssd1 vssd1 vccd1 vccd1 _11524_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10409__D line[65] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11454_ _11454_/A _11479_/Y vssd1 vssd1 vccd1 vccd1 _13694_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_156_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10405_ _10425_/CLK line[78] vssd1 vssd1 vccd1 vccd1 _10406_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12624__D line[54] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11385_ _11405_/CLK line[14] vssd1 vssd1 vccd1 vccd1 _11386_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_180_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07718__D line[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[14\].VALID\[2\].FF_D A[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13124_ _13938_/X vssd1 vssd1 vccd1 vccd1 _13124_/Y sky130_fd_sc_hd__inv_2
XDATA\[9\].CLKBUF\[0\] clk vssd1 vssd1 vccd1 vccd1 _13647_/CLK sky130_fd_sc_hd__clkbuf_4
X_10336_ _10336_/A _10359_/Y vssd1 vssd1 vccd1 vccd1 _13696_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_112_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10267_ _10285_/CLK line[15] vssd1 vssd1 vccd1 vccd1 _10268_/A sky130_fd_sc_hd__dfxtp_1
X_13055_ _13085_/CLK line[0] vssd1 vssd1 vccd1 vccd1 _13056_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_87_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08399__A _13913_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09933__D line[104] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12006_ _12006_/A _12039_/Y vssd1 vssd1 vccd1 vccd1 _13686_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_120_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10198_ _10198_/A _10219_/Y vssd1 vssd1 vccd1 vccd1 _13838_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[21\].CLKBUF\[0\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13957_ _13960_/A _13960_/B _13960_/C _13960_/D vssd1 vssd1 vccd1 vccd1 _13957_/X
+ sky130_fd_sc_hd__and4bb_4
XFILLER_74_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06069__D line[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12908_ _12910_/CLK line[56] vssd1 vssd1 vccd1 vccd1 _12909_/A sky130_fd_sc_hd__dfxtp_1
X_13888_ _13890_/CLK line[120] vssd1 vssd1 vccd1 vccd1 _13889_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_61_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XOVHB\[27\].VALID\[10\].FF OVHB\[27\].V/CLK A[17] vssd1 vssd1 vccd1 vccd1 OVHB\[27\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_12839_ _12839_/A _12844_/Y vssd1 vssd1 vccd1 vccd1 _13679_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_21_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13190__D line[57] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06360_ _06360_/A _06369_/Y vssd1 vssd1 vccd1 vccd1 _13640_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08284__D line[118] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05311_ _05315_/CLK line[39] vssd1 vssd1 vccd1 vccd1 _05312_/A sky130_fd_sc_hd__dfxtp_1
X_06291_ _06295_/CLK line[103] vssd1 vssd1 vccd1 vccd1 _06292_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[29\].CLKBUF\[4\] clk vssd1 vssd1 vccd1 vccd1 _10987_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA_OVHB\[5\].VALID\[9\].FF_D A[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08030_ _08030_/A _08049_/Y vssd1 vssd1 vccd1 vccd1 _13630_/Z sky130_fd_sc_hd__ebufn_2
X_05242_ _05242_/A _05249_/Y vssd1 vssd1 vccd1 vccd1 _13642_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_174_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XOVHB\[3\].VALID\[12\].TOBUF OVHB\[3\].VALID\[12\].FF/Q OVHB\[3\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04929_/B2 sky130_fd_sc_hd__ebufn_2
X_05173_ _05175_/CLK line[104] vssd1 vssd1 vccd1 vccd1 _05174_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12534__D line[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09693__A _13920_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06532__D line[85] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[30\].VALID\[8\].TOBUF OVHB\[30\].VALID\[8\].FF/Q OVHB\[30\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04931_/B2 sky130_fd_sc_hd__ebufn_2
X_09981_ _10005_/CLK line[12] vssd1 vssd1 vccd1 vccd1 _09982_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_116_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08932_ _08932_/A _08959_/Y vssd1 vssd1 vccd1 vccd1 _13692_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_115_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[9\].VALID\[1\].FF OVHB\[9\].V/CLK A[8] vssd1 vssd1 vccd1 vccd1 OVHB\[9\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XOVHB\[8\].VALID\[1\].TOBUF OVHB\[8\].VALID\[1\].FF/Q OVHB\[8\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04926_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__09843__D line[77] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08863_ _08885_/CLK line[13] vssd1 vssd1 vccd1 vccd1 _08864_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[17\].VALID\[12\].FF OVHB\[17\].V/CLK A[19] vssd1 vssd1 vccd1 vccd1 OVHB\[17\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13365__D line[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07814_ _07814_/A _07839_/Y vssd1 vssd1 vccd1 vccd1 _13694_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_123_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08459__D line[70] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08794_ _08794_/A _08819_/Y vssd1 vssd1 vccd1 vccd1 _13834_/Z sky130_fd_sc_hd__ebufn_2
X_04957_ _04965_/CLK line[5] vssd1 vssd1 vccd1 vccd1 _04958_/A sky130_fd_sc_hd__dfxtp_1
X_07745_ _07765_/CLK line[14] vssd1 vssd1 vccd1 vccd1 _07746_/A sky130_fd_sc_hd__dfxtp_1
X_07676_ _07676_/A _07699_/Y vssd1 vssd1 vccd1 vccd1 _13836_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_197_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09415_ _09445_/CLK line[0] vssd1 vssd1 vccd1 vccd1 _09416_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[14\].VALID\[14\].FF_D A[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12709__D line[107] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06627_ _06645_/CLK line[15] vssd1 vssd1 vccd1 vccd1 _06628_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10079__A _13922_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11613__D line[104] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08194__D line[91] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09346_ _09346_/A _09379_/Y vssd1 vssd1 vccd1 vccd1 _13826_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09868__A _13921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06707__D line[37] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06558_ _06558_/A _06579_/Y vssd1 vssd1 vccd1 vccd1 _13838_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_21_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05509_ _05525_/CLK line[1] vssd1 vssd1 vccd1 vccd1 _05510_/A sky130_fd_sc_hd__dfxtp_1
X_06489_ _06505_/CLK line[65] vssd1 vssd1 vccd1 vccd1 _06490_/A sky130_fd_sc_hd__dfxtp_1
X_09277_ _09305_/CLK line[74] vssd1 vssd1 vccd1 vccd1 _09278_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_138_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08228_ _08228_/A _08259_/Y vssd1 vssd1 vccd1 vccd1 _13828_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_193_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_OVHB\[27\].VALID\[2\].FF_D A[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08159_ _08185_/CLK line[75] vssd1 vssd1 vccd1 vccd1 _08160_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_162_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XDATA\[28\].CLKBUF\[1\] clk vssd1 vssd1 vccd1 vccd1 _10602_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__06442__D line[58] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11170_ _11170_/A _11199_/Y vssd1 vssd1 vccd1 vccd1 _13690_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[24\].VALID\[13\].FF_D A[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10121_ _10145_/CLK line[76] vssd1 vssd1 vccd1 vccd1 _10122_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[18\].CLKBUF\[7\] clk vssd1 vssd1 vccd1 vccd1 _07732_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__05058__D line[51] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10052_ _10052_/A _10079_/Y vssd1 vssd1 vccd1 vccd1 _13692_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10899__D line[33] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13275__D line[110] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08369__D line[43] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07273__D line[40] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13811_ _13811_/A _13824_/Y vssd1 vssd1 vccd1 vccd1 _13811_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[7\].VALID\[3\].FF OVHB\[7\].V/CLK A[10] vssd1 vssd1 vccd1 vccd1 OVHB\[7\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_44_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11373__A _13933_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13742_ _13750_/CLK line[53] vssd1 vssd1 vccd1 vccd1 _13743_/A sky130_fd_sc_hd__dfxtp_1
X_10954_ _13925_/X vssd1 vssd1 vccd1 vccd1 _10954_/Y sky130_fd_sc_hd__inv_2
X_13673_ _13673_/A _13684_/Y vssd1 vssd1 vccd1 vccd1 _13673_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11523__D line[77] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10885_ _10915_/CLK line[32] vssd1 vssd1 vccd1 vccd1 _10886_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06617__D line[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12624_ _12630_/CLK line[54] vssd1 vssd1 vccd1 vccd1 _12625_/A sky130_fd_sc_hd__dfxtp_1
XPHY_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05521__D line[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10139__D line[70] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12555_ _12555_/A _12564_/Y vssd1 vssd1 vccd1 vccd1 _13675_/Z sky130_fd_sc_hd__ebufn_2
XPHY_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11506_ _11510_/CLK line[55] vssd1 vssd1 vccd1 vccd1 _11507_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08832__D line[127] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12486_ _12490_/CLK line[119] vssd1 vssd1 vccd1 vccd1 _12487_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_184_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11437_ _11437_/A _11444_/Y vssd1 vssd1 vccd1 vccd1 _13677_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07448__D line[120] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11368_ _11370_/CLK line[120] vssd1 vssd1 vccd1 vccd1 _11369_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[26\].VALID\[14\].TOBUF OVHB\[26\].VALID\[14\].FF/Q OVHB\[26\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_98_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13107_ _13107_/A _13124_/Y vssd1 vssd1 vccd1 vccd1 _13667_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11548__A _13926_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10319_ _10319_/A _10324_/Y vssd1 vssd1 vccd1 vccd1 _13679_/Z sky130_fd_sc_hd__ebufn_2
X_11299_ _11299_/A _11304_/Y vssd1 vssd1 vccd1 vccd1 _13819_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[16\].VALID\[10\].FF_D A[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13038_ _13050_/CLK line[115] vssd1 vssd1 vccd1 vccd1 _13039_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_66_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05860_ _05860_/A _05879_/Y vssd1 vssd1 vccd1 vccd1 _13700_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07183__D line[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDATA\[17\].CLKBUF\[4\] clk vssd1 vssd1 vccd1 vccd1 _07347_/CLK sky130_fd_sc_hd__clkbuf_4
X_05791_ _05805_/CLK line[2] vssd1 vssd1 vccd1 vccd1 _05792_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_81_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07530_ _07530_/A _07559_/Y vssd1 vssd1 vccd1 vccd1 _13690_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_19_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07461_ _07485_/CLK line[12] vssd1 vssd1 vccd1 vccd1 _07462_/A sky130_fd_sc_hd__dfxtp_1
X_09200_ _09200_/CLK line[25] vssd1 vssd1 vccd1 vccd1 _09201_/A sky130_fd_sc_hd__dfxtp_1
X_06412_ _06412_/A _06439_/Y vssd1 vssd1 vccd1 vccd1 _13692_/Z sky130_fd_sc_hd__ebufn_2
X_07392_ _07392_/A _07419_/Y vssd1 vssd1 vccd1 vccd1 _13832_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_50_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05431__D line[108] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[6\].VALID\[6\].TOBUF OVHB\[6\].VALID\[6\].FF/Q OVHB\[6\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04923_/A2 sky130_fd_sc_hd__ebufn_2
XOVHB\[5\].VALID\[5\].FF OVHB\[5\].V/CLK A[12] vssd1 vssd1 vccd1 vccd1 OVHB\[5\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_06343_ _06365_/CLK line[13] vssd1 vssd1 vccd1 vccd1 _06344_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10049__D line[43] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09131_ _09131_/A _09134_/Y vssd1 vssd1 vccd1 vccd1 _13891_/Z sky130_fd_sc_hd__ebufn_2
X_09062_ _09062_/CLK _09063_/X vssd1 vssd1 vccd1 vccd1 _09060_/CLK sky130_fd_sc_hd__dlclkp_1
X_06274_ _06274_/A _06299_/Y vssd1 vssd1 vccd1 vccd1 _13834_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_175_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05225_ _05245_/CLK line[14] vssd1 vssd1 vccd1 vccd1 _05226_/A sky130_fd_sc_hd__dfxtp_1
X_08013_ _13912_/X wr vssd1 vssd1 vccd1 vccd1 _08013_/X sky130_fd_sc_hd__and2_1
XANTENNA__12264__D line[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07358__D line[93] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05156_ _05156_/A _05179_/Y vssd1 vssd1 vccd1 vccd1 _13836_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_131_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_OVHB\[29\].CG_CLK clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09964_ _09970_/CLK line[118] vssd1 vssd1 vccd1 vccd1 _09965_/A sky130_fd_sc_hd__dfxtp_1
X_05087_ _05105_/CLK line[79] vssd1 vssd1 vccd1 vccd1 _05088_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_103_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09573__D line[67] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08915_ _08915_/A _08924_/Y vssd1 vssd1 vccd1 vccd1 _13675_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_131_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09895_ _09895_/A _09904_/Y vssd1 vssd1 vccd1 vccd1 _13815_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_134_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10512__D line[127] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08846_ _08850_/CLK line[119] vssd1 vssd1 vccd1 vccd1 _08847_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05606__D line[60] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08777_ _08777_/A _08784_/Y vssd1 vssd1 vccd1 vccd1 _13817_/Z sky130_fd_sc_hd__ebufn_2
X_05989_ _06015_/CLK line[107] vssd1 vssd1 vccd1 vccd1 _05990_/A sky130_fd_sc_hd__dfxtp_1
X_07728_ _07730_/CLK line[120] vssd1 vssd1 vccd1 vccd1 _07729_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07821__D line[34] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12439__D line[97] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDATA\[16\].CLKBUF\[1\] clk vssd1 vssd1 vccd1 vccd1 _06962_/CLK sky130_fd_sc_hd__clkbuf_4
X_07659_ _07659_/A _07664_/Y vssd1 vssd1 vccd1 vccd1 _13819_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_80_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10670_ _10670_/CLK line[57] vssd1 vssd1 vccd1 vccd1 _10671_/A sky130_fd_sc_hd__dfxtp_1
XMUX.M\[2\].MUX\[1\] _13665_/Z _13735_/Z _13805_/Z _13875_/Z MUX.SEL0BUF\[2\]/X MUX.SEL1BUF\[2\]/X
+ vssd1 vssd1 vccd1 vccd1 Do[17] sky130_fd_sc_hd__mux4_1
X_09329_ _09329_/A _09344_/Y vssd1 vssd1 vccd1 vccd1 _13809_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_159_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09748__D line[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12340_ _12350_/CLK line[52] vssd1 vssd1 vccd1 vccd1 _12341_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_154_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[10\].VALID\[5\].FF_D A[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12271_ _12271_/A _12284_/Y vssd1 vssd1 vccd1 vccd1 _13671_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[13\].VALID\[10\].FF OVHB\[13\].V/CLK A[17] vssd1 vssd1 vccd1 vccd1 OVHB\[13\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11222_ _11230_/CLK line[53] vssd1 vssd1 vccd1 vccd1 _11223_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06172__D line[63] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[3\].VALID\[7\].FF OVHB\[3\].V/CLK A[14] vssd1 vssd1 vccd1 vccd1 OVHB\[3\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XOVHB\[13\].VALID\[1\].TOBUF OVHB\[13\].VALID\[1\].FF/Q OVHB\[13\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04926_/B2 sky130_fd_sc_hd__ebufn_2
X_11153_ _11153_/A _11164_/Y vssd1 vssd1 vccd1 vccd1 _13673_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12902__D line[53] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10104_ _10110_/CLK line[54] vssd1 vssd1 vccd1 vccd1 _10105_/A sky130_fd_sc_hd__dfxtp_1
X_11084_ _11090_/CLK line[118] vssd1 vssd1 vccd1 vccd1 _11085_/A sky130_fd_sc_hd__dfxtp_1
X_10035_ _10035_/A _10044_/Y vssd1 vssd1 vccd1 vccd1 _13675_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_103_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08099__D line[33] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_DATA\[18\].CLKBUF\[3\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11986_ _12000_/CLK line[18] vssd1 vssd1 vccd1 vccd1 _11987_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_63_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13725_ _13725_/A _13754_/Y vssd1 vssd1 vccd1 vccd1 _13725_/Z sky130_fd_sc_hd__ebufn_2
X_10937_ _10937_/A _10954_/Y vssd1 vssd1 vccd1 vccd1 _13737_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11253__D line[67] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06347__D line[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13656_ _13680_/CLK line[28] vssd1 vssd1 vccd1 vccd1 _13657_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_189_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10868_ _10880_/CLK line[19] vssd1 vssd1 vccd1 vccd1 _10869_/A sky130_fd_sc_hd__dfxtp_1
X_12607_ _12607_/A _12634_/Y vssd1 vssd1 vccd1 vccd1 _13727_/Z sky130_fd_sc_hd__ebufn_2
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13587_ _13587_/A _13614_/Y vssd1 vssd1 vccd1 vccd1 _13867_/Z sky130_fd_sc_hd__ebufn_2
X_10799_ _10799_/A _10814_/Y vssd1 vssd1 vccd1 vccd1 _13879_/Z sky130_fd_sc_hd__ebufn_2
XPHY_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08562__D line[117] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12538_ _12560_/CLK line[29] vssd1 vssd1 vccd1 vccd1 _12539_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_145_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12469_ _12469_/A _12494_/Y vssd1 vssd1 vccd1 vccd1 _13869_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[29\].V OVHB\[29\].V/CLK TIE/HI rst_n vssd1 vssd1 vccd1 vccd1 OVHB\[29\].V/Q
+ sky130_fd_sc_hd__dfrtp_1
XOVHB\[31\].VALID\[1\].FF OVHB\[31\].V/CLK A[8] vssd1 vssd1 vccd1 vccd1 OVHB\[31\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_05010_ _05010_/A _05039_/Y vssd1 vssd1 vccd1 vccd1 _13690_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_113_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12812__D line[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06810__D line[84] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06961_ _06961_/A _06964_/Y vssd1 vssd1 vccd1 vccd1 _13681_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_86_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XMUX.M\[1\].MUX\[3\] _13620_/Z _13690_/Z _13760_/Z _13830_/Z MUX.SEL0BUF\[1\]/X MUX.SEL1BUF\[1\]/X
+ vssd1 vssd1 vccd1 vccd1 Do[11] sky130_fd_sc_hd__mux4_1
XANTENNA__11428__D line[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08700_ _08710_/CLK line[52] vssd1 vssd1 vccd1 vccd1 _08701_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_100_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05912_ _05912_/CLK _05913_/X vssd1 vssd1 vccd1 vccd1 _05910_/CLK sky130_fd_sc_hd__dlclkp_1
X_09680_ _09690_/CLK line[116] vssd1 vssd1 vccd1 vccd1 _09681_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[16\].VOBUF OVHB\[16\].V/Q OVHB\[16\].INV/Y vssd1 vssd1 vccd1 vccd1 _04912_/B1
+ sky130_fd_sc_hd__ebufn_2
X_06892_ _06892_/CLK _06893_/X vssd1 vssd1 vccd1 vccd1 _06890_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_39_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XOVHB\[1\].VALID\[9\].FF OVHB\[1\].V/CLK A[16] vssd1 vssd1 vccd1 vccd1 OVHB\[1\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_08631_ _08631_/A _08644_/Y vssd1 vssd1 vccd1 vccd1 _13671_/Z sky130_fd_sc_hd__ebufn_2
X_05843_ _13902_/X wr vssd1 vssd1 vccd1 vccd1 _05843_/X sky130_fd_sc_hd__and2_1
XFILLER_54_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13643__D line[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[30\].VALID\[1\].FF_D A[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08737__D line[69] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08562_ _08570_/CLK line[117] vssd1 vssd1 vccd1 vccd1 _08563_/A sky130_fd_sc_hd__dfxtp_1
X_05774_ _13901_/X vssd1 vssd1 vccd1 vccd1 _05774_/Y sky130_fd_sc_hd__inv_2
X_07513_ _07513_/A _07524_/Y vssd1 vssd1 vccd1 vccd1 _13673_/Z sky130_fd_sc_hd__ebufn_2
X_08493_ _08493_/A _08504_/Y vssd1 vssd1 vccd1 vccd1 _13813_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07444_ _07450_/CLK line[118] vssd1 vssd1 vccd1 vccd1 _07445_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05161__D line[98] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07375_ _07375_/A _07384_/Y vssd1 vssd1 vccd1 vccd1 _13815_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[23\].VALID\[5\].FF_D A[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09114_ _09130_/CLK line[113] vssd1 vssd1 vccd1 vccd1 _09115_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08472__D line[90] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06326_ _06330_/CLK line[119] vssd1 vssd1 vccd1 vccd1 _06327_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_175_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09045_ _09045_/A _09064_/Y vssd1 vssd1 vccd1 vccd1 _13805_/Z sky130_fd_sc_hd__ebufn_2
X_06257_ _06257_/A _06264_/Y vssd1 vssd1 vccd1 vccd1 _13817_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07088__D line[83] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05208_ _05210_/CLK line[120] vssd1 vssd1 vccd1 vccd1 _05209_/A sky130_fd_sc_hd__dfxtp_1
X_06188_ _06190_/CLK line[56] vssd1 vssd1 vccd1 vccd1 _06189_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_89_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_OVHB\[16\].VALID\[9\].FF_D A[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13818__D line[88] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05139_ _05139_/A _05144_/Y vssd1 vssd1 vccd1 vccd1 _13819_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_1_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XOVHB\[8\].VALID\[12\].FF OVHB\[8\].V/CLK A[19] vssd1 vssd1 vccd1 vccd1 OVHB\[8\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_145_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06720__D line[48] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09947_ _09947_/A _09974_/Y vssd1 vssd1 vccd1 vccd1 _13867_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.M\[1\].MUX\[6\]_A2 _13766_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10242__D line[117] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09878_ _09900_/CLK line[93] vssd1 vssd1 vccd1 vccd1 _09879_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05336__D line[50] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05914__A _13902_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08829_ _08829_/A _08854_/Y vssd1 vssd1 vccd1 vccd1 _13869_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13553__D line[109] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11840_ _11860_/CLK line[94] vssd1 vssd1 vccd1 vccd1 _11841_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05633__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08647__D line[42] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_199_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07551__D line[39] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12169__D line[102] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11771_ _11771_/A _11794_/Y vssd1 vssd1 vccd1 vccd1 _13731_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_202_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[11\].VALID\[6\].TOBUF OVHB\[11\].VALID\[6\].FF/Q OVHB\[11\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04923_/A2 sky130_fd_sc_hd__ebufn_2
X_13510_ _13540_/CLK line[80] vssd1 vssd1 vccd1 vccd1 _13511_/A sky130_fd_sc_hd__dfxtp_1
X_10722_ _10740_/CLK line[95] vssd1 vssd1 vccd1 vccd1 _10723_/A sky130_fd_sc_hd__dfxtp_1
XMUX.M\[0\].MUX\[5\] _13638_/Z _13708_/Z _13778_/Z _13848_/Z MUX.SEL0BUF\[0\]/X MUX.SEL1BUF\[0\]/X
+ vssd1 vssd1 vccd1 vccd1 Do[5] sky130_fd_sc_hd__mux4_1
X_13441_ _13441_/A _13474_/Y vssd1 vssd1 vccd1 vccd1 _13721_/Z sky130_fd_sc_hd__ebufn_2
X_10653_ _10653_/A _10674_/Y vssd1 vssd1 vccd1 vccd1 _13733_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09478__D line[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11801__D line[76] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13372_ _13400_/CLK line[26] vssd1 vssd1 vccd1 vccd1 _13373_/A sky130_fd_sc_hd__dfxtp_1
X_10584_ _10600_/CLK line[17] vssd1 vssd1 vccd1 vccd1 _10585_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_70_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13578__A _13898_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12323_ _12323_/A _12354_/Y vssd1 vssd1 vccd1 vccd1 _13723_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10417__D line[69] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12254_ _12280_/CLK line[27] vssd1 vssd1 vccd1 vccd1 _12255_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_142_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13728__D line[61] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11205_ _11205_/A _11234_/Y vssd1 vssd1 vccd1 vccd1 _13725_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05808__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12185_ _12185_/A _12214_/Y vssd1 vssd1 vccd1 vccd1 _13865_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07726__D line[119] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[28\].VALID\[4\].FF OVHB\[28\].V/CLK A[11] vssd1 vssd1 vccd1 vccd1 OVHB\[28\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_11136_ _11160_/CLK line[28] vssd1 vssd1 vccd1 vccd1 _11137_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_150_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[4\].VALID\[0\].FF_D A[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10152__D line[90] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11067_ _11067_/A _11094_/Y vssd1 vssd1 vccd1 vccd1 _13867_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_95_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10018_ _10040_/CLK line[29] vssd1 vssd1 vccd1 vccd1 _10019_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_209_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[10\].VALID\[1\].FF OVHB\[10\].V/CLK A[8] vssd1 vssd1 vccd1 vccd1 OVHB\[10\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07461__D line[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12079__D line[75] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11969_ _13934_/X vssd1 vssd1 vccd1 vccd1 _11969_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06077__D line[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13708_ _13708_/A _13719_/Y vssd1 vssd1 vccd1 vccd1 _13708_/Z sky130_fd_sc_hd__ebufn_2
X_05490_ _05490_/CLK line[121] vssd1 vssd1 vccd1 vccd1 _05491_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_32_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13639_ _13645_/CLK line[6] vssd1 vssd1 vccd1 vccd1 _13640_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[16\].CLKBUF\[5\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09388__D line[125] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07160_ _07170_/CLK line[116] vssd1 vssd1 vccd1 vccd1 _07161_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_157_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06111_ _06111_/A _06124_/Y vssd1 vssd1 vccd1 vccd1 _13671_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_157_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07091_ _07091_/A _07104_/Y vssd1 vssd1 vccd1 vccd1 _13811_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10327__D line[42] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[29\].VALID\[9\].FF_D A[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06042_ _06050_/CLK line[117] vssd1 vssd1 vccd1 vccd1 _06043_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[16\].VALID\[12\].TOBUF OVHB\[16\].VALID\[12\].FF/Q OVHB\[16\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04929_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__12542__D line[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07636__D line[92] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09801_ _09801_/A _09834_/Y vssd1 vssd1 vccd1 vccd1 _13721_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06540__D line[89] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07993_ _07993_/A _08014_/Y vssd1 vssd1 vccd1 vccd1 _13873_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11158__D line[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09732_ _09760_/CLK line[26] vssd1 vssd1 vccd1 vccd1 _09733_/A sky130_fd_sc_hd__dfxtp_1
X_06944_ _06960_/CLK line[17] vssd1 vssd1 vccd1 vccd1 _06945_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_67_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09851__D line[66] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[9\].CLKBUF\[5\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09663_ _09663_/A _09694_/Y vssd1 vssd1 vccd1 vccd1 _13863_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_27_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06875_ _06875_/A _06894_/Y vssd1 vssd1 vccd1 vccd1 _13875_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_55_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08614_ _08640_/CLK line[27] vssd1 vssd1 vccd1 vccd1 _08615_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_131_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13951__A A_h[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05826_ _05840_/CLK line[18] vssd1 vssd1 vccd1 vccd1 _05827_/A sky130_fd_sc_hd__dfxtp_1
X_09594_ _09620_/CLK line[91] vssd1 vssd1 vccd1 vccd1 _09595_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_43_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XOVHB\[26\].VALID\[6\].FF OVHB\[26\].V/CLK A[13] vssd1 vssd1 vccd1 vccd1 OVHB\[26\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08545_ _08545_/A _08574_/Y vssd1 vssd1 vccd1 vccd1 _13865_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05757_ _05757_/A _05774_/Y vssd1 vssd1 vccd1 vccd1 _13877_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08476_ _08500_/CLK line[92] vssd1 vssd1 vccd1 vccd1 _08477_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05688_ _05700_/CLK line[83] vssd1 vssd1 vccd1 vccd1 _05689_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12717__D line[111] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07427_ _07427_/A _07454_/Y vssd1 vssd1 vccd1 vccd1 _13867_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_211_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06715__D line[41] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07358_ _07380_/CLK line[93] vssd1 vssd1 vccd1 vccd1 _07359_/A sky130_fd_sc_hd__dfxtp_1
X_06309_ _06309_/A _06334_/Y vssd1 vssd1 vccd1 vccd1 _13869_/Z sky130_fd_sc_hd__ebufn_2
X_07289_ _07289_/A _07314_/Y vssd1 vssd1 vccd1 vccd1 _13729_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_191_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09028_ _13915_/X wr vssd1 vssd1 vccd1 vccd1 _09028_/X sky130_fd_sc_hd__and2_1
XFILLER_151_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06450__D line[62] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11068__D line[125] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05066__D line[55] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12941_ _12945_/CLK line[71] vssd1 vssd1 vccd1 vccd1 _12942_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_18_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13283__D line[99] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MUX.M\[0\].MUX\[7\]_A0 _13642_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08377__D line[47] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12872_ _12872_/A _12879_/Y vssd1 vssd1 vccd1 vccd1 _13712_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[7\].CLKBUF\[5\] clk vssd1 vssd1 vccd1 vccd1 _13262_/CLK sky130_fd_sc_hd__clkbuf_4
X_11823_ _11825_/CLK line[72] vssd1 vssd1 vccd1 vccd1 _11824_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_60_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XOVHB\[26\].VALID\[0\].TOBUF OVHB\[26\].VALID\[0\].FF/Q OVHB\[26\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04924_/B2 sky130_fd_sc_hd__ebufn_2
X_11754_ _11754_/A _11759_/Y vssd1 vssd1 vccd1 vccd1 _13714_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10705_ _10705_/CLK line[73] vssd1 vssd1 vccd1 vccd1 _10706_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11685_ _11685_/CLK line[9] vssd1 vssd1 vccd1 vccd1 _11686_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11531__D line[66] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[24\].VALID\[8\].FF OVHB\[24\].V/CLK A[15] vssd1 vssd1 vccd1 vccd1 OVHB\[24\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_13424_ _13424_/A _13439_/Y vssd1 vssd1 vccd1 vccd1 _13704_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06625__D line[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10636_ _10636_/A _10639_/Y vssd1 vssd1 vccd1 vccd1 _13716_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[4\].VALID\[10\].FF OVHB\[4\].V/CLK A[17] vssd1 vssd1 vccd1 vccd1 OVHB\[4\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__09001__D line[76] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13355_ _13365_/CLK line[4] vssd1 vssd1 vccd1 vccd1 _13356_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_139_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10567_ _10567_/CLK _10568_/X vssd1 vssd1 vccd1 vccd1 _10565_/CLK sky130_fd_sc_hd__dlclkp_1
X_12306_ _12306_/A _12319_/Y vssd1 vssd1 vccd1 vccd1 _13706_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08840__D line[116] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13286_ _13286_/A _13299_/Y vssd1 vssd1 vccd1 vccd1 _13846_/Z sky130_fd_sc_hd__ebufn_2
X_10498_ _13923_/X wr vssd1 vssd1 vccd1 vccd1 _10498_/X sky130_fd_sc_hd__and2_1
XANTENNA__13458__D line[51] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12237_ _12245_/CLK line[5] vssd1 vssd1 vccd1 vccd1 _12238_/A sky130_fd_sc_hd__dfxtp_1
X_12168_ _12168_/A _12179_/Y vssd1 vssd1 vccd1 vccd1 _13848_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_110_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11119_ _11125_/CLK line[6] vssd1 vssd1 vccd1 vccd1 _11120_/A sky130_fd_sc_hd__dfxtp_1
X_04990_ _05000_/CLK line[20] vssd1 vssd1 vccd1 vccd1 _04991_/A sky130_fd_sc_hd__dfxtp_1
X_12099_ _12105_/CLK line[70] vssd1 vssd1 vccd1 vccd1 _12100_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[24\].CGAND _13920_/Y wr vssd1 vssd1 vccd1 vccd1 OVHB\[24\].CGAND/X sky130_fd_sc_hd__and2_4
XFILLER_77_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11706__D line[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06660_ _06680_/CLK line[30] vssd1 vssd1 vccd1 vccd1 _06661_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07191__D line[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05611_ _05611_/A _05634_/Y vssd1 vssd1 vccd1 vccd1 _13731_/Z sky130_fd_sc_hd__ebufn_2
X_06591_ _06591_/A _06614_/Y vssd1 vssd1 vccd1 vccd1 _13871_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_91_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08330_ _08360_/CLK line[16] vssd1 vssd1 vccd1 vccd1 _08331_/A sky130_fd_sc_hd__dfxtp_1
X_05542_ _05560_/CLK line[31] vssd1 vssd1 vccd1 vccd1 _05543_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[6\].CLKBUF\[2\] clk vssd1 vssd1 vccd1 vccd1 _12877_/CLK sky130_fd_sc_hd__clkbuf_4
X_05473_ _05473_/A _05494_/Y vssd1 vssd1 vccd1 vccd1 _13873_/Z sky130_fd_sc_hd__ebufn_2
X_08261_ _08261_/A _08294_/Y vssd1 vssd1 vccd1 vccd1 _13861_/Z sky130_fd_sc_hd__ebufn_2
X_07212_ _07240_/CLK line[26] vssd1 vssd1 vccd1 vccd1 _07213_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[18\].VALID\[6\].TOBUF OVHB\[18\].VALID\[6\].FF/Q OVHB\[18\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04923_/A2 sky130_fd_sc_hd__ebufn_2
X_08192_ _08220_/CLK line[90] vssd1 vssd1 vccd1 vccd1 _08193_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_118_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07143_ _07143_/A _07174_/Y vssd1 vssd1 vccd1 vccd1 _13863_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10057__D line[47] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07074_ _07100_/CLK line[91] vssd1 vssd1 vccd1 vccd1 _07075_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_118_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08750__D line[80] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_DATA\[14\].CLKBUF\[7\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12272__D line[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06025_ _06025_/A _06054_/Y vssd1 vssd1 vccd1 vccd1 _13865_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_160_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07366__D line[82] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07944__A _13912_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[1\].VALID\[13\].FF_D A[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07663__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07976_ _07976_/A _07979_/Y vssd1 vssd1 vccd1 vccd1 _13856_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_75_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09581__D line[71] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09715_ _09725_/CLK line[4] vssd1 vssd1 vccd1 vccd1 _09716_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_19_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06927_ _06927_/CLK _06928_/X vssd1 vssd1 vccd1 vccd1 _06925_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_142_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10520__D line[116] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09646_ _09646_/A _09659_/Y vssd1 vssd1 vccd1 vccd1 _13846_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[26\].CLKBUF\[6\] clk vssd1 vssd1 vccd1 vccd1 _10217_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_28_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06858_ _13905_/X wr vssd1 vssd1 vccd1 vccd1 _06858_/X sky130_fd_sc_hd__and2_1
XFILLER_43_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05614__D line[49] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05809_ _13902_/X vssd1 vssd1 vccd1 vccd1 _05809_/Y sky130_fd_sc_hd__inv_2
X_09577_ _09585_/CLK line[69] vssd1 vssd1 vccd1 vccd1 _09578_/A sky130_fd_sc_hd__dfxtp_1
X_06789_ _13905_/X vssd1 vssd1 vccd1 vccd1 _06789_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13831__D line[108] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08528_ _08528_/A _08539_/Y vssd1 vssd1 vccd1 vccd1 _13848_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[7\].CLKBUF\[7\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08925__D line[32] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[18\].VALID\[10\].FF OVHB\[18\].V/CLK A[17] vssd1 vssd1 vccd1 vccd1 OVHB\[18\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12447__D line[101] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08459_ _08465_/CLK line[70] vssd1 vssd1 vccd1 vccd1 _08460_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11470_ _11470_/A _11479_/Y vssd1 vssd1 vccd1 vccd1 _13710_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10421_ _10425_/CLK line[71] vssd1 vssd1 vccd1 vccd1 _10422_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_167_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07838__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09756__D line[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13140_ _13140_/A _13159_/Y vssd1 vssd1 vccd1 vccd1 _13700_/Z sky130_fd_sc_hd__ebufn_2
X_10352_ _10352_/A _10359_/Y vssd1 vssd1 vccd1 vccd1 _13712_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12182__D line[122] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[0\].VALID\[3\].FF_D A[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13071_ _13085_/CLK line[2] vssd1 vssd1 vccd1 vccd1 _13072_/A sky130_fd_sc_hd__dfxtp_1
X_10283_ _10285_/CLK line[8] vssd1 vssd1 vccd1 vccd1 _10284_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_151_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06180__D line[52] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12022_ _12022_/A _12039_/Y vssd1 vssd1 vccd1 vccd1 _13702_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[24\].VALID\[5\].TOBUF OVHB\[24\].VALID\[5\].FF/Q OVHB\[24\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04927_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_104_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12910__D line[57] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09491__D line[44] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13973_ A_h[1] vssd1 vssd1 vccd1 vccd1 _13982_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_18_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10430__D line[80] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12924_ _12924_/A _12949_/Y vssd1 vssd1 vccd1 vccd1 _13764_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_19_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12855_ _12875_/CLK line[46] vssd1 vssd1 vccd1 vccd1 _12856_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_73_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[10\].CGAND_B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11806_ _11806_/A _11829_/Y vssd1 vssd1 vccd1 vccd1 _13766_/Z sky130_fd_sc_hd__ebufn_2
X_12786_ _12786_/A _12809_/Y vssd1 vssd1 vccd1 vccd1 _13626_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_92_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XDATA\[25\].CLKBUF\[3\] clk vssd1 vssd1 vccd1 vccd1 _09832_/CLK sky130_fd_sc_hd__clkbuf_4
XPHY_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12357__D line[74] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11737_ _11755_/CLK line[47] vssd1 vssd1 vccd1 vccd1 _11738_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_159_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11261__D line[71] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_OVHB\[14\].CGAND_A _13904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06355__D line[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11668_ _11668_/A _11689_/Y vssd1 vssd1 vccd1 vccd1 _13628_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_174_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13407_ _13435_/CLK line[42] vssd1 vssd1 vccd1 vccd1 _13408_/A sky130_fd_sc_hd__dfxtp_1
X_10619_ _10635_/CLK line[33] vssd1 vssd1 vccd1 vccd1 _10620_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11599_ _11615_/CLK line[97] vssd1 vssd1 vccd1 vccd1 _11600_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09666__D line[124] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13338_ _13338_/A _13369_/Y vssd1 vssd1 vccd1 vccd1 _13618_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08570__D line[121] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13188__D line[56] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10605__D line[32] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13269_ _13295_/CLK line[107] vssd1 vssd1 vccd1 vccd1 _13270_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06090__D line[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12820__D line[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07830_ _07830_/A _07839_/Y vssd1 vssd1 vccd1 vccd1 _13710_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_110_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07914__D line[91] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05284__A _13900_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07761_ _07765_/CLK line[7] vssd1 vssd1 vccd1 vccd1 _07762_/A sky130_fd_sc_hd__dfxtp_1
X_04973_ _04973_/A _05004_/Y vssd1 vssd1 vccd1 vccd1 _13653_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11436__D line[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09500_ _09500_/A _09519_/Y vssd1 vssd1 vccd1 vccd1 _13700_/Z sky130_fd_sc_hd__ebufn_2
X_06712_ _06712_/A _06719_/Y vssd1 vssd1 vccd1 vccd1 _13712_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[15\].VALID\[0\].FF_D A[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07692_ _07692_/A _07699_/Y vssd1 vssd1 vccd1 vccd1 _13852_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_65_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09431_ _09445_/CLK line[2] vssd1 vssd1 vccd1 vccd1 _09432_/A sky130_fd_sc_hd__dfxtp_1
X_06643_ _06645_/CLK line[8] vssd1 vssd1 vccd1 vccd1 _06644_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[30\].VALID\[4\].TOBUF OVHB\[30\].VALID\[4\].FF/Q OVHB\[30\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04925_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_80_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09362_ _09362_/A _09379_/Y vssd1 vssd1 vccd1 vccd1 _13842_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09203__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08745__D line[73] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06574_ _06574_/A _06579_/Y vssd1 vssd1 vccd1 vccd1 _13854_/Z sky130_fd_sc_hd__ebufn_2
X_08313_ _08325_/CLK line[3] vssd1 vssd1 vccd1 vccd1 _08314_/A sky130_fd_sc_hd__dfxtp_1
X_05525_ _05525_/CLK line[9] vssd1 vssd1 vccd1 vccd1 _05526_/A sky130_fd_sc_hd__dfxtp_1
X_09293_ _09305_/CLK line[67] vssd1 vssd1 vccd1 vccd1 _09294_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11171__D line[44] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08244_ _08244_/A _08259_/Y vssd1 vssd1 vccd1 vccd1 _13844_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06265__D line[96] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05456_ _05456_/A _05459_/Y vssd1 vssd1 vccd1 vccd1 _13856_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_119_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08175_ _08185_/CLK line[68] vssd1 vssd1 vccd1 vccd1 _08176_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_193_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XDATA\[24\].CLKBUF\[0\] clk vssd1 vssd1 vccd1 vccd1 _09447_/CLK sky130_fd_sc_hd__clkbuf_4
X_05387_ _05387_/CLK _05388_/X vssd1 vssd1 vccd1 vccd1 _05385_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA_DATA\[28\].CLKBUF\[1\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07126_ _07126_/A _07139_/Y vssd1 vssd1 vccd1 vccd1 _13846_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08480__D line[94] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05459__A _13900_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13098__D line[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XDATA\[14\].CLKBUF\[6\] clk vssd1 vssd1 vccd1 vccd1 _06577_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__05178__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07057_ _07065_/CLK line[69] vssd1 vssd1 vccd1 vccd1 _07058_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_133_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07096__D line[87] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06008_ _06008_/A _06019_/Y vssd1 vssd1 vccd1 vccd1 _13848_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[6\].VALID\[7\].FF_D A[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07959_ _07975_/CLK line[97] vssd1 vssd1 vccd1 vccd1 _07960_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DEC.DEC0.AND1_A_N A[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11346__D line[124] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10250__D line[121] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[14\].CG clk OVHB\[14\].CGAND/X vssd1 vssd1 vccd1 vccd1 OVHB\[14\].V/CLK sky130_fd_sc_hd__dlclkp_1
X_10970_ _10970_/A _10989_/Y vssd1 vssd1 vccd1 vccd1 _13770_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05344__D line[54] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09629_ _09655_/CLK line[107] vssd1 vssd1 vccd1 vccd1 _09630_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_15_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13561__D line[98] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MUX.M\[0\].MUX\[4\]_A3 _13846_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12640_ _12640_/A _12669_/Y vssd1 vssd1 vccd1 vccd1 _13760_/Z sky130_fd_sc_hd__ebufn_2
XPHY_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08655__D line[46] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12571_ _12595_/CLK line[44] vssd1 vssd1 vccd1 vccd1 _12572_/A sky130_fd_sc_hd__dfxtp_1
XPHY_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11522_ _11522_/A _11549_/Y vssd1 vssd1 vccd1 vccd1 _13762_/Z sky130_fd_sc_hd__ebufn_2
XPHY_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06753__A _13905_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11453_ _11475_/CLK line[45] vssd1 vssd1 vccd1 vccd1 _11454_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_109_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XOVHB\[6\].VALID\[14\].TOBUF OVHB\[6\].VALID\[14\].FF/Q OVHB\[6\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/B2 sky130_fd_sc_hd__ebufn_2
X_10404_ _10404_/A _10429_/Y vssd1 vssd1 vccd1 vccd1 _13764_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06903__D line[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11384_ _11384_/A _11409_/Y vssd1 vssd1 vccd1 vccd1 _13624_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_164_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__04930__A1_N A_h[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13123_ _13938_/X wr vssd1 vssd1 vccd1 vccd1 _13123_/X sky130_fd_sc_hd__and2_1
XFILLER_194_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10425__D line[73] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10335_ _10355_/CLK line[46] vssd1 vssd1 vccd1 vccd1 _10336_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_124_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_DATA\[1\].CLKBUF\[0\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05519__D line[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13054_ _13937_/X vssd1 vssd1 vccd1 vccd1 _13054_/Y sky130_fd_sc_hd__inv_2
X_10266_ _10266_/A _10289_/Y vssd1 vssd1 vccd1 vccd1 _13626_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13736__D line[50] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12005_ _12035_/CLK line[32] vssd1 vssd1 vccd1 vccd1 _12006_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_87_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XDATA\[13\].CLKBUF\[3\] clk vssd1 vssd1 vccd1 vccd1 _06192_/CLK sky130_fd_sc_hd__clkbuf_4
X_10197_ _10215_/CLK line[111] vssd1 vssd1 vccd1 vccd1 _10198_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[28\].VALID\[0\].FF_D A[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10160__D line[94] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[8\].VALID\[13\].FF_D A[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05254__D line[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13956_ _13960_/C _13960_/B _13960_/A _13960_/D vssd1 vssd1 vccd1 vccd1 _13956_/X
+ sky130_fd_sc_hd__and4b_4
XANTENNA__06928__A _13909_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12907_ _12907_/A _12914_/Y vssd1 vssd1 vccd1 vccd1 _13747_/Z sky130_fd_sc_hd__ebufn_2
X_13887_ _13887_/A _13894_/Y vssd1 vssd1 vccd1 vccd1 _13887_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[26\].VALID\[10\].TOBUF OVHB\[26\].VALID\[10\].FF/Q OVHB\[26\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04932_/B2 sky130_fd_sc_hd__ebufn_2
X_12838_ _12840_/CLK line[24] vssd1 vssd1 vccd1 vccd1 _12839_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_210_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12087__D line[79] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12769_ _12769_/A _12774_/Y vssd1 vssd1 vccd1 vccd1 _13889_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06085__D line[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05310_ _05310_/A _05319_/Y vssd1 vssd1 vccd1 vccd1 _13710_/Z sky130_fd_sc_hd__ebufn_2
X_06290_ _06290_/A _06299_/Y vssd1 vssd1 vccd1 vccd1 _13850_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_175_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05241_ _05245_/CLK line[7] vssd1 vssd1 vccd1 vccd1 _05242_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_128_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09396__D line[114] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09974__A _13921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05172_ _05172_/A _05179_/Y vssd1 vssd1 vccd1 vccd1 _13852_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[19\].V_RESET_B rst_n vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10335__D line[46] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09693__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09980_ _09980_/A _10009_/Y vssd1 vssd1 vccd1 vccd1 _13620_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05429__D line[107] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08931_ _08955_/CLK line[44] vssd1 vssd1 vccd1 vccd1 _08932_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_143_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__04911__A A_h[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12550__D line[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[6\].VALID\[2\].TOBUF OVHB\[6\].VALID\[2\].FF/Q OVHB\[6\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04930_/B2 sky130_fd_sc_hd__ebufn_2
X_08862_ _08862_/A _08889_/Y vssd1 vssd1 vccd1 vccd1 _13622_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07644__D line[81] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07813_ _07835_/CLK line[45] vssd1 vssd1 vccd1 vccd1 _07814_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_29_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08793_ _08815_/CLK line[109] vssd1 vssd1 vccd1 vccd1 _08794_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_123_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07744_ _07744_/A _07769_/Y vssd1 vssd1 vccd1 vccd1 _13624_/Z sky130_fd_sc_hd__ebufn_2
X_04956_ _04956_/A _04969_/Y vssd1 vssd1 vccd1 vccd1 _13636_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_65_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XDATA\[12\].CLKBUF\[0\] clk vssd1 vssd1 vccd1 vccd1 _05807_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07675_ _07695_/CLK line[110] vssd1 vssd1 vccd1 vccd1 _07676_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[9\].CG clk OVHB\[9\].CGAND/X vssd1 vssd1 vccd1 vccd1 OVHB\[9\].V/CLK sky130_fd_sc_hd__dlclkp_1
X_09414_ _13916_/X vssd1 vssd1 vccd1 vccd1 _09414_/Y sky130_fd_sc_hd__inv_2
X_06626_ _06626_/A _06649_/Y vssd1 vssd1 vccd1 vccd1 _13626_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_80_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09345_ _09375_/CLK line[96] vssd1 vssd1 vccd1 vccd1 _09346_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09868__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06557_ _06575_/CLK line[111] vssd1 vssd1 vccd1 vccd1 _06558_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_166_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05508_ _05508_/A _05529_/Y vssd1 vssd1 vccd1 vccd1 _13628_/Z sky130_fd_sc_hd__ebufn_2
X_09276_ _09276_/A _09309_/Y vssd1 vssd1 vccd1 vccd1 _13756_/Z sky130_fd_sc_hd__ebufn_2
X_06488_ _06488_/A _06509_/Y vssd1 vssd1 vccd1 vccd1 _13768_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_21_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08227_ _08255_/CLK line[106] vssd1 vssd1 vccd1 vccd1 _08228_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12725__D line[100] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05439_ _05455_/CLK line[97] vssd1 vssd1 vccd1 vccd1 _05440_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07819__D line[33] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08158_ _08158_/A _08189_/Y vssd1 vssd1 vccd1 vccd1 _13758_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_146_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07109_ _07135_/CLK line[107] vssd1 vssd1 vccd1 vccd1 _07110_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_134_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08089_ _08115_/CLK line[43] vssd1 vssd1 vccd1 vccd1 _08090_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_106_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10120_ _10120_/A _10149_/Y vssd1 vssd1 vccd1 vccd1 _13760_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_0_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_DATA\[26\].CLKBUF\[3\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12460__D line[112] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10051_ _10075_/CLK line[44] vssd1 vssd1 vccd1 vccd1 _10052_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_196_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11076__D line[114] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11654__A _13926_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13810_ _13820_/CLK line[84] vssd1 vssd1 vccd1 vccd1 _13811_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_91_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13741_ _13741_/A _13754_/Y vssd1 vssd1 vccd1 vccd1 _13741_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_90_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11373__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10953_ _13925_/X wr vssd1 vssd1 vccd1 vccd1 _10953_/X sky130_fd_sc_hd__and2_1
XANTENNA__13291__D line[103] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[9\].VALID\[10\].FF OVHB\[9\].V/CLK A[17] vssd1 vssd1 vccd1 vccd1 OVHB\[9\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08385__D line[36] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13672_ _13680_/CLK line[21] vssd1 vssd1 vccd1 vccd1 _13673_/A sky130_fd_sc_hd__dfxtp_1
X_10884_ _13925_/X vssd1 vssd1 vccd1 vccd1 _10884_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12623_ _12623_/A _12634_/Y vssd1 vssd1 vccd1 vccd1 _13743_/Z sky130_fd_sc_hd__ebufn_2
XPHY_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12554_ _12560_/CLK line[22] vssd1 vssd1 vccd1 vccd1 _12555_/A sky130_fd_sc_hd__dfxtp_1
XPHY_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11505_ _11505_/A _11514_/Y vssd1 vssd1 vccd1 vccd1 _13745_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_157_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12635__D line[64] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12485_ _12485_/A _12494_/Y vssd1 vssd1 vccd1 vccd1 _13885_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06633__D line[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11436_ _11440_/CLK line[23] vssd1 vssd1 vccd1 vccd1 _11437_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_125_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11829__A _13927_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11367_ _11367_/A _11374_/Y vssd1 vssd1 vccd1 vccd1 _13887_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09944__D line[123] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13106_ _13120_/CLK line[18] vssd1 vssd1 vccd1 vccd1 _13107_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_3_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10318_ _10320_/CLK line[24] vssd1 vssd1 vccd1 vccd1 _10319_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11548__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11298_ _11300_/CLK line[88] vssd1 vssd1 vccd1 vccd1 _11299_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13466__D line[55] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13037_ _13037_/A _13054_/Y vssd1 vssd1 vccd1 vccd1 _13877_/Z sky130_fd_sc_hd__ebufn_2
X_10249_ _10249_/A _10254_/Y vssd1 vssd1 vccd1 vccd1 _13889_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_39_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_OVHB\[11\].VALID\[3\].FF_D A[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09031__TE_B _09064_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05790_ _05790_/A _05809_/Y vssd1 vssd1 vccd1 vccd1 _13630_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_207_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13939_ A_h[0] vssd1 vssd1 vccd1 vccd1 _13949_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__11714__D line[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08295__D line[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07460_ _07460_/A _07489_/Y vssd1 vssd1 vccd1 vccd1 _13620_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06808__D line[83] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06411_ _06435_/CLK line[44] vssd1 vssd1 vccd1 vccd1 _06412_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_50_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07391_ _07415_/CLK line[108] vssd1 vssd1 vccd1 vccd1 _07392_/A sky130_fd_sc_hd__dfxtp_1
X_09130_ _09130_/CLK line[121] vssd1 vssd1 vccd1 vccd1 _09131_/A sky130_fd_sc_hd__dfxtp_1
X_06342_ _06342_/A _06369_/Y vssd1 vssd1 vccd1 vccd1 _13622_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07489__A _13911_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XOVHB\[4\].VALID\[7\].TOBUF OVHB\[4\].VALID\[7\].FF/Q OVHB\[4\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/A2 sky130_fd_sc_hd__ebufn_2
XOVHB\[12\].VOBUF OVHB\[12\].V/Q OVHB\[12\].INV/Y vssd1 vssd1 vccd1 vccd1 _04912_/B1
+ sky130_fd_sc_hd__ebufn_2
X_09061_ _09061_/A _09064_/Y vssd1 vssd1 vccd1 vccd1 _13821_/Z sky130_fd_sc_hd__ebufn_2
X_06273_ _06295_/CLK line[109] vssd1 vssd1 vccd1 vccd1 _06274_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_147_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08012_ _08012_/CLK _08013_/X vssd1 vssd1 vccd1 vccd1 _08010_/CLK sky130_fd_sc_hd__dlclkp_1
X_05224_ _05224_/A _05249_/Y vssd1 vssd1 vccd1 vccd1 _13624_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_190_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10065__D line[36] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05155_ _05175_/CLK line[110] vssd1 vssd1 vccd1 vccd1 _05156_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05159__D line[97] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09963_ _09963_/A _09974_/Y vssd1 vssd1 vccd1 vccd1 _13883_/Z sky130_fd_sc_hd__ebufn_2
X_05086_ _05086_/A _05109_/Y vssd1 vssd1 vccd1 vccd1 _13766_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[10\].VALID\[11\].FF_D A[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13376__D line[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12280__D line[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08914_ _08920_/CLK line[22] vssd1 vssd1 vccd1 vccd1 _08915_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__04998__D line[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09894_ _09900_/CLK line[86] vssd1 vssd1 vccd1 vccd1 _09895_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07374__D line[86] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08845_ _08845_/A _08854_/Y vssd1 vssd1 vccd1 vccd1 _13885_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_85_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08776_ _08780_/CLK line[87] vssd1 vssd1 vccd1 vccd1 _08777_/A sky130_fd_sc_hd__dfxtp_1
X_05988_ _05988_/A _06019_/Y vssd1 vssd1 vccd1 vccd1 _13828_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_150_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07727_ _07727_/A _07734_/Y vssd1 vssd1 vccd1 vccd1 _13887_/Z sky130_fd_sc_hd__ebufn_2
X_04939_ _04965_/CLK line[11] vssd1 vssd1 vccd1 vccd1 _04940_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_53_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11624__D line[123] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07658_ _07660_/CLK line[88] vssd1 vssd1 vccd1 vccd1 _07659_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05622__D line[53] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08783__A _13914_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[20\].VALID\[10\].FF_D A[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06609_ _06609_/A _06614_/Y vssd1 vssd1 vccd1 vccd1 _13889_/Z sky130_fd_sc_hd__ebufn_2
X_07589_ _07589_/A _07594_/Y vssd1 vssd1 vccd1 vccd1 _13749_/Z sky130_fd_sc_hd__ebufn_2
X_09328_ _09340_/CLK line[83] vssd1 vssd1 vccd1 vccd1 _09329_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08933__D line[45] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[19\].VALID\[0\].FF OVHB\[19\].V/CLK A[7] vssd1 vssd1 vccd1 vccd1 OVHB\[19\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_09259_ _09259_/A _09274_/Y vssd1 vssd1 vccd1 vccd1 _13739_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12455__D line[105] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07549__D line[38] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12270_ _12280_/CLK line[20] vssd1 vssd1 vccd1 vccd1 _12271_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11221_ _11221_/A _11234_/Y vssd1 vssd1 vccd1 vccd1 _13741_/Z sky130_fd_sc_hd__ebufn_2
X_11152_ _11160_/CLK line[21] vssd1 vssd1 vccd1 vccd1 _11153_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[24\].VALID\[3\].FF_D A[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[11\].VALID\[2\].TOBUF OVHB\[11\].VALID\[2\].FF/Q OVHB\[11\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04930_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_0_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12190__D line[126] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10103_ _10103_/A _10114_/Y vssd1 vssd1 vccd1 vccd1 _13743_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10703__D line[72] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11083_ _11083_/A _11094_/Y vssd1 vssd1 vccd1 vccd1 _13883_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07284__D line[59] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08958__A _13915_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10034_ _10040_/CLK line[22] vssd1 vssd1 vccd1 vccd1 _10035_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_48_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_OVHB\[17\].VALID\[7\].FF_D A[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[24\].CLKBUF\[5\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11985_ _11985_/A _12004_/Y vssd1 vssd1 vccd1 vccd1 _13665_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_44_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13724_ _13750_/CLK line[59] vssd1 vssd1 vccd1 vccd1 _13725_/A sky130_fd_sc_hd__dfxtp_1
X_10936_ _10950_/CLK line[50] vssd1 vssd1 vccd1 vccd1 _10937_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_204_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05532__D line[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10867_ _10867_/A _10884_/Y vssd1 vssd1 vccd1 vccd1 _13667_/Z sky130_fd_sc_hd__ebufn_2
X_13655_ _13655_/A _13684_/Y vssd1 vssd1 vccd1 vccd1 _13655_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_32_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12606_ _12630_/CLK line[60] vssd1 vssd1 vccd1 vccd1 _12607_/A sky130_fd_sc_hd__dfxtp_1
X_13586_ _13610_/CLK line[124] vssd1 vssd1 vccd1 vccd1 _13587_/A sky130_fd_sc_hd__dfxtp_1
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10798_ _10810_/CLK line[115] vssd1 vssd1 vccd1 vccd1 _10799_/A sky130_fd_sc_hd__dfxtp_1
XPHY_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12537_ _12537_/A _12564_/Y vssd1 vssd1 vccd1 vccd1 _13657_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12365__D line[78] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07459__D line[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06363__D line[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12468_ _12490_/CLK line[125] vssd1 vssd1 vccd1 vccd1 _12469_/A sky130_fd_sc_hd__dfxtp_1
X_11419_ _11419_/A _11444_/Y vssd1 vssd1 vccd1 vccd1 _13659_/Z sky130_fd_sc_hd__ebufn_2
X_12399_ _12399_/A _12424_/Y vssd1 vssd1 vccd1 vccd1 _13799_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10463__A _13923_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09674__D line[113] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[19\].V_D TIE/HI vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09029__A _13915_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[17\].VALID\[2\].FF OVHB\[17\].V/CLK A[9] vssd1 vssd1 vccd1 vccd1 OVHB\[17\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XDATA\[4\].CLKBUF\[7\] clk vssd1 vssd1 vccd1 vccd1 _12492_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__10613__D line[45] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06960_ _06960_/CLK line[25] vssd1 vssd1 vccd1 vccd1 _06961_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_100_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05707__D line[106] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05911_ _05911_/A _05914_/Y vssd1 vssd1 vccd1 vccd1 _13751_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_39_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06891_ _06891_/A _06894_/Y vssd1 vssd1 vccd1 vccd1 _13891_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_67_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08630_ _08640_/CLK line[20] vssd1 vssd1 vccd1 vccd1 _08631_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_55_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05842_ _05842_/CLK _05843_/X vssd1 vssd1 vccd1 vccd1 _05840_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__07922__D line[95] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08561_ _08561_/A _08574_/Y vssd1 vssd1 vccd1 vccd1 _13881_/Z sky130_fd_sc_hd__ebufn_2
X_05773_ _13901_/X wr vssd1 vssd1 vccd1 vccd1 _05773_/X sky130_fd_sc_hd__and2_1
XFILLER_35_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07512_ _07520_/CLK line[21] vssd1 vssd1 vccd1 vccd1 _07513_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06538__D line[88] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08492_ _08500_/CLK line[85] vssd1 vssd1 vccd1 vccd1 _08493_/A sky130_fd_sc_hd__dfxtp_1
X_07443_ _07443_/A _07454_/Y vssd1 vssd1 vccd1 vccd1 _13883_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_168_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10638__A _13924_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09849__D line[65] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07374_ _07380_/CLK line[86] vssd1 vssd1 vccd1 vccd1 _07375_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_13_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09113_ _09113_/A _09134_/Y vssd1 vssd1 vccd1 vccd1 _13873_/Z sky130_fd_sc_hd__ebufn_2
X_06325_ _06325_/A _06334_/Y vssd1 vssd1 vccd1 vccd1 _13885_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[19\].CGAND _13912_/X wr vssd1 vssd1 vccd1 vccd1 OVHB\[19\].CGAND/X sky130_fd_sc_hd__and2_4
XFILLER_129_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09044_ _09060_/CLK line[81] vssd1 vssd1 vccd1 vccd1 _09045_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06273__D line[109] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06256_ _06260_/CLK line[87] vssd1 vssd1 vccd1 vccd1 _06257_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_190_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05207_ _05207_/A _05214_/Y vssd1 vssd1 vccd1 vccd1 _13887_/Z sky130_fd_sc_hd__ebufn_2
X_06187_ _06187_/A _06194_/Y vssd1 vssd1 vccd1 vccd1 _13747_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_104_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05138_ _05140_/CLK line[88] vssd1 vssd1 vccd1 vccd1 _05139_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_1_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13684__A _13899_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[25\].VALID\[14\].FF_D A[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09946_ _09970_/CLK line[124] vssd1 vssd1 vccd1 vccd1 _09947_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_77_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05069_ _05069_/A _05074_/Y vssd1 vssd1 vccd1 vccd1 _13749_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_58_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_MUX.M\[1\].MUX\[6\]_A3 _13836_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09877_ _09877_/A _09904_/Y vssd1 vssd1 vccd1 vccd1 _13797_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_97_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XDATA\[3\].CLKBUF\[4\] clk vssd1 vssd1 vccd1 vccd1 _12107_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_161_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08828_ _08850_/CLK line[125] vssd1 vssd1 vccd1 vccd1 _08829_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06298__A _13903_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[15\].VALID\[4\].FF OVHB\[15\].V/CLK A[11] vssd1 vssd1 vccd1 vccd1 OVHB\[15\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_08759_ _08759_/A _08784_/Y vssd1 vssd1 vccd1 vccd1 _13799_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11354__D line[113] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06448__D line[61] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11770_ _11790_/CLK line[62] vssd1 vssd1 vccd1 vccd1 _11771_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_53_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10721_ _10721_/A _10744_/Y vssd1 vssd1 vccd1 vccd1 _13801_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_54_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XOVHB\[31\].VALID\[13\].FF OVHB\[31\].V/CLK A[20] vssd1 vssd1 vccd1 vccd1 OVHB\[31\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_14_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13440_ _13470_/CLK line[48] vssd1 vssd1 vccd1 vccd1 _13441_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08663__D line[35] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10652_ _10670_/CLK line[63] vssd1 vssd1 vccd1 vccd1 _10653_/A sky130_fd_sc_hd__dfxtp_1
X_13371_ _13371_/A _13404_/Y vssd1 vssd1 vccd1 vccd1 _13651_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13859__A _13899_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10583_ _10583_/A _10604_/Y vssd1 vssd1 vccd1 vccd1 _13663_/Z sky130_fd_sc_hd__ebufn_2
X_12322_ _12350_/CLK line[58] vssd1 vssd1 vccd1 vccd1 _12323_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13578__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12253_ _12253_/A _12284_/Y vssd1 vssd1 vccd1 vccd1 _13653_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_181_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[19\].VALID\[14\].TOBUF OVHB\[19\].VALID\[14\].FF/Q OVHB\[19\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/B2 sky130_fd_sc_hd__ebufn_2
X_11204_ _11230_/CLK line[59] vssd1 vssd1 vccd1 vccd1 _11205_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06911__D line[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12184_ _12210_/CLK line[123] vssd1 vssd1 vccd1 vccd1 _12185_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11529__D line[65] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11135_ _11135_/A _11164_/Y vssd1 vssd1 vccd1 vccd1 _13655_/Z sky130_fd_sc_hd__ebufn_2
X_11066_ _11090_/CLK line[124] vssd1 vssd1 vccd1 vccd1 _11067_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[17\].VALID\[11\].FF_D A[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13744__D line[54] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10017_ _10017_/A _10044_/Y vssd1 vssd1 vccd1 vccd1 _13657_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08838__D line[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12003__A _13934_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11968_ _13934_/X wr vssd1 vssd1 vccd1 vccd1 _11968_/X sky130_fd_sc_hd__and2_1
XDATA\[2\].CLKBUF\[1\] clk vssd1 vssd1 vccd1 vccd1 _11162_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__05262__D line[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13707_ _13715_/CLK line[37] vssd1 vssd1 vccd1 vccd1 _13708_/A sky130_fd_sc_hd__dfxtp_1
X_10919_ _13925_/X vssd1 vssd1 vccd1 vccd1 _10919_/Y sky130_fd_sc_hd__inv_2
X_11899_ _13927_/X vssd1 vssd1 vccd1 vccd1 _11899_/Y sky130_fd_sc_hd__inv_2
XFILLER_189_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[12\].VALID\[13\].TOBUF OVHB\[12\].VALID\[13\].FF/Q OVHB\[12\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04916_/B2 sky130_fd_sc_hd__ebufn_2
XOVHB\[13\].VALID\[6\].FF OVHB\[13\].V/CLK A[13] vssd1 vssd1 vccd1 vccd1 OVHB\[13\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_13638_ _13638_/A _13649_/Y vssd1 vssd1 vccd1 vccd1 _13638_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_158_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[27\].VALID\[10\].FF_D A[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[22\].CLKBUF\[7\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12095__D line[68] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[20\].CGAND _13913_/X wr vssd1 vssd1 vccd1 vccd1 OVHB\[20\].CGAND/X sky130_fd_sc_hd__and2_4
X_13569_ _13575_/CLK line[102] vssd1 vssd1 vccd1 vccd1 _13570_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07189__D line[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06110_ _06120_/CLK line[20] vssd1 vssd1 vccd1 vccd1 _06111_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_8_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07090_ _07100_/CLK line[84] vssd1 vssd1 vccd1 vccd1 _07091_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_172_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06041_ _06041_/A _06054_/Y vssd1 vssd1 vccd1 vccd1 _13881_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_160_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10343__D line[35] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09800_ _09830_/CLK line[48] vssd1 vssd1 vccd1 vccd1 _09801_/A sky130_fd_sc_hd__dfxtp_1
X_07992_ _08010_/CLK line[127] vssd1 vssd1 vccd1 vccd1 _07993_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05437__D line[111] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09731_ _09731_/A _09764_/Y vssd1 vssd1 vccd1 vccd1 _13651_/Z sky130_fd_sc_hd__ebufn_2
X_06943_ _06943_/A _06964_/Y vssd1 vssd1 vccd1 vccd1 _13663_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[18\].VALID\[2\].TOBUF OVHB\[18\].VALID\[2\].FF/Q OVHB\[18\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04930_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__13654__D line[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDATA\[22\].CLKBUF\[5\] clk vssd1 vssd1 vccd1 vccd1 _09062_/CLK sky130_fd_sc_hd__clkbuf_4
X_09662_ _09690_/CLK line[122] vssd1 vssd1 vccd1 vccd1 _09663_/A sky130_fd_sc_hd__dfxtp_1
X_06874_ _06890_/CLK line[113] vssd1 vssd1 vccd1 vccd1 _06875_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_28_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07652__D line[85] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08613_ _08613_/A _08644_/Y vssd1 vssd1 vccd1 vccd1 _13653_/Z sky130_fd_sc_hd__ebufn_2
X_05825_ _05825_/A _05844_/Y vssd1 vssd1 vccd1 vccd1 _13665_/Z sky130_fd_sc_hd__ebufn_2
X_09593_ _09593_/A _09624_/Y vssd1 vssd1 vccd1 vccd1 _13793_/Z sky130_fd_sc_hd__ebufn_2
X_08544_ _08570_/CLK line[123] vssd1 vssd1 vccd1 vccd1 _08545_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05756_ _05770_/CLK line[114] vssd1 vssd1 vccd1 vccd1 _05757_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08475_ _08475_/A _08504_/Y vssd1 vssd1 vccd1 vccd1 _13795_/Z sky130_fd_sc_hd__ebufn_2
X_05687_ _05687_/A _05704_/Y vssd1 vssd1 vccd1 vccd1 _13807_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11902__D line[122] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09579__D line[70] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07426_ _07450_/CLK line[124] vssd1 vssd1 vccd1 vccd1 _07427_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05900__D line[52] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07357_ _07357_/A _07384_/Y vssd1 vssd1 vccd1 vccd1 _13797_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10518__D line[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06308_ _06330_/CLK line[125] vssd1 vssd1 vccd1 vccd1 _06309_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_176_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07288_ _07310_/CLK line[61] vssd1 vssd1 vccd1 vccd1 _07289_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_191_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13829__D line[107] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09027_ _09027_/CLK _09028_/X vssd1 vssd1 vccd1 vccd1 _09025_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__11199__A _13933_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12733__D line[104] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06239_ _06239_/A _06264_/Y vssd1 vssd1 vccd1 vccd1 _13799_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[20\].VALID\[6\].FF_D A[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[11\].VALID\[8\].FF OVHB\[11\].V/CLK A[15] vssd1 vssd1 vccd1 vccd1 OVHB\[11\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07827__D line[37] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[13\].CG_CLK clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09929_ _09935_/CLK line[102] vssd1 vssd1 vccd1 vccd1 _09930_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_105_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12940_ _12940_/A _12949_/Y vssd1 vssd1 vccd1 vccd1 _13780_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07562__D line[58] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MUX.M\[0\].MUX\[7\]_A1 _13712_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11084__D line[118] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12871_ _12875_/CLK line[39] vssd1 vssd1 vccd1 vccd1 _12872_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06178__D line[51] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11822_ _11822_/A _11829_/Y vssd1 vssd1 vccd1 vccd1 _13782_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[21\].CLKBUF\[2\] clk vssd1 vssd1 vccd1 vccd1 _08677_/CLK sky130_fd_sc_hd__clkbuf_4
XPHY_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11753_ _11755_/CLK line[40] vssd1 vssd1 vccd1 vccd1 _11754_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12908__D line[56] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[24\].VALID\[1\].TOBUF OVHB\[24\].VALID\[1\].FF/Q OVHB\[24\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04926_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_41_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09489__D line[43] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10704_ _10704_/A _10709_/Y vssd1 vssd1 vccd1 vccd1 _13784_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08393__D line[40] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11684_ _11684_/A _11689_/Y vssd1 vssd1 vccd1 vccd1 _13644_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05810__D line[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10635_ _10635_/CLK line[41] vssd1 vssd1 vccd1 vccd1 _10636_/A sky130_fd_sc_hd__dfxtp_1
X_13423_ _13435_/CLK line[35] vssd1 vssd1 vccd1 vccd1 _13424_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12493__A _13935_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13354_ _13354_/A _13369_/Y vssd1 vssd1 vccd1 vccd1 _13634_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_139_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10566_ _10566_/A _10569_/Y vssd1 vssd1 vccd1 vccd1 _13646_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_127_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12305_ _12315_/CLK line[36] vssd1 vssd1 vccd1 vccd1 _12306_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_6_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12643__D line[77] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13285_ _13295_/CLK line[100] vssd1 vssd1 vccd1 vccd1 _13286_/A sky130_fd_sc_hd__dfxtp_1
X_10497_ _10497_/CLK _10498_/X vssd1 vssd1 vccd1 vccd1 _10495_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__07737__D line[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06641__D line[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12236_ _12236_/A _12249_/Y vssd1 vssd1 vccd1 vccd1 _13636_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_5_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11259__D line[70] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12167_ _12175_/CLK line[101] vssd1 vssd1 vccd1 vccd1 _12168_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09952__D line[127] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11118_ _11118_/A _11129_/Y vssd1 vssd1 vccd1 vccd1 _13638_/Z sky130_fd_sc_hd__ebufn_2
X_12098_ _12098_/A _12109_/Y vssd1 vssd1 vccd1 vccd1 _13778_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_49_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08568__D line[120] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11049_ _11055_/CLK line[102] vssd1 vssd1 vccd1 vccd1 _11050_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[1\].VALID\[1\].FF_D A[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12668__A _13936_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05610_ _05630_/CLK line[62] vssd1 vssd1 vccd1 vccd1 _05611_/A sky130_fd_sc_hd__dfxtp_1
X_06590_ _06610_/CLK line[126] vssd1 vssd1 vccd1 vccd1 _06591_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_33_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05541_ _05541_/A _05564_/Y vssd1 vssd1 vccd1 vccd1 _13661_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12818__D line[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08260_ _08290_/CLK line[112] vssd1 vssd1 vccd1 vccd1 _08261_/A sky130_fd_sc_hd__dfxtp_1
X_05472_ _05490_/CLK line[127] vssd1 vssd1 vccd1 vccd1 _05473_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06816__D line[87] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07211_ _07211_/A _07244_/Y vssd1 vssd1 vccd1 vccd1 _13651_/Z sky130_fd_sc_hd__ebufn_2
X_08191_ _08191_/A _08224_/Y vssd1 vssd1 vccd1 vccd1 _13791_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[16\].VALID\[7\].TOBUF OVHB\[16\].VALID\[7\].FF/Q OVHB\[16\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/A2 sky130_fd_sc_hd__ebufn_2
X_07142_ _07170_/CLK line[122] vssd1 vssd1 vccd1 vccd1 _07143_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[10\].CLKBUF\[5\] clk vssd1 vssd1 vccd1 vccd1 _05422_/CLK sky130_fd_sc_hd__clkbuf_4
X_07073_ _07073_/A _07104_/Y vssd1 vssd1 vccd1 vccd1 _13793_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_105_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06551__D line[108] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06024_ _06050_/CLK line[123] vssd1 vssd1 vccd1 vccd1 _06025_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[30\].VALID\[0\].TOBUF OVHB\[30\].VALID\[0\].FF/Q OVHB\[30\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04924_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__11169__D line[43] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10073__D line[40] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05167__D line[101] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07975_ _07975_/CLK line[105] vssd1 vssd1 vccd1 vccd1 _07976_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13384__D line[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13962__A A_h[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06926_ _06926_/A _06929_/Y vssd1 vssd1 vccd1 vccd1 _13646_/Z sky130_fd_sc_hd__ebufn_2
X_09714_ _09714_/A _09729_/Y vssd1 vssd1 vccd1 vccd1 _13634_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_142_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08478__D line[93] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09645_ _09655_/CLK line[100] vssd1 vssd1 vccd1 vccd1 _09646_/A sky130_fd_sc_hd__dfxtp_1
X_06857_ _06857_/CLK _06858_/X vssd1 vssd1 vccd1 vccd1 _06855_/CLK sky130_fd_sc_hd__dlclkp_1
X_05808_ _13902_/X wr vssd1 vssd1 vccd1 vccd1 _05808_/X sky130_fd_sc_hd__and2_1
XFILLER_83_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09576_ _09576_/A _09589_/Y vssd1 vssd1 vccd1 vccd1 _13776_/Z sky130_fd_sc_hd__ebufn_2
X_06788_ _13905_/X wr vssd1 vssd1 vccd1 vccd1 _06788_/X sky130_fd_sc_hd__and2_1
XFILLER_35_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08527_ _08535_/CLK line[101] vssd1 vssd1 vccd1 vccd1 _08528_/A sky130_fd_sc_hd__dfxtp_1
XPHY_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05739_ _13901_/X vssd1 vssd1 vccd1 vccd1 _05739_/Y sky130_fd_sc_hd__inv_2
XANTENNA__04930__B1 A_h[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11632__D line[127] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08458_ _08458_/A _08469_/Y vssd1 vssd1 vccd1 vccd1 _13778_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06726__D line[60] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05630__D line[57] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09102__D line[122] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07409_ _07415_/CLK line[102] vssd1 vssd1 vccd1 vccd1 _07410_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10248__D line[120] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08389_ _08395_/CLK line[38] vssd1 vssd1 vccd1 vccd1 _08390_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10420_ _10420_/A _10429_/Y vssd1 vssd1 vccd1 vccd1 _13780_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08941__D line[34] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13559__D line[97] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10351_ _10355_/CLK line[39] vssd1 vssd1 vccd1 vccd1 _10352_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_152_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13070_ _13070_/A _13089_/Y vssd1 vssd1 vccd1 vccd1 _13630_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_183_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10282_ _10282_/A _10289_/Y vssd1 vssd1 vccd1 vccd1 _13642_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XOVHB\[4\].VALID\[1\].FF OVHB\[4\].V/CLK A[8] vssd1 vssd1 vccd1 vccd1 OVHB\[4\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_183_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12021_ _12035_/CLK line[34] vssd1 vssd1 vccd1 vccd1 _12022_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_151_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05077__D line[74] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[22\].VALID\[6\].TOBUF OVHB\[22\].VALID\[6\].FF/Q OVHB\[22\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04923_/A2 sky130_fd_sc_hd__ebufn_2
XANTENNA__11807__D line[79] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13972_ A_h[0] vssd1 vssd1 vccd1 vccd1 _13982_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__05805__D line[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07292__D line[63] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12923_ _12945_/CLK line[77] vssd1 vssd1 vccd1 vccd1 _12924_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_18_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XOVHB\[6\].VALID\[10\].TOBUF OVHB\[6\].VALID\[10\].FF/Q OVHB\[6\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04932_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_18_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12854_ _12854_/A _12879_/Y vssd1 vssd1 vccd1 vccd1 _13694_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_61_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11805_ _11825_/CLK line[78] vssd1 vssd1 vccd1 vccd1 _11806_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[7\].VALID\[5\].FF_D A[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12785_ _12805_/CLK line[14] vssd1 vssd1 vccd1 vccd1 _12786_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_159_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11736_ _11736_/A _11759_/Y vssd1 vssd1 vccd1 vccd1 _13696_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05540__D line[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[14\].CGAND_B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10158__D line[93] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11667_ _11685_/CLK line[15] vssd1 vssd1 vccd1 vccd1 _11668_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13406_ _13406_/A _13439_/Y vssd1 vssd1 vccd1 vccd1 _13686_/Z sky130_fd_sc_hd__ebufn_2
X_10618_ _10618_/A _10639_/Y vssd1 vssd1 vccd1 vccd1 _13698_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11598_ _11598_/A _11619_/Y vssd1 vssd1 vccd1 vccd1 _13838_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_128_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_OVHB\[18\].CGAND_A _13911_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[18\].V_RESET_B rst_n vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12373__D line[67] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10549_ _10565_/CLK line[1] vssd1 vssd1 vccd1 vccd1 _10550_/A sky130_fd_sc_hd__dfxtp_1
X_13337_ _13365_/CLK line[10] vssd1 vssd1 vccd1 vccd1 _13338_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07467__D line[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13268_ _13268_/A _13299_/Y vssd1 vssd1 vccd1 vccd1 _13828_/Z sky130_fd_sc_hd__ebufn_2
X_12219_ _12245_/CLK line[11] vssd1 vssd1 vccd1 vccd1 _12220_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[15\].CLKBUF\[1\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13199_ _13225_/CLK line[75] vssd1 vssd1 vccd1 vccd1 _13200_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09682__D line[117] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10621__D line[34] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07760_ _07760_/A _07769_/Y vssd1 vssd1 vccd1 vccd1 _13640_/Z sky130_fd_sc_hd__ebufn_2
X_04972_ _05000_/CLK line[26] vssd1 vssd1 vccd1 vccd1 _04973_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_49_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05715__D line[110] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06711_ _06715_/CLK line[39] vssd1 vssd1 vccd1 vccd1 _06712_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_37_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[2\].VALID\[3\].FF OVHB\[2\].V/CLK A[10] vssd1 vssd1 vccd1 vccd1 OVHB\[2\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_07691_ _07695_/CLK line[103] vssd1 vssd1 vccd1 vccd1 _07692_/A sky130_fd_sc_hd__dfxtp_1
X_09430_ _09430_/A _09449_/Y vssd1 vssd1 vccd1 vccd1 _13630_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_37_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06642_ _06642_/A _06649_/Y vssd1 vssd1 vccd1 vccd1 _13642_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_80_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07930__D line[84] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09361_ _09375_/CLK line[98] vssd1 vssd1 vccd1 vccd1 _09362_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__04912__B1 _04912_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12548__D line[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06573_ _06575_/CLK line[104] vssd1 vssd1 vccd1 vccd1 _06574_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_80_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08312_ _08312_/A _08329_/Y vssd1 vssd1 vccd1 vccd1 _13632_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_178_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05524_ _05524_/A _05529_/Y vssd1 vssd1 vccd1 vccd1 _13644_/Z sky130_fd_sc_hd__ebufn_2
X_09292_ _09292_/A _09309_/Y vssd1 vssd1 vccd1 vccd1 _13772_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[8\].CLKBUF\[1\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08243_ _08255_/CLK line[99] vssd1 vssd1 vccd1 vccd1 _08244_/A sky130_fd_sc_hd__dfxtp_1
X_05455_ _05455_/CLK line[105] vssd1 vssd1 vccd1 vccd1 _05456_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_138_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09857__D line[69] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08174_ _08174_/A _08189_/Y vssd1 vssd1 vccd1 vccd1 _13774_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_21_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05386_ _05386_/A _05389_/Y vssd1 vssd1 vccd1 vccd1 _13786_/Z sky130_fd_sc_hd__ebufn_2
X_07125_ _07135_/CLK line[100] vssd1 vssd1 vccd1 vccd1 _07126_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_137_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06281__D line[98] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07056_ _07056_/A _07069_/Y vssd1 vssd1 vccd1 vccd1 _13776_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_173_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06007_ _06015_/CLK line[101] vssd1 vssd1 vccd1 vccd1 _06008_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09592__D line[90] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07958_ _07958_/A _07979_/Y vssd1 vssd1 vccd1 vccd1 _13838_/Z sky130_fd_sc_hd__ebufn_2
X_06909_ _06925_/CLK line[1] vssd1 vssd1 vccd1 vccd1 _06910_/A sky130_fd_sc_hd__dfxtp_1
X_07889_ _07905_/CLK line[65] vssd1 vssd1 vccd1 vccd1 _07890_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_56_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09628_ _09628_/A _09659_/Y vssd1 vssd1 vccd1 vccd1 _13828_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07840__D line[48] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XOVHB\[29\].VALID\[12\].TOBUF OVHB\[29\].VALID\[12\].FF/Q OVHB\[29\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04929_/B2 sky130_fd_sc_hd__ebufn_2
XPHY_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09559_ _09585_/CLK line[75] vssd1 vssd1 vccd1 vccd1 _09560_/A sky130_fd_sc_hd__dfxtp_1
XPHY_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11362__D line[117] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06456__D line[50] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12570_ _12570_/A _12599_/Y vssd1 vssd1 vccd1 vccd1 _13690_/Z sky130_fd_sc_hd__ebufn_2
XPHY_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[0\].VALID\[5\].FF OVHB\[0\].V/CLK A[12] vssd1 vssd1 vccd1 vccd1 OVHB\[0\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11521_ _11545_/CLK line[76] vssd1 vssd1 vccd1 vccd1 _11522_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_178_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09767__D line[42] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06753__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11452_ _11452_/A _11479_/Y vssd1 vssd1 vccd1 vccd1 _13692_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08671__D line[39] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13289__D line[102] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10403_ _10425_/CLK line[77] vssd1 vssd1 vccd1 vccd1 _10404_/A sky130_fd_sc_hd__dfxtp_1
X_11383_ _11405_/CLK line[13] vssd1 vssd1 vccd1 vccd1 _11384_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_125_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13122_ _13122_/CLK _13123_/X vssd1 vssd1 vccd1 vccd1 _13120_/CLK sky130_fd_sc_hd__dlclkp_1
X_10334_ _10334_/A _10359_/Y vssd1 vssd1 vccd1 vccd1 _13694_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_11_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12921__D line[76] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13053_ _13937_/X wr vssd1 vssd1 vccd1 vccd1 _13053_/X sky130_fd_sc_hd__and2_1
X_10265_ _10285_/CLK line[14] vssd1 vssd1 vccd1 vccd1 _10266_/A sky130_fd_sc_hd__dfxtp_1
X_12004_ _13934_/X vssd1 vssd1 vccd1 vccd1 _12004_/Y sky130_fd_sc_hd__inv_2
X_10196_ _10196_/A _10219_/Y vssd1 vssd1 vccd1 vccd1 _13836_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11537__D line[69] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__04927__A2_N _04927_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XOVHB\[22\].VALID\[11\].TOBUF OVHB\[22\].VALID\[11\].FF/Q OVHB\[22\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04915_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__09007__D line[79] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13955_ _13960_/C _13960_/A _13960_/B _13960_/D vssd1 vssd1 vccd1 vccd1 _13955_/X
+ sky130_fd_sc_hd__and4bb_4
XFILLER_19_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06928__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12906_ _12910_/CLK line[55] vssd1 vssd1 vccd1 vccd1 _12907_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_47_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08846__D line[119] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13886_ _13890_/CLK line[119] vssd1 vssd1 vccd1 vccd1 _13887_/A sky130_fd_sc_hd__dfxtp_1
X_12837_ _12837_/A _12844_/Y vssd1 vssd1 vccd1 vccd1 _13677_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11272__D line[90] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05270__D line[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12768_ _12770_/CLK line[120] vssd1 vssd1 vccd1 vccd1 _12769_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11719_ _11719_/A _11724_/Y vssd1 vssd1 vccd1 vccd1 _13679_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_159_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12699_ _12699_/A _12704_/Y vssd1 vssd1 vccd1 vccd1 _13819_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08581__D line[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05240_ _05240_/A _05249_/Y vssd1 vssd1 vccd1 vccd1 _13640_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_30_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13199__D line[75] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05171_ _05175_/CLK line[103] vssd1 vssd1 vccd1 vccd1 _05172_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07197__D line[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08930_ _08930_/A _08959_/Y vssd1 vssd1 vccd1 vccd1 _13690_/Z sky130_fd_sc_hd__ebufn_2
X_08861_ _08885_/CLK line[12] vssd1 vssd1 vccd1 vccd1 _08862_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11447__D line[42] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10351__D line[39] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[4\].VALID\[3\].TOBUF OVHB\[4\].VALID\[3\].FF/Q OVHB\[4\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04919_/B2 sky130_fd_sc_hd__ebufn_2
X_07812_ _07812_/A _07839_/Y vssd1 vssd1 vccd1 vccd1 _13692_/Z sky130_fd_sc_hd__ebufn_2
X_08792_ _08792_/A _08819_/Y vssd1 vssd1 vccd1 vccd1 _13832_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05445__D line[100] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[2\].VALID\[14\].FF_D A[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[29\].VALID\[6\].TOBUF OVHB\[29\].VALID\[6\].FF/Q OVHB\[29\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04923_/A2 sky130_fd_sc_hd__ebufn_2
XFILLER_38_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07743_ _07765_/CLK line[13] vssd1 vssd1 vccd1 vccd1 _07744_/A sky130_fd_sc_hd__dfxtp_1
X_04955_ _04965_/CLK line[4] vssd1 vssd1 vccd1 vccd1 _04956_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_84_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13662__D line[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[13\].CLKBUF\[3\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08756__D line[92] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07674_ _07674_/A _07699_/Y vssd1 vssd1 vccd1 vccd1 _13834_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07660__D line[89] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[27\].VALID\[0\].FF OVHB\[27\].V/CLK A[7] vssd1 vssd1 vccd1 vccd1 OVHB\[27\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_09413_ _13916_/X wr vssd1 vssd1 vccd1 vccd1 _09413_/X sky130_fd_sc_hd__and2_1
X_06625_ _06645_/CLK line[14] vssd1 vssd1 vccd1 vccd1 _06626_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12278__D line[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[12\].VALID\[1\].FF_D A[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09344_ _13916_/X vssd1 vssd1 vccd1 vccd1 _09344_/Y sky130_fd_sc_hd__inv_2
X_06556_ _06556_/A _06579_/Y vssd1 vssd1 vccd1 vccd1 _13836_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05180__D line[112] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05507_ _05525_/CLK line[15] vssd1 vssd1 vccd1 vccd1 _05508_/A sky130_fd_sc_hd__dfxtp_1
X_09275_ _09305_/CLK line[64] vssd1 vssd1 vccd1 vccd1 _09276_/A sky130_fd_sc_hd__dfxtp_1
X_06487_ _06505_/CLK line[79] vssd1 vssd1 vccd1 vccd1 _06488_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11910__D line[126] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08226_ _08226_/A _08259_/Y vssd1 vssd1 vccd1 vccd1 _13826_/Z sky130_fd_sc_hd__ebufn_2
X_05438_ _05438_/A _05459_/Y vssd1 vssd1 vccd1 vccd1 _13838_/Z sky130_fd_sc_hd__ebufn_2
X_08157_ _08185_/CLK line[74] vssd1 vssd1 vccd1 vccd1 _08158_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10526__D line[119] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05369_ _05385_/CLK line[65] vssd1 vssd1 vccd1 vccd1 _05370_/A sky130_fd_sc_hd__dfxtp_1
X_07108_ _07108_/A _07139_/Y vssd1 vssd1 vccd1 vccd1 _13828_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[6\].CLKBUF\[3\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08088_ _08088_/A _08119_/Y vssd1 vssd1 vccd1 vccd1 _13688_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13837__D line[111] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07039_ _07065_/CLK line[75] vssd1 vssd1 vccd1 vccd1 _07040_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07835__D line[41] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10050_ _10050_/A _10079_/Y vssd1 vssd1 vccd1 vccd1 _13690_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_0_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10261__D line[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05355__D line[64] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XDATA\[31\].CLKBUF\[7\] clk vssd1 vssd1 vccd1 vccd1 _11932_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_28_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_OVHB\[3\].VALID\[8\].FF_D A[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13740_ _13750_/CLK line[52] vssd1 vssd1 vccd1 vccd1 _13741_/A sky130_fd_sc_hd__dfxtp_1
X_10952_ _10952_/CLK _10953_/X vssd1 vssd1 vccd1 vccd1 _10950_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__07570__D line[62] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12188__D line[125] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13671_ _13671_/A _13684_/Y vssd1 vssd1 vccd1 vccd1 _13671_/Z sky130_fd_sc_hd__ebufn_2
X_10883_ _13925_/X wr vssd1 vssd1 vccd1 vccd1 _10883_/X sky130_fd_sc_hd__and2_1
XPHY_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06186__D line[55] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12622_ _12630_/CLK line[53] vssd1 vssd1 vccd1 vccd1 _12623_/A sky130_fd_sc_hd__dfxtp_1
XPHY_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12553_ _12553_/A _12564_/Y vssd1 vssd1 vccd1 vccd1 _13673_/Z sky130_fd_sc_hd__ebufn_2
XPHY_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09497__D line[47] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11504_ _11510_/CLK line[54] vssd1 vssd1 vccd1 vccd1 _11505_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[25\].VALID\[2\].FF OVHB\[25\].V/CLK A[9] vssd1 vssd1 vccd1 vccd1 OVHB\[25\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12484_ _12490_/CLK line[118] vssd1 vssd1 vccd1 vccd1 _12485_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10436__D line[92] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11435_ _11435_/A _11444_/Y vssd1 vssd1 vccd1 vccd1 _13675_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[4\].VALID\[10\].FF_D A[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XDATA\[0\].CLKBUF\[6\] clk vssd1 vssd1 vccd1 vccd1 _05177_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_98_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11366_ _11370_/CLK line[119] vssd1 vssd1 vccd1 vccd1 _11367_/A sky130_fd_sc_hd__dfxtp_1
X_13105_ _13105_/A _13124_/Y vssd1 vssd1 vccd1 vccd1 _13665_/Z sky130_fd_sc_hd__ebufn_2
X_10317_ _10317_/A _10324_/Y vssd1 vssd1 vccd1 vccd1 _13677_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12651__D line[66] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11297_ _11297_/A _11304_/Y vssd1 vssd1 vccd1 vccd1 _13817_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07745__D line[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10248_ _10250_/CLK line[120] vssd1 vssd1 vccd1 vccd1 _10249_/A sky130_fd_sc_hd__dfxtp_1
X_13036_ _13050_/CLK line[114] vssd1 vssd1 vccd1 vccd1 _13037_/A sky130_fd_sc_hd__dfxtp_1
X_10179_ _10179_/A _10184_/Y vssd1 vssd1 vccd1 vccd1 _13819_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09960__D line[116] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05843__A _13902_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13938_ _13938_/A _13938_/B _13938_/C _13938_/D vssd1 vssd1 vccd1 vccd1 _13938_/X
+ sky130_fd_sc_hd__and4_4
XANTENNA_OVHB\[25\].VALID\[1\].FF_D A[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13869_ _13869_/A _13894_/Y vssd1 vssd1 vccd1 vccd1 _13869_/Z sky130_fd_sc_hd__ebufn_2
X_06410_ _06410_/A _06439_/Y vssd1 vssd1 vccd1 vccd1 _13690_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[30\].CLKBUF\[4\] clk vssd1 vssd1 vccd1 vccd1 _11547_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_179_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06096__D line[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07390_ _07390_/A _07419_/Y vssd1 vssd1 vccd1 vccd1 _13830_/Z sky130_fd_sc_hd__ebufn_2
X_06341_ _06365_/CLK line[12] vssd1 vssd1 vccd1 vccd1 _06342_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12826__D line[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XOVHB\[22\].VALID\[13\].FF OVHB\[22\].V/CLK A[20] vssd1 vssd1 vccd1 vccd1 OVHB\[22\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_09060_ _09060_/CLK line[89] vssd1 vssd1 vccd1 vccd1 _09061_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[18\].VALID\[5\].FF_D A[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[2\].VALID\[8\].TOBUF OVHB\[2\].VALID\[8\].FF/Q OVHB\[2\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04931_/B2 sky130_fd_sc_hd__ebufn_2
X_06272_ _06272_/A _06299_/Y vssd1 vssd1 vccd1 vccd1 _13832_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09200__D line[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08011_ _08011_/A _08014_/Y vssd1 vssd1 vccd1 vccd1 _13891_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_163_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05223_ _05245_/CLK line[13] vssd1 vssd1 vccd1 vccd1 _05224_/A sky130_fd_sc_hd__dfxtp_1
X_05154_ _05154_/A _05179_/Y vssd1 vssd1 vccd1 vccd1 _13834_/Z sky130_fd_sc_hd__ebufn_2
XMUX.SEL1BUF\[3\] A[1] vssd1 vssd1 vccd1 vccd1 MUX.SEL1BUF\[3\]/X sky130_fd_sc_hd__clkbuf_2
XFILLER_143_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09962_ _09970_/CLK line[117] vssd1 vssd1 vccd1 vccd1 _09963_/A sky130_fd_sc_hd__dfxtp_1
X_05085_ _05105_/CLK line[78] vssd1 vssd1 vccd1 vccd1 _05086_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_171_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XOVHB\[23\].VALID\[4\].FF OVHB\[23\].V/CLK A[11] vssd1 vssd1 vccd1 vccd1 OVHB\[23\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_08913_ _08913_/A _08924_/Y vssd1 vssd1 vccd1 vccd1 _13673_/Z sky130_fd_sc_hd__ebufn_2
X_09893_ _09893_/A _09904_/Y vssd1 vssd1 vccd1 vccd1 _13813_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11177__D line[47] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08844_ _08850_/CLK line[118] vssd1 vssd1 vccd1 vccd1 _08845_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05175__D line[105] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09870__D line[80] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XOVHB\[15\].CGAND _13905_/X wr vssd1 vssd1 vccd1 vccd1 OVHB\[15\].CGAND/X sky130_fd_sc_hd__and2_4
XFILLER_27_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05987_ _06015_/CLK line[106] vssd1 vssd1 vccd1 vccd1 _05988_/A sky130_fd_sc_hd__dfxtp_1
X_08775_ _08775_/A _08784_/Y vssd1 vssd1 vccd1 vccd1 _13815_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13392__D line[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_04938_ _04938_/A _04969_/Y vssd1 vssd1 vccd1 vccd1 _13618_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08486__D line[82] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07726_ _07730_/CLK line[119] vssd1 vssd1 vccd1 vccd1 _07727_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_84_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07657_ _07657_/A _07664_/Y vssd1 vssd1 vccd1 vccd1 _13817_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08783__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06608_ _06610_/CLK line[120] vssd1 vssd1 vccd1 vccd1 _06609_/A sky130_fd_sc_hd__dfxtp_1
X_07588_ _07590_/CLK line[56] vssd1 vssd1 vccd1 vccd1 _07589_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_43_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_DATA\[11\].CLKBUF\[5\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09327_ _09327_/A _09344_/Y vssd1 vssd1 vccd1 vccd1 _13807_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_40_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06539_ _06539_/A _06544_/Y vssd1 vssd1 vccd1 vccd1 _13819_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_178_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11640__D line[116] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06734__D line[49] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09258_ _09270_/CLK line[51] vssd1 vssd1 vccd1 vccd1 _09259_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09110__D line[126] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08209_ _08209_/A _08224_/Y vssd1 vssd1 vccd1 vccd1 _13809_/Z sky130_fd_sc_hd__ebufn_2
X_09189_ _09189_/A _09204_/Y vssd1 vssd1 vccd1 vccd1 _13669_/Z sky130_fd_sc_hd__ebufn_2
X_11220_ _11230_/CLK line[52] vssd1 vssd1 vccd1 vccd1 _11221_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13567__D line[101] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11151_ _11151_/A _11164_/Y vssd1 vssd1 vccd1 vccd1 _13671_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_108_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10102_ _10110_/CLK line[53] vssd1 vssd1 vccd1 vccd1 _10103_/A sky130_fd_sc_hd__dfxtp_1
X_11082_ _11090_/CLK line[117] vssd1 vssd1 vccd1 vccd1 _11083_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08958__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10033_ _10033_/A _10044_/Y vssd1 vssd1 vccd1 vccd1 _13673_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[4\].CLKBUF\[5\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05085__D line[78] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11815__D line[68] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XOVHB\[21\].VALID\[6\].FF OVHB\[21\].V/CLK A[13] vssd1 vssd1 vccd1 vccd1 OVHB\[21\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06909__D line[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11984_ _12000_/CLK line[17] vssd1 vssd1 vccd1 vccd1 _11985_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[9\].VALID\[14\].FF_D A[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[30\].CLKBUF\[7\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[19\].VALID\[10\].TOBUF OVHB\[19\].VALID\[10\].FF/Q OVHB\[19\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04932_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_189_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13723_ _13723_/A _13754_/Y vssd1 vssd1 vccd1 vccd1 _13723_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_17_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10935_ _10935_/A _10954_/Y vssd1 vssd1 vccd1 vccd1 _13735_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_16_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13654_ _13680_/CLK line[27] vssd1 vssd1 vccd1 vccd1 _13655_/A sky130_fd_sc_hd__dfxtp_1
X_10866_ _10880_/CLK line[18] vssd1 vssd1 vccd1 vccd1 _10867_/A sky130_fd_sc_hd__dfxtp_1
X_12605_ _12605_/A _12634_/Y vssd1 vssd1 vccd1 vccd1 _13725_/Z sky130_fd_sc_hd__ebufn_2
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11550__D line[80] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13585_ _13585_/A _13614_/Y vssd1 vssd1 vccd1 vccd1 _13865_/Z sky130_fd_sc_hd__ebufn_2
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XOVHB\[27\].CG clk OVHB\[27\].CGAND/X vssd1 vssd1 vccd1 vccd1 OVHB\[27\].V/CLK sky130_fd_sc_hd__dlclkp_1
X_10797_ _10797_/A _10814_/Y vssd1 vssd1 vccd1 vccd1 _13877_/Z sky130_fd_sc_hd__ebufn_2
XPHY_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12536_ _12560_/CLK line[28] vssd1 vssd1 vccd1 vccd1 _12537_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_157_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10166__D line[82] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10744__A _13924_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12467_ _12467_/A _12494_/Y vssd1 vssd1 vccd1 vccd1 _13867_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_157_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11418_ _11440_/CLK line[29] vssd1 vssd1 vccd1 vccd1 _11419_/A sky130_fd_sc_hd__dfxtp_1
X_12398_ _12420_/CLK line[93] vssd1 vssd1 vccd1 vccd1 _12399_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10463__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13477__D line[74] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12381__D line[71] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11349_ _11349_/A _11374_/Y vssd1 vssd1 vccd1 vccd1 _13869_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07475__D line[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05910_ _05910_/CLK line[57] vssd1 vssd1 vccd1 vccd1 _05911_/A sky130_fd_sc_hd__dfxtp_1
X_13019_ _13937_/X vssd1 vssd1 vccd1 vccd1 _13019_/Y sky130_fd_sc_hd__inv_2
X_06890_ _06890_/CLK line[121] vssd1 vssd1 vccd1 vccd1 _06891_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09690__D line[121] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05841_ _05841_/A _05844_/Y vssd1 vssd1 vccd1 vccd1 _13681_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_55_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11725__D line[32] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08560_ _08570_/CLK line[116] vssd1 vssd1 vccd1 vccd1 _08561_/A sky130_fd_sc_hd__dfxtp_1
X_05772_ _05772_/CLK _05773_/X vssd1 vssd1 vccd1 vccd1 _05770_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__05723__D line[99] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07511_ _07511_/A _07524_/Y vssd1 vssd1 vccd1 vccd1 _13671_/Z sky130_fd_sc_hd__ebufn_2
X_08491_ _08491_/A _08504_/Y vssd1 vssd1 vccd1 vccd1 _13811_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10919__A _13925_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07442_ _07450_/CLK line[117] vssd1 vssd1 vccd1 vccd1 _07443_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_62_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10638__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12556__D line[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07373_ _07373_/A _07384_/Y vssd1 vssd1 vccd1 vccd1 _13813_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_13_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06324_ _06330_/CLK line[118] vssd1 vssd1 vccd1 vccd1 _06325_/A sky130_fd_sc_hd__dfxtp_1
X_09112_ _09130_/CLK line[127] vssd1 vssd1 vccd1 vccd1 _09113_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_129_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09043_ _09043_/A _09064_/Y vssd1 vssd1 vccd1 vccd1 _13803_/Z sky130_fd_sc_hd__ebufn_2
X_06255_ _06255_/A _06264_/Y vssd1 vssd1 vccd1 vccd1 _13815_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09865__D line[73] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05206_ _05210_/CLK line[119] vssd1 vssd1 vccd1 vccd1 _05207_/A sky130_fd_sc_hd__dfxtp_1
X_06186_ _06190_/CLK line[55] vssd1 vssd1 vccd1 vccd1 _06187_/A sky130_fd_sc_hd__dfxtp_1
X_05137_ _05137_/A _05144_/Y vssd1 vssd1 vccd1 vccd1 _13817_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10804__D line[118] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12291__D line[44] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XOVHB\[9\].VOBUF OVHB\[9\].V/Q OVHB\[9\].INV/Y vssd1 vssd1 vccd1 vccd1 _04912_/B1
+ sky130_fd_sc_hd__ebufn_2
XANTENNA__07385__D line[96] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09945_ _09945_/A _09974_/Y vssd1 vssd1 vccd1 vccd1 _13865_/Z sky130_fd_sc_hd__ebufn_2
X_05068_ _05070_/CLK line[56] vssd1 vssd1 vccd1 vccd1 _05069_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_77_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09876_ _09900_/CLK line[92] vssd1 vssd1 vccd1 vccd1 _09877_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06579__A _13904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08827_ _08827_/A _08854_/Y vssd1 vssd1 vccd1 vccd1 _13867_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_18_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06298__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08758_ _08780_/CLK line[93] vssd1 vssd1 vccd1 vccd1 _08759_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_73_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07709_ _07709_/A _07734_/Y vssd1 vssd1 vccd1 vccd1 _13869_/Z sky130_fd_sc_hd__ebufn_2
X_08689_ _08689_/A _08714_/Y vssd1 vssd1 vccd1 vccd1 _13729_/Z sky130_fd_sc_hd__ebufn_2
X_10720_ _10740_/CLK line[94] vssd1 vssd1 vccd1 vccd1 _10721_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_110_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XOVHB\[18\].VALID\[9\].FF OVHB\[18\].V/CLK A[16] vssd1 vssd1 vccd1 vccd1 OVHB\[18\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12466__D line[124] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10651_ _10651_/A _10674_/Y vssd1 vssd1 vccd1 vccd1 _13731_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11370__D line[121] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06464__D line[54] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13370_ _13400_/CLK line[16] vssd1 vssd1 vccd1 vccd1 _13371_/A sky130_fd_sc_hd__dfxtp_1
X_10582_ _10600_/CLK line[31] vssd1 vssd1 vccd1 vccd1 _10583_/A sky130_fd_sc_hd__dfxtp_1
X_12321_ _12321_/A _12354_/Y vssd1 vssd1 vccd1 vccd1 _13721_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_5_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09775__D line[46] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[9\].VALID\[8\].TOBUF OVHB\[9\].VALID\[8\].FF/Q OVHB\[9\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04931_/B2 sky130_fd_sc_hd__ebufn_2
X_12252_ _12280_/CLK line[26] vssd1 vssd1 vccd1 vccd1 _12253_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_5_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11203_ _11203_/A _11234_/Y vssd1 vssd1 vccd1 vccd1 _13723_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.M\[3\].MUX\[0\]_A0 _13679_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12183_ _12183_/A _12214_/Y vssd1 vssd1 vccd1 vccd1 _13863_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10714__D line[91] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09045__TE_B _09064_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07873__A _13912_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11134_ _11160_/CLK line[27] vssd1 vssd1 vccd1 vccd1 _11135_/A sky130_fd_sc_hd__dfxtp_1
X_11065_ _11065_/A _11094_/Y vssd1 vssd1 vccd1 vccd1 _13865_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_103_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10016_ _10040_/CLK line[28] vssd1 vssd1 vccd1 vccd1 _10017_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_48_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_OVHB\[21\].VALID\[4\].FF_D A[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12003__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11545__D line[73] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[2\].CG_CLK clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06639__D line[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09015__D line[68] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11967_ _11967_/CLK _11968_/X vssd1 vssd1 vccd1 vccd1 _11965_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA_DATA\[2\].CLKBUF\[7\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13706_ _13706_/A _13719_/Y vssd1 vssd1 vccd1 vccd1 _13706_/Z sky130_fd_sc_hd__ebufn_2
X_10918_ _13925_/X wr vssd1 vssd1 vccd1 vccd1 _10918_/X sky130_fd_sc_hd__and2_1
X_11898_ _13927_/X wr vssd1 vssd1 vccd1 vccd1 _11898_/X sky130_fd_sc_hd__and2_1
XANTENNA_OVHB\[14\].VALID\[8\].FF_D A[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13637_ _13645_/CLK line[5] vssd1 vssd1 vccd1 vccd1 _13638_/A sky130_fd_sc_hd__dfxtp_1
X_10849_ _13925_/X vssd1 vssd1 vccd1 vccd1 _10849_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11280__D line[94] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06374__D line[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13568_ _13568_/A _13579_/Y vssd1 vssd1 vccd1 vccd1 _13848_/Z sky130_fd_sc_hd__ebufn_2
X_12519_ _12525_/CLK line[6] vssd1 vssd1 vccd1 vccd1 _12520_/A sky130_fd_sc_hd__dfxtp_1
X_13499_ _13505_/CLK line[70] vssd1 vssd1 vccd1 vccd1 _13500_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06040_ _06050_/CLK line[116] vssd1 vssd1 vccd1 vccd1 _06041_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_173_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07991_ _07991_/A _08014_/Y vssd1 vssd1 vccd1 vccd1 _13871_/Z sky130_fd_sc_hd__ebufn_2
X_09730_ _09760_/CLK line[16] vssd1 vssd1 vccd1 vccd1 _09731_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[11\].VALID\[12\].FF_D A[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06942_ _06960_/CLK line[31] vssd1 vssd1 vccd1 vccd1 _06943_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_39_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09661_ _09661_/A _09694_/Y vssd1 vssd1 vccd1 vccd1 _13861_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[16\].VALID\[3\].TOBUF OVHB\[16\].VALID\[3\].FF/Q OVHB\[16\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04919_/B2 sky130_fd_sc_hd__ebufn_2
X_06873_ _06873_/A _06894_/Y vssd1 vssd1 vccd1 vccd1 _13873_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11455__D line[46] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08612_ _08640_/CLK line[26] vssd1 vssd1 vccd1 vccd1 _08613_/A sky130_fd_sc_hd__dfxtp_1
X_05824_ _05840_/CLK line[17] vssd1 vssd1 vccd1 vccd1 _05825_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06549__D line[107] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09592_ _09620_/CLK line[90] vssd1 vssd1 vccd1 vccd1 _09593_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05453__D line[104] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08543_ _08543_/A _08574_/Y vssd1 vssd1 vccd1 vccd1 _13863_/Z sky130_fd_sc_hd__ebufn_2
X_05755_ _05755_/A _05774_/Y vssd1 vssd1 vccd1 vccd1 _13875_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13670__D line[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08764__D line[81] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05686_ _05700_/CLK line[82] vssd1 vssd1 vccd1 vccd1 _05687_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08474_ _08500_/CLK line[91] vssd1 vssd1 vccd1 vccd1 _08475_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08119__A _13932_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07425_ _07425_/A _07454_/Y vssd1 vssd1 vccd1 vccd1 _13865_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[21\].VALID\[11\].FF_D A[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07356_ _07380_/CLK line[92] vssd1 vssd1 vccd1 vccd1 _07357_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_176_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06307_ _06307_/A _06334_/Y vssd1 vssd1 vccd1 vccd1 _13867_/Z sky130_fd_sc_hd__ebufn_2
X_07287_ _07287_/A _07314_/Y vssd1 vssd1 vccd1 vccd1 _13727_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_136_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09026_ _09026_/A _09029_/Y vssd1 vssd1 vccd1 vccd1 _13786_/Z sky130_fd_sc_hd__ebufn_2
X_06238_ _06260_/CLK line[93] vssd1 vssd1 vccd1 vccd1 _06239_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_123_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06169_ _06169_/A _06194_/Y vssd1 vssd1 vccd1 vccd1 _13729_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05628__D line[56] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08004__D line[118] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13845__D line[100] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[31\].VALID\[10\].FF_D A[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09928_ _09928_/A _09939_/Y vssd1 vssd1 vccd1 vccd1 _13848_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08939__D line[33] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09859_ _09865_/CLK line[70] vssd1 vssd1 vccd1 vccd1 _09860_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_85_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MUX.M\[0\].MUX\[7\]_A2 _13782_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12870_ _12870_/A _12879_/Y vssd1 vssd1 vccd1 vccd1 _13710_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05363__D line[77] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09413__A _13916_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11821_ _11825_/CLK line[71] vssd1 vssd1 vccd1 vccd1 _11822_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[27\].VALID\[8\].FF_D A[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13580__D line[112] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11752_ _11752_/A _11759_/Y vssd1 vssd1 vccd1 vccd1 _13712_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[18\].V_D TIE/HI vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12196__D line[114] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10703_ _10705_/CLK line[72] vssd1 vssd1 vccd1 vccd1 _10704_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11683_ _11685_/CLK line[8] vssd1 vssd1 vccd1 vccd1 _11684_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[22\].VALID\[2\].TOBUF OVHB\[22\].VALID\[2\].FF/Q OVHB\[22\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04930_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__12774__A _13936_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13422_ _13422_/A _13439_/Y vssd1 vssd1 vccd1 vccd1 _13702_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10634_ _10634_/A _10639_/Y vssd1 vssd1 vccd1 vccd1 _13714_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12493__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13353_ _13365_/CLK line[3] vssd1 vssd1 vccd1 vccd1 _13354_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_6_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_DATA\[23\].CLKBUF\[1\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[17\].V_RESET_B rst_n vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10565_ _10565_/CLK line[9] vssd1 vssd1 vccd1 vccd1 _10566_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_154_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12304_ _12304_/A _12319_/Y vssd1 vssd1 vccd1 vccd1 _13704_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05388__A _13900_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13284_ _13284_/A _13299_/Y vssd1 vssd1 vccd1 vccd1 _13844_/Z sky130_fd_sc_hd__ebufn_2
X_10496_ _10496_/A _10499_/Y vssd1 vssd1 vccd1 vccd1 _13856_/Z sky130_fd_sc_hd__ebufn_2
X_12235_ _12245_/CLK line[4] vssd1 vssd1 vccd1 vccd1 _12236_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10444__D line[81] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05538__D line[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12166_ _12166_/A _12179_/Y vssd1 vssd1 vccd1 vccd1 _13846_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13755__D line[64] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11117_ _11125_/CLK line[5] vssd1 vssd1 vccd1 vccd1 _11118_/A sky130_fd_sc_hd__dfxtp_1
X_12097_ _12105_/CLK line[69] vssd1 vssd1 vccd1 vccd1 _12098_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07753__D line[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11048_ _11048_/A _11059_/Y vssd1 vssd1 vccd1 vccd1 _13848_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12949__A _13937_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XOVHB\[27\].VALID\[13\].FF OVHB\[27\].V/CLK A[20] vssd1 vssd1 vccd1 vccd1 OVHB\[27\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12668__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12999_ _13015_/CLK line[97] vssd1 vssd1 vccd1 vccd1 _13000_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_33_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05540_ _05560_/CLK line[30] vssd1 vssd1 vccd1 vccd1 _05541_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10619__D line[33] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05471_ _05471_/A _05494_/Y vssd1 vssd1 vccd1 vccd1 _13871_/Z sky130_fd_sc_hd__ebufn_2
X_07210_ _07240_/CLK line[16] vssd1 vssd1 vccd1 vccd1 _07211_/A sky130_fd_sc_hd__dfxtp_1
X_08190_ _08220_/CLK line[80] vssd1 vssd1 vccd1 vccd1 _08191_/A sky130_fd_sc_hd__dfxtp_1
X_07141_ _07141_/A _07174_/Y vssd1 vssd1 vccd1 vccd1 _13861_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[5\].V OVHB\[5\].V/CLK TIE/HI rst_n vssd1 vssd1 vccd1 vccd1 OVHB\[5\].V/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12834__D line[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[14\].VALID\[8\].TOBUF OVHB\[14\].VALID\[8\].FF/Q OVHB\[14\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04931_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__07928__D line[83] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07072_ _07100_/CLK line[90] vssd1 vssd1 vccd1 vccd1 _07073_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_145_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[8\].VALID\[3\].FF_D A[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06023_ _06023_/A _06054_/Y vssd1 vssd1 vccd1 vccd1 _13863_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_126_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XOVHB\[9\].VALID\[4\].FF OVHB\[9\].V/CLK A[11] vssd1 vssd1 vccd1 vccd1 OVHB\[9\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_114_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07974_ _07974_/A _07979_/Y vssd1 vssd1 vccd1 vccd1 _13854_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_19_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09713_ _09725_/CLK line[3] vssd1 vssd1 vccd1 vccd1 _09714_/A sky130_fd_sc_hd__dfxtp_1
X_06925_ _06925_/CLK line[9] vssd1 vssd1 vccd1 vccd1 _06926_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11185__D line[36] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09644_ _09644_/A _09659_/Y vssd1 vssd1 vccd1 vccd1 _13844_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06279__D line[97] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06856_ _06856_/A _06859_/Y vssd1 vssd1 vccd1 vccd1 _13856_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[9\].VALID\[12\].TOBUF OVHB\[9\].VALID\[12\].FF/Q OVHB\[9\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04929_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_35_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05807_ _05807_/CLK _05808_/X vssd1 vssd1 vccd1 vccd1 _05805_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_82_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09575_ _09585_/CLK line[68] vssd1 vssd1 vccd1 vccd1 _09576_/A sky130_fd_sc_hd__dfxtp_1
X_06787_ _06787_/CLK _06788_/X vssd1 vssd1 vccd1 vccd1 _06785_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__08494__D line[86] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08526_ _08526_/A _08539_/Y vssd1 vssd1 vccd1 vccd1 _13846_/Z sky130_fd_sc_hd__ebufn_2
XPHY_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05738_ _13901_/X wr vssd1 vssd1 vccd1 vccd1 _05738_/X sky130_fd_sc_hd__and2_1
XANTENNA__04930__B2 _04930_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08457_ _08465_/CLK line[69] vssd1 vssd1 vccd1 vccd1 _08458_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05669_ _13901_/X vssd1 vssd1 vccd1 vccd1 _05669_/Y sky130_fd_sc_hd__inv_2
XPHY_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07408_ _07408_/A _07419_/Y vssd1 vssd1 vccd1 vccd1 _13848_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_50_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08388_ _08388_/A _08399_/Y vssd1 vssd1 vccd1 vccd1 _13708_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07339_ _07345_/CLK line[70] vssd1 vssd1 vccd1 vccd1 _07340_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12744__D line[123] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06742__D line[53] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10350_ _10350_/A _10359_/Y vssd1 vssd1 vccd1 vccd1 _13710_/Z sky130_fd_sc_hd__ebufn_2
X_09009_ _09025_/CLK line[65] vssd1 vssd1 vccd1 vccd1 _09010_/A sky130_fd_sc_hd__dfxtp_1
X_10281_ _10285_/CLK line[7] vssd1 vssd1 vccd1 vccd1 _10282_/A sky130_fd_sc_hd__dfxtp_1
X_12020_ _12020_/A _12039_/Y vssd1 vssd1 vccd1 vccd1 _13700_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XOVHB\[2\].VALID\[11\].TOBUF OVHB\[2\].VALID\[11\].FF/Q OVHB\[2\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04915_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_183_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13575__D line[105] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08669__D line[38] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[20\].VALID\[7\].TOBUF OVHB\[20\].VALID\[7\].FF/Q OVHB\[20\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/A2 sky130_fd_sc_hd__ebufn_2
X_13971_ _13971_/A _13971_/B _13971_/C _13971_/D vssd1 vssd1 vccd1 vccd1 _13971_/X
+ sky130_fd_sc_hd__and4_4
XANTENNA__11095__D line[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[7\].VALID\[6\].FF OVHB\[7\].V/CLK A[13] vssd1 vssd1 vccd1 vccd1 OVHB\[7\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_86_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12922_ _12922_/A _12949_/Y vssd1 vssd1 vccd1 vccd1 _13762_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[18\].VALID\[12\].FF_D A[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05093__D line[67] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12919__D line[75] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12853_ _12875_/CLK line[45] vssd1 vssd1 vccd1 vccd1 _12854_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_33_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10289__A _13923_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11823__D line[72] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11804_ _11804_/A _11829_/Y vssd1 vssd1 vccd1 vccd1 _13764_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_33_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06917__D line[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12784_ _12784_/A _12809_/Y vssd1 vssd1 vccd1 vccd1 _13624_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__04921__B2 _04923_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11735_ _11755_/CLK line[46] vssd1 vssd1 vccd1 vccd1 _11736_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11666_ _11666_/A _11689_/Y vssd1 vssd1 vccd1 vccd1 _13626_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13405_ _13435_/CLK line[32] vssd1 vssd1 vccd1 vccd1 _13406_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_186_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10617_ _10635_/CLK line[47] vssd1 vssd1 vccd1 vccd1 _10618_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_174_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_OVHB\[28\].VALID\[11\].FF_D A[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11597_ _11615_/CLK line[111] vssd1 vssd1 vccd1 vccd1 _11598_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[18\].CGAND_B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13336_ _13336_/A _13369_/Y vssd1 vssd1 vccd1 vccd1 _13616_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06652__D line[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10548_ _10548_/A _10569_/Y vssd1 vssd1 vccd1 vccd1 _13628_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10174__D line[86] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13267_ _13295_/CLK line[106] vssd1 vssd1 vccd1 vccd1 _13268_/A sky130_fd_sc_hd__dfxtp_1
X_10479_ _10495_/CLK line[97] vssd1 vssd1 vccd1 vccd1 _10480_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05268__D line[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12218_ _12218_/A _12249_/Y vssd1 vssd1 vccd1 vccd1 _13618_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_170_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_DATA\[21\].CLKBUF\[3\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13198_ _13198_/A _13229_/Y vssd1 vssd1 vccd1 vccd1 _13758_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13485__D line[78] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12149_ _12175_/CLK line[107] vssd1 vssd1 vccd1 vccd1 _12150_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08579__D line[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07483__D line[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_04971_ _04971_/A _05004_/Y vssd1 vssd1 vccd1 vccd1 _13651_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11583__A _13926_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06710_ _06710_/A _06719_/Y vssd1 vssd1 vccd1 vccd1 _13710_/Z sky130_fd_sc_hd__ebufn_2
X_07690_ _07690_/A _07699_/Y vssd1 vssd1 vccd1 vccd1 _13850_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_92_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XOVHB\[10\].V OVHB\[10\].V/CLK TIE/HI rst_n vssd1 vssd1 vccd1 vccd1 OVHB\[10\].V/Q
+ sky130_fd_sc_hd__dfrtp_1
X_06641_ _06645_/CLK line[7] vssd1 vssd1 vccd1 vccd1 _06642_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11733__D line[45] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09360_ _09360_/A _09379_/Y vssd1 vssd1 vccd1 vccd1 _13840_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06827__D line[106] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06572_ _06572_/A _06579_/Y vssd1 vssd1 vccd1 vccd1 _13852_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05731__D line[103] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08311_ _08325_/CLK line[2] vssd1 vssd1 vccd1 vccd1 _08312_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[5\].VALID\[8\].FF OVHB\[5\].V/CLK A[15] vssd1 vssd1 vccd1 vccd1 OVHB\[5\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_05523_ _05525_/CLK line[8] vssd1 vssd1 vccd1 vccd1 _05524_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10349__D line[38] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09291_ _09305_/CLK line[66] vssd1 vssd1 vccd1 vccd1 _09292_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_178_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05454_ _05454_/A _05459_/Y vssd1 vssd1 vccd1 vccd1 _13854_/Z sky130_fd_sc_hd__ebufn_2
X_08242_ _08242_/A _08259_/Y vssd1 vssd1 vccd1 vccd1 _13842_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_193_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05385_ _05385_/CLK line[73] vssd1 vssd1 vccd1 vccd1 _05386_/A sky130_fd_sc_hd__dfxtp_1
X_08173_ _08185_/CLK line[67] vssd1 vssd1 vccd1 vccd1 _08174_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[29\].VALID\[2\].TOBUF OVHB\[29\].VALID\[2\].FF/Q OVHB\[29\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04930_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__07658__D line[88] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07124_ _07124_/A _07139_/Y vssd1 vssd1 vccd1 vccd1 _13844_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_118_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10084__D line[59] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07055_ _07065_/CLK line[68] vssd1 vssd1 vccd1 vccd1 _07056_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11758__A _13927_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06006_ _06006_/A _06019_/Y vssd1 vssd1 vccd1 vccd1 _13846_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[30\].VALID\[7\].FF_D A[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11908__D line[125] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[23\].VALID\[11\].FF OVHB\[23\].V/CLK A[18] vssd1 vssd1 vccd1 vccd1 OVHB\[23\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13973__A A_h[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07393__D line[109] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05906__D line[55] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[25\].VALID\[13\].TOBUF OVHB\[25\].VALID\[13\].FF/Q OVHB\[25\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04916_/B2 sky130_fd_sc_hd__ebufn_2
X_07957_ _07975_/CLK line[111] vssd1 vssd1 vccd1 vccd1 _07958_/A sky130_fd_sc_hd__dfxtp_1
X_06908_ _06908_/A _06929_/Y vssd1 vssd1 vccd1 vccd1 _13628_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_101_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07888_ _07888_/A _07909_/Y vssd1 vssd1 vccd1 vccd1 _13768_/Z sky130_fd_sc_hd__ebufn_2
X_09627_ _09655_/CLK line[106] vssd1 vssd1 vccd1 vccd1 _09628_/A sky130_fd_sc_hd__dfxtp_1
X_06839_ _06855_/CLK line[97] vssd1 vssd1 vccd1 vccd1 _06840_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_15_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09558_ _09558_/A _09589_/Y vssd1 vssd1 vccd1 vccd1 _13758_/Z sky130_fd_sc_hd__ebufn_2
XPHY_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05641__D line[76] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10259__D line[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08509_ _08535_/CLK line[107] vssd1 vssd1 vccd1 vccd1 _08510_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_196_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09489_ _09515_/CLK line[43] vssd1 vssd1 vccd1 vccd1 _09490_/A sky130_fd_sc_hd__dfxtp_1
XPHY_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11520_ _11520_/A _11549_/Y vssd1 vssd1 vccd1 vccd1 _13760_/Z sky130_fd_sc_hd__ebufn_2
XPHY_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12474__D line[113] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11451_ _11475_/CLK line[44] vssd1 vssd1 vccd1 vccd1 _11452_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_168_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[13\].VALID\[13\].FF OVHB\[13\].V/CLK A[20] vssd1 vssd1 vccd1 vccd1 OVHB\[13\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07568__D line[61] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10402_ _10402_/A _10429_/Y vssd1 vssd1 vccd1 vccd1 _13762_/Z sky130_fd_sc_hd__ebufn_2
X_11382_ _11382_/A _11409_/Y vssd1 vssd1 vccd1 vccd1 _13622_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_124_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13121_ _13121_/A _13124_/Y vssd1 vssd1 vccd1 vccd1 _13681_/Z sky130_fd_sc_hd__ebufn_2
X_10333_ _10355_/CLK line[45] vssd1 vssd1 vccd1 vccd1 _10334_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_125_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09783__D line[35] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13052_ _13052_/CLK _13053_/X vssd1 vssd1 vccd1 vccd1 _13050_/CLK sky130_fd_sc_hd__dlclkp_1
X_10264_ _10264_/A _10289_/Y vssd1 vssd1 vccd1 vccd1 _13624_/Z sky130_fd_sc_hd__ebufn_2
X_12003_ _13934_/X wr vssd1 vssd1 vccd1 vccd1 _12003_/X sky130_fd_sc_hd__and2_1
XANTENNA__10722__D line[95] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10195_ _10215_/CLK line[110] vssd1 vssd1 vccd1 vccd1 _10196_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05816__D line[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13954_ _13960_/C _13960_/B _13960_/A _13960_/D vssd1 vssd1 vccd1 vccd1 _13954_/X
+ sky130_fd_sc_hd__and4bb_4
X_12905_ _12905_/A _12914_/Y vssd1 vssd1 vccd1 vccd1 _13745_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12649__D line[65] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13885_ _13885_/A _13894_/Y vssd1 vssd1 vccd1 vccd1 _13885_/Z sky130_fd_sc_hd__ebufn_2
X_12836_ _12840_/CLK line[23] vssd1 vssd1 vccd1 vccd1 _12837_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09023__D line[72] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12767_ _12767_/A _12774_/Y vssd1 vssd1 vccd1 vccd1 _13887_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09958__D line[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13123__A _13938_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11718_ _11720_/CLK line[24] vssd1 vssd1 vccd1 vccd1 _11719_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[14\].VALID\[0\].FF OVHB\[14\].V/CLK A[7] vssd1 vssd1 vccd1 vccd1 OVHB\[14\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_12698_ _12700_/CLK line[88] vssd1 vssd1 vccd1 vccd1 _12699_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_30_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[4\].VALID\[6\].FF_D A[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11649_ _11649_/A _11654_/Y vssd1 vssd1 vccd1 vccd1 _13889_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_175_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[31\].VALID\[4\].FF OVHB\[31\].V/CLK A[11] vssd1 vssd1 vccd1 vccd1 OVHB\[31\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_05170_ _05170_/A _05179_/Y vssd1 vssd1 vccd1 vccd1 _13850_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06382__D line[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13319_ _13319_/A _13334_/Y vssd1 vssd1 vccd1 vccd1 _13879_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_170_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08860_ _08860_/A _08889_/Y vssd1 vssd1 vccd1 vccd1 _13620_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_97_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07811_ _07835_/CLK line[44] vssd1 vssd1 vccd1 vccd1 _07812_/A sky130_fd_sc_hd__dfxtp_1
X_08791_ _08815_/CLK line[108] vssd1 vssd1 vccd1 vccd1 _08792_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_84_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XOVHB\[2\].VALID\[4\].TOBUF OVHB\[2\].VALID\[4\].FF/Q OVHB\[2\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04925_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07742_ _07742_/A _07769_/Y vssd1 vssd1 vccd1 vccd1 _13622_/Z sky130_fd_sc_hd__ebufn_2
X_04954_ _04954_/A _04969_/Y vssd1 vssd1 vccd1 vccd1 _13634_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[27\].VALID\[7\].TOBUF OVHB\[27\].VALID\[7\].FF/Q OVHB\[27\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/A2 sky130_fd_sc_hd__ebufn_2
XFILLER_203_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07673_ _07695_/CLK line[109] vssd1 vssd1 vccd1 vccd1 _07674_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11463__D line[35] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09412_ _09412_/CLK _09413_/X vssd1 vssd1 vccd1 vccd1 _09410_/CLK sky130_fd_sc_hd__dlclkp_1
X_06624_ _06624_/A _06649_/Y vssd1 vssd1 vccd1 vccd1 _13624_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06557__D line[111] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09343_ _13916_/X wr vssd1 vssd1 vccd1 vccd1 _09343_/X sky130_fd_sc_hd__and2_1
X_06555_ _06575_/CLK line[110] vssd1 vssd1 vccd1 vccd1 _06556_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_80_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05506_ _05506_/A _05529_/Y vssd1 vssd1 vccd1 vccd1 _13626_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08772__D line[85] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09274_ _13916_/X vssd1 vssd1 vccd1 vccd1 _09274_/Y sky130_fd_sc_hd__inv_2
XFILLER_178_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06486_ _06486_/A _06509_/Y vssd1 vssd1 vccd1 vccd1 _13766_/Z sky130_fd_sc_hd__ebufn_2
X_08225_ _08255_/CLK line[96] vssd1 vssd1 vccd1 vccd1 _08226_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[11\].CGAND _13901_/X wr vssd1 vssd1 vccd1 vccd1 OVHB\[11\].CGAND/X sky130_fd_sc_hd__and2_4
X_05437_ _05455_/CLK line[111] vssd1 vssd1 vccd1 vccd1 _05438_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_165_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05368_ _05368_/A _05389_/Y vssd1 vssd1 vccd1 vccd1 _13768_/Z sky130_fd_sc_hd__ebufn_2
X_08156_ _08156_/A _08189_/Y vssd1 vssd1 vccd1 vccd1 _13756_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_180_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07107_ _07135_/CLK line[106] vssd1 vssd1 vccd1 vccd1 _07108_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_106_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05299_ _05315_/CLK line[33] vssd1 vssd1 vccd1 vccd1 _05300_/A sky130_fd_sc_hd__dfxtp_1
X_08087_ _08115_/CLK line[42] vssd1 vssd1 vccd1 vccd1 _08088_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_134_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XOVHB\[12\].VALID\[2\].FF OVHB\[12\].V/CLK A[9] vssd1 vssd1 vccd1 vccd1 OVHB\[12\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_164_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07038_ _07038_/A _07069_/Y vssd1 vssd1 vccd1 vccd1 _13758_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_134_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11638__D line[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[19\].VALID\[3\].FF_D A[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09108__D line[125] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08989_ _08989_/A _08994_/Y vssd1 vssd1 vccd1 vccd1 _13749_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13853__D line[104] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08947__D line[37] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10951_ _10951_/A _10954_/Y vssd1 vssd1 vccd1 vccd1 _13751_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_56_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13670_ _13680_/CLK line[20] vssd1 vssd1 vccd1 vccd1 _13671_/A sky130_fd_sc_hd__dfxtp_1
X_10882_ _10882_/CLK _10883_/X vssd1 vssd1 vccd1 vccd1 _10880_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__05371__D line[66] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12621_ _12621_/A _12634_/Y vssd1 vssd1 vccd1 vccd1 _13741_/Z sky130_fd_sc_hd__ebufn_2
XPHY_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12552_ _12560_/CLK line[21] vssd1 vssd1 vccd1 vccd1 _12553_/A sky130_fd_sc_hd__dfxtp_1
XPHY_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08682__D line[58] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11503_ _11503_/A _11514_/Y vssd1 vssd1 vccd1 vccd1 _13743_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12483_ _12483_/A _12494_/Y vssd1 vssd1 vccd1 vccd1 _13883_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07298__D line[51] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11434_ _11440_/CLK line[22] vssd1 vssd1 vccd1 vccd1 _11435_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_165_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11365_ _11365_/A _11374_/Y vssd1 vssd1 vccd1 vccd1 _13885_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_98_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13104_ _13120_/CLK line[17] vssd1 vssd1 vccd1 vccd1 _13105_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_98_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06930__D line[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10316_ _10320_/CLK line[23] vssd1 vssd1 vccd1 vccd1 _10317_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_98_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XOVHB\[28\].VALID\[7\].FF OVHB\[28\].V/CLK A[14] vssd1 vssd1 vccd1 vccd1 OVHB\[28\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_125_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11296_ _11300_/CLK line[87] vssd1 vssd1 vccd1 vccd1 _11297_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10452__D line[85] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13035_ _13035_/A _13054_/Y vssd1 vssd1 vccd1 vccd1 _13875_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_3_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10247_ _10247_/A _10254_/Y vssd1 vssd1 vccd1 vccd1 _13887_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_121_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05546__D line[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10178_ _10180_/CLK line[88] vssd1 vssd1 vccd1 vccd1 _10179_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13763__D line[77] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[18\].CLKBUF\[6\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05843__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08857__D line[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[10\].VALID\[4\].FF OVHB\[10\].V/CLK A[11] vssd1 vssd1 vccd1 vccd1 OVHB\[10\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_82_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07761__D line[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12379__D line[70] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13937_ _13938_/A _13938_/B _13938_/C _13938_/D vssd1 vssd1 vccd1 vccd1 _13937_/X
+ sky130_fd_sc_hd__and4b_4
XFILLER_34_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13868_ _13890_/CLK line[125] vssd1 vssd1 vccd1 vccd1 _13869_/A sky130_fd_sc_hd__dfxtp_1
X_12819_ _12819_/A _12844_/Y vssd1 vssd1 vccd1 vccd1 _13659_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_62_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13799_ _13799_/A _13824_/Y vssd1 vssd1 vccd1 vccd1 _13799_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09688__D line[120] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06340_ _06340_/A _06369_/Y vssd1 vssd1 vccd1 vccd1 _13620_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_203_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13788__A _13899_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10627__D line[37] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06271_ _06295_/CLK line[108] vssd1 vssd1 vccd1 vccd1 _06272_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_30_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XDATA\[29\].CLKBUF\[2\] clk vssd1 vssd1 vccd1 vccd1 _10917_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__13003__D line[99] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[0\].VALID\[9\].TOBUF OVHB\[0\].VALID\[9\].FF/Q OVHB\[0\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04914_/B2 sky130_fd_sc_hd__ebufn_2
X_05222_ _05222_/A _05249_/Y vssd1 vssd1 vccd1 vccd1 _13622_/Z sky130_fd_sc_hd__ebufn_2
X_08010_ _08010_/CLK line[121] vssd1 vssd1 vccd1 vccd1 _08011_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_190_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05153_ _05175_/CLK line[109] vssd1 vssd1 vccd1 vccd1 _05154_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07936__D line[87] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09961_ _09961_/A _09974_/Y vssd1 vssd1 vccd1 vccd1 _13881_/Z sky130_fd_sc_hd__ebufn_2
X_05084_ _05084_/A _05109_/Y vssd1 vssd1 vccd1 vccd1 _13764_/Z sky130_fd_sc_hd__ebufn_2
X_08912_ _08920_/CLK line[21] vssd1 vssd1 vccd1 vccd1 _08913_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10362__D line[58] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09892_ _09900_/CLK line[85] vssd1 vssd1 vccd1 vccd1 _09893_/A sky130_fd_sc_hd__dfxtp_1
X_08843_ _08843_/A _08854_/Y vssd1 vssd1 vccd1 vccd1 _13883_/Z sky130_fd_sc_hd__ebufn_2
X_08774_ _08780_/CLK line[86] vssd1 vssd1 vccd1 vccd1 _08775_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_27_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05986_ _05986_/A _06019_/Y vssd1 vssd1 vccd1 vccd1 _13826_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07671__D line[108] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[26\].VALID\[9\].FF OVHB\[26\].V/CLK A[16] vssd1 vssd1 vccd1 vccd1 OVHB\[26\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12289__D line[43] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07725_ _07725_/A _07734_/Y vssd1 vssd1 vccd1 vccd1 _13885_/Z sky130_fd_sc_hd__ebufn_2
X_04937_ _04965_/CLK line[10] vssd1 vssd1 vccd1 vccd1 _04938_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11193__D line[40] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06287__D line[101] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07656_ _07660_/CLK line[87] vssd1 vssd1 vccd1 vccd1 _07657_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[5\].VOBUF OVHB\[5\].V/Q OVHB\[5\].INV/Y vssd1 vssd1 vccd1 vccd1 _04912_/B1
+ sky130_fd_sc_hd__ebufn_2
XFILLER_43_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06607_ _06607_/A _06614_/Y vssd1 vssd1 vccd1 vccd1 _13887_/Z sky130_fd_sc_hd__ebufn_2
X_07587_ _07587_/A _07594_/Y vssd1 vssd1 vccd1 vccd1 _13747_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_179_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09598__D line[93] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09326_ _09340_/CLK line[82] vssd1 vssd1 vccd1 vccd1 _09327_/A sky130_fd_sc_hd__dfxtp_1
X_06538_ _06540_/CLK line[88] vssd1 vssd1 vccd1 vccd1 _06539_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10537__D line[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09257_ _09257_/A _09274_/Y vssd1 vssd1 vccd1 vccd1 _13737_/Z sky130_fd_sc_hd__ebufn_2
X_06469_ _06469_/A _06474_/Y vssd1 vssd1 vccd1 vccd1 _13749_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__04926__A2_N _04926_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08208_ _08220_/CLK line[83] vssd1 vssd1 vccd1 vccd1 _08209_/A sky130_fd_sc_hd__dfxtp_1
X_09188_ _09200_/CLK line[19] vssd1 vssd1 vccd1 vccd1 _09189_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_193_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08139_ _08139_/A _08154_/Y vssd1 vssd1 vccd1 vccd1 _13739_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12752__D line[127] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07846__D line[60] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11150_ _11160_/CLK line[20] vssd1 vssd1 vccd1 vccd1 _11151_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06750__D line[57] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11368__D line[120] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10101_ _10101_/A _10114_/Y vssd1 vssd1 vccd1 vccd1 _13741_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_108_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11081_ _11081_/A _11094_/Y vssd1 vssd1 vccd1 vccd1 _13881_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[18\].CLKBUF\[5\] clk vssd1 vssd1 vccd1 vccd1 _07662_/CLK sky130_fd_sc_hd__clkbuf_4
XOVHB\[15\].VALID\[11\].TOBUF OVHB\[15\].VALID\[11\].FF/Q OVHB\[15\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04915_/B2 sky130_fd_sc_hd__ebufn_2
X_10032_ _10040_/CLK line[21] vssd1 vssd1 vccd1 vccd1 _10033_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_102_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11983_ _11983_/A _12004_/Y vssd1 vssd1 vccd1 vccd1 _13663_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_90_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[9\].VALID\[4\].TOBUF OVHB\[9\].VALID\[4\].FF/Q OVHB\[9\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04925_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_16_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13722_ _13750_/CLK line[58] vssd1 vssd1 vccd1 vccd1 _13723_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06197__D line[74] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10934_ _10950_/CLK line[49] vssd1 vssd1 vccd1 vccd1 _10935_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_189_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13653_ _13653_/A _13684_/Y vssd1 vssd1 vccd1 vccd1 _13653_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12927__D line[79] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10865_ _10865_/A _10884_/Y vssd1 vssd1 vccd1 vccd1 _13665_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[0\].VALID\[9\].FF_D A[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12604_ _12630_/CLK line[59] vssd1 vssd1 vccd1 vccd1 _12605_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06925__D line[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XOVHB\[4\].VALID\[13\].FF OVHB\[4\].V/CLK A[20] vssd1 vssd1 vccd1 vccd1 OVHB\[4\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_13584_ _13610_/CLK line[123] vssd1 vssd1 vccd1 vccd1 _13585_/A sky130_fd_sc_hd__dfxtp_1
X_10796_ _10810_/CLK line[114] vssd1 vssd1 vccd1 vccd1 _10797_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09301__D line[71] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12535_ _12535_/A _12564_/Y vssd1 vssd1 vccd1 vccd1 _13655_/Z sky130_fd_sc_hd__ebufn_2
XPHY_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12466_ _12490_/CLK line[124] vssd1 vssd1 vccd1 vccd1 _12467_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_138_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11417_ _11417_/A _11444_/Y vssd1 vssd1 vccd1 vccd1 _13657_/Z sky130_fd_sc_hd__ebufn_2
X_12397_ _12397_/A _12424_/Y vssd1 vssd1 vccd1 vccd1 _13797_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06660__D line[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11348_ _11370_/CLK line[125] vssd1 vssd1 vccd1 vccd1 _11349_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_99_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11278__D line[93] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11279_ _11279_/A _11304_/Y vssd1 vssd1 vccd1 vccd1 _13799_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05276__D line[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13018_ _13937_/X wr vssd1 vssd1 vccd1 vccd1 _13018_/X sky130_fd_sc_hd__and2_1
XANTENNA__13493__D line[67] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05840_ _05840_/CLK line[25] vssd1 vssd1 vccd1 vccd1 _05841_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08587__D line[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XDATA\[17\].CLKBUF\[2\] clk vssd1 vssd1 vccd1 vccd1 _07277_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_82_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05771_ _05771_/A _05774_/Y vssd1 vssd1 vccd1 vccd1 _13891_/Z sky130_fd_sc_hd__ebufn_2
X_07510_ _07520_/CLK line[20] vssd1 vssd1 vccd1 vccd1 _07511_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_63_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08490_ _08500_/CLK line[84] vssd1 vssd1 vccd1 vccd1 _08491_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_23_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07441_ _07441_/A _07454_/Y vssd1 vssd1 vccd1 vccd1 _13881_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11741__D line[34] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06835__D line[110] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07372_ _07380_/CLK line[85] vssd1 vssd1 vccd1 vccd1 _07373_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_188_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09211__D line[44] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[22\].VALID\[2\].FF_D A[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09111_ _09111_/A _09134_/Y vssd1 vssd1 vccd1 vccd1 _13871_/Z sky130_fd_sc_hd__ebufn_2
X_06323_ _06323_/A _06334_/Y vssd1 vssd1 vccd1 vccd1 _13883_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_175_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09042_ _09060_/CLK line[95] vssd1 vssd1 vccd1 vccd1 _09043_/A sky130_fd_sc_hd__dfxtp_1
X_06254_ _06260_/CLK line[86] vssd1 vssd1 vccd1 vccd1 _06255_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[28\].VALID\[11\].FF OVHB\[28\].V/CLK A[18] vssd1 vssd1 vccd1 vccd1 OVHB\[28\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_135_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13668__D line[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05205_ _05205_/A _05214_/Y vssd1 vssd1 vccd1 vccd1 _13885_/Z sky130_fd_sc_hd__ebufn_2
X_06185_ _06185_/A _06194_/Y vssd1 vssd1 vccd1 vccd1 _13745_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_190_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_OVHB\[15\].VALID\[6\].FF_D A[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05136_ _05140_/CLK line[87] vssd1 vssd1 vccd1 vccd1 _05137_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_144_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10092__D line[63] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09944_ _09970_/CLK line[123] vssd1 vssd1 vccd1 vccd1 _09945_/A sky130_fd_sc_hd__dfxtp_1
X_05067_ _05067_/A _05074_/Y vssd1 vssd1 vccd1 vccd1 _13747_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05186__D line[124] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09875_ _09875_/A _09904_/Y vssd1 vssd1 vccd1 vccd1 _13795_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_112_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11916__D line[114] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08826_ _08850_/CLK line[124] vssd1 vssd1 vccd1 vccd1 _08827_/A sky130_fd_sc_hd__dfxtp_1
X_08757_ _08757_/A _08784_/Y vssd1 vssd1 vccd1 vccd1 _13797_/Z sky130_fd_sc_hd__ebufn_2
X_05969_ _05969_/A _05984_/Y vssd1 vssd1 vccd1 vccd1 _13809_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_38_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07708_ _07730_/CLK line[125] vssd1 vssd1 vccd1 vccd1 _07709_/A sky130_fd_sc_hd__dfxtp_1
X_08688_ _08710_/CLK line[61] vssd1 vssd1 vccd1 vccd1 _08689_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[31\].CLKBUF\[1\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[18\].VALID\[13\].FF OVHB\[18\].V/CLK A[20] vssd1 vssd1 vccd1 vccd1 OVHB\[18\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_07639_ _07639_/A _07664_/Y vssd1 vssd1 vccd1 vccd1 _13799_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_202_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10650_ _10670_/CLK line[62] vssd1 vssd1 vccd1 vccd1 _10651_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_167_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05004__A _13931_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09309_ _13916_/X vssd1 vssd1 vccd1 vccd1 _09309_/Y sky130_fd_sc_hd__inv_2
XANTENNA__10267__D line[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10581_ _10581_/A _10604_/Y vssd1 vssd1 vccd1 vccd1 _13661_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[16\].V_RESET_B rst_n vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12320_ _12350_/CLK line[48] vssd1 vssd1 vccd1 vccd1 _12321_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08960__D line[48] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12251_ _12251_/A _12284_/Y vssd1 vssd1 vccd1 vccd1 _13651_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_119_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12482__D line[117] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07576__D line[50] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[7\].VALID\[9\].TOBUF OVHB\[7\].VALID\[9\].FF/Q OVHB\[7\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04914_/B2 sky130_fd_sc_hd__ebufn_2
X_11202_ _11230_/CLK line[58] vssd1 vssd1 vccd1 vccd1 _11203_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[5\].VALID\[11\].FF_D A[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12182_ _12210_/CLK line[122] vssd1 vssd1 vccd1 vccd1 _12183_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.M\[3\].MUX\[0\]_A1 _13749_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11133_ _11133_/A _11164_/Y vssd1 vssd1 vccd1 vccd1 _13653_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07873__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09791__D line[39] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11064_ _11090_/CLK line[123] vssd1 vssd1 vccd1 vccd1 _11065_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_95_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10730__D line[84] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10015_ _10015_/A _10044_/Y vssd1 vssd1 vccd1 vccd1 _13655_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_48_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05824__D line[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08200__D line[94] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_DEC.DEC0.AND3_A A[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11966_ _11966_/A _11969_/Y vssd1 vssd1 vccd1 vccd1 _13646_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_44_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13705_ _13715_/CLK line[36] vssd1 vssd1 vccd1 vccd1 _13706_/A sky130_fd_sc_hd__dfxtp_1
X_10917_ _10917_/CLK _10918_/X vssd1 vssd1 vccd1 vccd1 _10915_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__12657__D line[69] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11897_ _11897_/CLK _11898_/X vssd1 vssd1 vccd1 vccd1 _11895_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_71_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13636_ _13636_/A _13649_/Y vssd1 vssd1 vccd1 vccd1 _13636_/Z sky130_fd_sc_hd__ebufn_2
X_10848_ _13925_/X wr vssd1 vssd1 vccd1 vccd1 _10848_/X sky130_fd_sc_hd__and2_1
X_13567_ _13575_/CLK line[101] vssd1 vssd1 vccd1 vccd1 _13568_/A sky130_fd_sc_hd__dfxtp_1
X_10779_ _13924_/X vssd1 vssd1 vccd1 vccd1 _10779_/Y sky130_fd_sc_hd__inv_2
XANTENNA__09966__D line[119] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12518_ _12518_/A _12529_/Y vssd1 vssd1 vccd1 vccd1 _13638_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_117_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13498_ _13498_/A _13509_/Y vssd1 vssd1 vccd1 vccd1 _13778_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[28\].VALID\[6\].FF_D A[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12392__D line[90] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10905__D line[36] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12449_ _12455_/CLK line[102] vssd1 vssd1 vccd1 vccd1 _12450_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_145_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06390__D line[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07990_ _08010_/CLK line[126] vssd1 vssd1 vccd1 vccd1 _07991_/A sky130_fd_sc_hd__dfxtp_1
X_06941_ _06941_/A _06964_/Y vssd1 vssd1 vccd1 vccd1 _13661_/Z sky130_fd_sc_hd__ebufn_2
XMUX.M\[1\].MUX\[1\] _13646_/Z _13716_/Z _13786_/Z _13856_/Z MUX.SEL0BUF\[1\]/X MUX.SEL1BUF\[1\]/X
+ vssd1 vssd1 vccd1 vccd1 Do[9] sky130_fd_sc_hd__mux4_1
XANTENNA__10640__D line[48] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09660_ _09690_/CLK line[112] vssd1 vssd1 vccd1 vccd1 _09661_/A sky130_fd_sc_hd__dfxtp_1
X_06872_ _06890_/CLK line[127] vssd1 vssd1 vccd1 vccd1 _06873_/A sky130_fd_sc_hd__dfxtp_1
X_08611_ _08611_/A _08644_/Y vssd1 vssd1 vccd1 vccd1 _13651_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[14\].VALID\[4\].TOBUF OVHB\[14\].VALID\[4\].FF/Q OVHB\[14\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04925_/B2 sky130_fd_sc_hd__ebufn_2
XOVHB\[0\].VALID\[11\].FF OVHB\[0\].V/CLK A[18] vssd1 vssd1 vccd1 vccd1 OVHB\[0\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_05823_ _05823_/A _05844_/Y vssd1 vssd1 vccd1 vccd1 _13663_/Z sky130_fd_sc_hd__ebufn_2
X_09591_ _09591_/A _09624_/Y vssd1 vssd1 vccd1 vccd1 _13791_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_36_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08542_ _08570_/CLK line[122] vssd1 vssd1 vccd1 vccd1 _08543_/A sky130_fd_sc_hd__dfxtp_1
X_05754_ _05770_/CLK line[113] vssd1 vssd1 vccd1 vccd1 _05755_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_211_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12567__D line[42] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08473_ _08473_/A _08504_/Y vssd1 vssd1 vccd1 vccd1 _13793_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11471__D line[39] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05685_ _05685_/A _05704_/Y vssd1 vssd1 vccd1 vccd1 _13805_/Z sky130_fd_sc_hd__ebufn_2
X_07424_ _07450_/CLK line[123] vssd1 vssd1 vccd1 vccd1 _07425_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06565__D line[100] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07355_ _07355_/A _07384_/Y vssd1 vssd1 vccd1 vccd1 _13795_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_148_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09876__D line[92] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06306_ _06330_/CLK line[124] vssd1 vssd1 vccd1 vccd1 _06307_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08780__D line[89] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07286_ _07310_/CLK line[60] vssd1 vssd1 vccd1 vccd1 _07287_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13398__D line[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09025_ _09025_/CLK line[73] vssd1 vssd1 vccd1 vccd1 _09026_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10815__D line[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06237_ _06237_/A _06264_/Y vssd1 vssd1 vccd1 vccd1 _13797_/Z sky130_fd_sc_hd__ebufn_2
X_06168_ _06190_/CLK line[61] vssd1 vssd1 vccd1 vccd1 _06169_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[10\].CLKBUF\[1\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05119_ _05119_/A _05144_/Y vssd1 vssd1 vccd1 vccd1 _13799_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_131_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06099_ _06099_/A _06124_/Y vssd1 vssd1 vccd1 vccd1 _13659_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_49_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05494__A _13900_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09927_ _09935_/CLK line[101] vssd1 vssd1 vccd1 vccd1 _09928_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11646__D line[119] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09858_ _09858_/A _09869_/Y vssd1 vssd1 vccd1 vccd1 _13778_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[17\].CG clk OVHB\[17\].CGAND/X vssd1 vssd1 vccd1 vccd1 OVHB\[17\].V/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA_OVHB\[9\].VALID\[1\].FF_D A[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09116__D line[114] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08809_ _08815_/CLK line[102] vssd1 vssd1 vccd1 vccd1 _08810_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_45_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09789_ _09795_/CLK line[38] vssd1 vssd1 vccd1 vccd1 _09790_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.M\[0\].MUX\[7\]_A3 _13852_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11820_ _11820_/A _11829_/Y vssd1 vssd1 vccd1 vccd1 _13780_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09413__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08955__D line[41] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11751_ _11755_/CLK line[39] vssd1 vssd1 vccd1 vccd1 _11752_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[22\].CG_CLK clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11381__D line[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_DATA\[3\].CLKBUF\[1\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10702_ _10702_/A _10709_/Y vssd1 vssd1 vccd1 vccd1 _13782_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06475__D line[64] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11682_ _11682_/A _11689_/Y vssd1 vssd1 vccd1 vccd1 _13642_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMUX.M\[0\].MUX\[3\] _13634_/Z _13704_/Z _13774_/Z _13844_/Z MUX.SEL0BUF\[0\]/X MUX.SEL1BUF\[0\]/X
+ vssd1 vssd1 vccd1 vccd1 Do[3] sky130_fd_sc_hd__mux4_1
XFILLER_197_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13421_ _13435_/CLK line[34] vssd1 vssd1 vccd1 vccd1 _13422_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10633_ _10635_/CLK line[40] vssd1 vssd1 vccd1 vccd1 _10634_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[20\].VALID\[3\].TOBUF OVHB\[20\].VALID\[3\].FF/Q OVHB\[20\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04919_/B2 sky130_fd_sc_hd__ebufn_2
XPHY_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13352_ _13352_/A _13369_/Y vssd1 vssd1 vccd1 vccd1 _13632_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05669__A _13901_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08690__D line[62] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10564_ _10564_/A _10569_/Y vssd1 vssd1 vccd1 vccd1 _13644_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_155_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12303_ _12315_/CLK line[35] vssd1 vssd1 vccd1 vccd1 _12304_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_6_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13283_ _13295_/CLK line[99] vssd1 vssd1 vccd1 vccd1 _13284_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05388__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10495_ _10495_/CLK line[105] vssd1 vssd1 vccd1 vccd1 _10496_/A sky130_fd_sc_hd__dfxtp_1
X_12234_ _12234_/A _12249_/Y vssd1 vssd1 vccd1 vccd1 _13634_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_146_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12165_ _12175_/CLK line[100] vssd1 vssd1 vccd1 vccd1 _12166_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_122_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11116_ _11116_/A _11129_/Y vssd1 vssd1 vccd1 vccd1 _13636_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_110_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12096_ _12096_/A _12109_/Y vssd1 vssd1 vccd1 vccd1 _13776_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11556__D line[92] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[14\].VALID\[11\].FF OVHB\[14\].V/CLK A[18] vssd1 vssd1 vccd1 vccd1 OVHB\[14\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10460__D line[89] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11047_ _11055_/CLK line[101] vssd1 vssd1 vccd1 vccd1 _11048_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05554__D line[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13771__D line[66] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08865__D line[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12998_ _12998_/A _13019_/Y vssd1 vssd1 vccd1 vccd1 _13838_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_33_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11949_ _11965_/CLK line[1] vssd1 vssd1 vccd1 vccd1 _11950_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_178_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05470_ _05490_/CLK line[126] vssd1 vssd1 vccd1 vccd1 _05471_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06963__A _13909_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13619_ _13645_/CLK line[11] vssd1 vssd1 vccd1 vccd1 _13620_/A sky130_fd_sc_hd__dfxtp_1
X_07140_ _07170_/CLK line[112] vssd1 vssd1 vccd1 vccd1 _07141_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[11\].VALID\[9\].FF_D A[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10635__D line[41] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[12\].VALID\[9\].TOBUF OVHB\[12\].VALID\[9\].FF/Q OVHB\[12\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04914_/B2 sky130_fd_sc_hd__ebufn_2
X_07071_ _07071_/A _07104_/Y vssd1 vssd1 vccd1 vccd1 _13791_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13011__D line[103] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05729__D line[102] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06022_ _06050_/CLK line[122] vssd1 vssd1 vccd1 vccd1 _06023_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08105__D line[36] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[5\].VALID\[13\].TOBUF OVHB\[5\].VALID\[13\].FF/Q OVHB\[5\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04916_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_206_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07973_ _07975_/CLK line[104] vssd1 vssd1 vccd1 vccd1 _07974_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_206_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09712_ _09712_/A _09729_/Y vssd1 vssd1 vccd1 vccd1 _13632_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10370__D line[62] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDATA\[8\].CLKBUF\[6\] clk vssd1 vssd1 vccd1 vccd1 _13577_/CLK sky130_fd_sc_hd__clkbuf_4
X_06924_ _06924_/A _06929_/Y vssd1 vssd1 vccd1 vccd1 _13644_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_19_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05464__D line[123] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09643_ _09655_/CLK line[99] vssd1 vssd1 vccd1 vccd1 _09644_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_27_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06855_ _06855_/CLK line[105] vssd1 vssd1 vccd1 vccd1 _06856_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_67_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05806_ _05806_/A _05809_/Y vssd1 vssd1 vccd1 vccd1 _13646_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_55_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09574_ _09574_/A _09589_/Y vssd1 vssd1 vccd1 vccd1 _13774_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_82_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06786_ _06786_/A _06789_/Y vssd1 vssd1 vccd1 vccd1 _13786_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_35_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07034__A _13909_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08525_ _08535_/CLK line[100] vssd1 vssd1 vccd1 vccd1 _08526_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12297__D line[47] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05737_ _05737_/CLK _05738_/X vssd1 vssd1 vccd1 vccd1 _05735_/CLK sky130_fd_sc_hd__dlclkp_1
XPHY_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06295__D line[105] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08456_ _08456_/A _08469_/Y vssd1 vssd1 vccd1 vccd1 _13776_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_168_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05668_ _13901_/X wr vssd1 vssd1 vccd1 vccd1 _05668_/X sky130_fd_sc_hd__and2_1
XPHY_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07407_ _07415_/CLK line[101] vssd1 vssd1 vccd1 vccd1 _07408_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_23_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08387_ _08395_/CLK line[37] vssd1 vssd1 vccd1 vccd1 _08388_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05599_ _13901_/X vssd1 vssd1 vccd1 vccd1 _05599_/Y sky130_fd_sc_hd__inv_2
XANTENNA_DATA\[28\].CLKBUF\[4\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07338_ _07338_/A _07349_/Y vssd1 vssd1 vccd1 vccd1 _13778_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_192_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09059__TE_B _09064_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10545__D line[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07269_ _07275_/CLK line[38] vssd1 vssd1 vccd1 vccd1 _07270_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05639__D line[75] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09008_ _09008_/A _09029_/Y vssd1 vssd1 vccd1 vccd1 _13768_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08015__D line[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10280_ _10280_/A _10289_/Y vssd1 vssd1 vccd1 vccd1 _13640_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_164_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12760__D line[116] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07854__D line[49] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07209__A _13910_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13970_ _13971_/A _13971_/B _13971_/C _13971_/D vssd1 vssd1 vccd1 vccd1 _13970_/X
+ sky130_fd_sc_hd__and4b_4
XFILLER_59_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12921_ _12945_/CLK line[76] vssd1 vssd1 vccd1 vccd1 _12922_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_86_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XOVHB\[9\].VALID\[13\].FF OVHB\[9\].V/CLK A[20] vssd1 vssd1 vccd1 vccd1 OVHB\[9\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[31\].VALID\[5\].FF_D A[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12852_ _12852_/A _12879_/Y vssd1 vssd1 vccd1 vccd1 _13692_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[22\].VALID\[0\].FF OVHB\[22\].V/CLK A[7] vssd1 vssd1 vccd1 vccd1 OVHB\[22\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XDATA\[7\].CLKBUF\[3\] clk vssd1 vssd1 vccd1 vccd1 _13192_/CLK sky130_fd_sc_hd__clkbuf_4
X_11803_ _11825_/CLK line[77] vssd1 vssd1 vccd1 vccd1 _11804_/A sky130_fd_sc_hd__dfxtp_1
X_12783_ _12805_/CLK line[13] vssd1 vssd1 vccd1 vccd1 _12784_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_92_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__04921__A2 _04922_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12000__D line[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11734_ _11734_/A _11759_/Y vssd1 vssd1 vccd1 vccd1 _13694_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11665_ _11685_/CLK line[14] vssd1 vssd1 vccd1 vccd1 _11666_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12935__D line[68] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[24\].VALID\[9\].FF_D A[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13404_ _13898_/Y vssd1 vssd1 vccd1 vccd1 _13404_/Y sky130_fd_sc_hd__inv_2
X_10616_ _10616_/A _10639_/Y vssd1 vssd1 vccd1 vccd1 _13696_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11596_ _11596_/A _11619_/Y vssd1 vssd1 vccd1 vccd1 _13836_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13335_ _13365_/CLK line[0] vssd1 vssd1 vccd1 vccd1 _13336_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_41_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10547_ _10565_/CLK line[15] vssd1 vssd1 vccd1 vccd1 _10548_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[1\].CLKBUF\[3\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13266_ _13266_/A _13299_/Y vssd1 vssd1 vccd1 vccd1 _13826_/Z sky130_fd_sc_hd__ebufn_2
X_10478_ _10478_/A _10499_/Y vssd1 vssd1 vccd1 vccd1 _13838_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08503__A _13913_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12670__D line[80] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12217_ _12245_/CLK line[10] vssd1 vssd1 vccd1 vccd1 _12218_/A sky130_fd_sc_hd__dfxtp_1
X_13197_ _13225_/CLK line[74] vssd1 vssd1 vccd1 vccd1 _13198_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_111_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12148_ _12148_/A _12179_/Y vssd1 vssd1 vccd1 vccd1 _13828_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_150_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11286__D line[82] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11864__A _13927_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDATA\[27\].CLKBUF\[7\] clk vssd1 vssd1 vccd1 vccd1 _10532_/CLK sky130_fd_sc_hd__clkbuf_4
X_04970_ _05000_/CLK line[16] vssd1 vssd1 vccd1 vccd1 _04971_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_2_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12079_ _12105_/CLK line[75] vssd1 vssd1 vccd1 vccd1 _12080_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[12\].VALID\[13\].FF_D A[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11583__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08595__D line[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06640_ _06640_/A _06649_/Y vssd1 vssd1 vccd1 vccd1 _13640_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_25_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06571_ _06575_/CLK line[103] vssd1 vssd1 vccd1 vccd1 _06572_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__04912__A2 _04914_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08310_ _08310_/A _08329_/Y vssd1 vssd1 vccd1 vccd1 _13630_/Z sky130_fd_sc_hd__ebufn_2
X_05522_ _05522_/A _05529_/Y vssd1 vssd1 vccd1 vccd1 _13642_/Z sky130_fd_sc_hd__ebufn_2
X_09290_ _09290_/A _09309_/Y vssd1 vssd1 vccd1 vccd1 _13770_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_33_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07004__D line[59] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XDATA\[6\].CLKBUF\[0\] clk vssd1 vssd1 vccd1 vccd1 _12807_/CLK sky130_fd_sc_hd__clkbuf_4
X_08241_ _08255_/CLK line[98] vssd1 vssd1 vccd1 vccd1 _08242_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12845__D line[32] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05453_ _05455_/CLK line[104] vssd1 vssd1 vccd1 vccd1 _05454_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_193_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[20\].VALID\[2\].FF OVHB\[20\].V/CLK A[9] vssd1 vssd1 vccd1 vccd1 OVHB\[20\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_119_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XOVHB\[2\].VALID\[0\].TOBUF OVHB\[2\].VALID\[0\].FF/Q OVHB\[2\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04924_/B2 sky130_fd_sc_hd__ebufn_2
X_08172_ _08172_/A _08189_/Y vssd1 vssd1 vccd1 vccd1 _13772_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[22\].VALID\[12\].FF_D A[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06843__D line[99] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05384_ _05384_/A _05389_/Y vssd1 vssd1 vccd1 vccd1 _13784_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_174_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07123_ _07135_/CLK line[99] vssd1 vssd1 vccd1 vccd1 _07124_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_118_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[27\].VALID\[3\].TOBUF OVHB\[27\].VALID\[3\].FF/Q OVHB\[27\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04919_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_106_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07054_ _07054_/A _07069_/Y vssd1 vssd1 vccd1 vccd1 _13774_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11758__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[21\].VALID\[14\].TOBUF OVHB\[21\].VALID\[14\].FF/Q OVHB\[21\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__13676__D line[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06005_ _06015_/CLK line[100] vssd1 vssd1 vccd1 vccd1 _06006_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[17\].V_D TIE/HI vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[5\].VALID\[4\].FF_D A[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07956_ _07956_/A _07979_/Y vssd1 vssd1 vccd1 vccd1 _13836_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05194__D line[113] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06907_ _06925_/CLK line[15] vssd1 vssd1 vccd1 vccd1 _06908_/A sky130_fd_sc_hd__dfxtp_1
X_07887_ _07905_/CLK line[79] vssd1 vssd1 vccd1 vccd1 _07888_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11924__D line[118] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09626_ _09626_/A _09659_/Y vssd1 vssd1 vccd1 vccd1 _13826_/Z sky130_fd_sc_hd__ebufn_2
X_06838_ _06838_/A _06859_/Y vssd1 vssd1 vccd1 vccd1 _13838_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_71_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XDATA\[26\].CLKBUF\[4\] clk vssd1 vssd1 vccd1 vccd1 _10147_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_204_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09557_ _09585_/CLK line[74] vssd1 vssd1 vccd1 vccd1 _09558_/A sky130_fd_sc_hd__dfxtp_1
X_06769_ _06785_/CLK line[65] vssd1 vssd1 vccd1 vccd1 _06770_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_102_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08508_ _08508_/A _08539_/Y vssd1 vssd1 vccd1 vccd1 _13828_/Z sky130_fd_sc_hd__ebufn_2
XPHY_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07699__A _13911_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09488_ _09488_/A _09519_/Y vssd1 vssd1 vccd1 vccd1 _13688_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_23_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[19\].VALID\[3\].FF OVHB\[19\].V/CLK A[10] vssd1 vssd1 vccd1 vccd1 OVHB\[19\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08439_ _08465_/CLK line[75] vssd1 vssd1 vccd1 vccd1 _08440_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11450_ _11450_/A _11479_/Y vssd1 vssd1 vccd1 vccd1 _13690_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10401_ _10425_/CLK line[76] vssd1 vssd1 vccd1 vccd1 _10402_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10275__D line[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11381_ _11405_/CLK line[12] vssd1 vssd1 vccd1 vccd1 _11382_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05369__D line[65] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13120_ _13120_/CLK line[25] vssd1 vssd1 vccd1 vccd1 _13121_/A sky130_fd_sc_hd__dfxtp_1
X_10332_ _10332_/A _10359_/Y vssd1 vssd1 vccd1 vccd1 _13692_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13586__D line[124] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[26\].CLKBUF\[6\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12490__D line[121] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13051_ _13051_/A _13054_/Y vssd1 vssd1 vccd1 vccd1 _13891_/Z sky130_fd_sc_hd__ebufn_2
X_10263_ _10285_/CLK line[13] vssd1 vssd1 vccd1 vccd1 _10264_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[19\].VALID\[9\].TOBUF OVHB\[19\].VALID\[9\].FF/Q OVHB\[19\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04914_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_105_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07584__D line[54] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12002_ _12002_/CLK _12003_/X vssd1 vssd1 vccd1 vccd1 _12000_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_78_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10194_ _10194_/A _10219_/Y vssd1 vssd1 vccd1 vccd1 _13834_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_120_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13953_ _13960_/A _13960_/B _13960_/C _13960_/D vssd1 vssd1 vccd1 vccd1 _13953_/Y
+ sky130_fd_sc_hd__nor4b_4
XANTENNA__11834__D line[91] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12904_ _12910_/CLK line[54] vssd1 vssd1 vccd1 vccd1 _12905_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05832__D line[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08993__A _13915_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13884_ _13890_/CLK line[118] vssd1 vssd1 vccd1 vccd1 _13885_/A sky130_fd_sc_hd__dfxtp_1
X_12835_ _12835_/A _12844_/Y vssd1 vssd1 vccd1 vccd1 _13675_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13404__A _13898_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12766_ _12770_/CLK line[119] vssd1 vssd1 vccd1 vccd1 _12767_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XDATA\[25\].CLKBUF\[1\] clk vssd1 vssd1 vccd1 vccd1 _09762_/CLK sky130_fd_sc_hd__clkbuf_4
XPHY_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11717_ _11717_/A _11724_/Y vssd1 vssd1 vccd1 vccd1 _13677_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13123__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12665__D line[73] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12697_ _12697_/A _12704_/Y vssd1 vssd1 vccd1 vccd1 _13817_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_175_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07759__D line[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11648_ _11650_/CLK line[120] vssd1 vssd1 vccd1 vccd1 _11649_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[15\].CLKBUF\[7\] clk vssd1 vssd1 vccd1 vccd1 _06892_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__06018__A _13902_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10185__D line[96] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11579_ _11579_/A _11584_/Y vssd1 vssd1 vccd1 vccd1 _13819_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_116_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13318_ _13330_/CLK line[115] vssd1 vssd1 vccd1 vccd1 _13319_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[17\].VALID\[5\].FF OVHB\[17\].V/CLK A[12] vssd1 vssd1 vccd1 vccd1 OVHB\[17\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_155_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10913__D line[40] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13249_ _13249_/A _13264_/Y vssd1 vssd1 vccd1 vccd1 _13809_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07494__D line[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[5\].VALID\[11\].FF OVHB\[5\].V/CLK A[18] vssd1 vssd1 vccd1 vccd1 OVHB\[5\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_123_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07810_ _07810_/A _07839_/Y vssd1 vssd1 vccd1 vccd1 _13690_/Z sky130_fd_sc_hd__ebufn_2
X_08790_ _08790_/A _08819_/Y vssd1 vssd1 vccd1 vccd1 _13830_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_38_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07741_ _07765_/CLK line[12] vssd1 vssd1 vccd1 vccd1 _07742_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09064__A _13915_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[0\].VALID\[5\].TOBUF OVHB\[0\].VALID\[5\].FF/Q OVHB\[0\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04927_/B2 sky130_fd_sc_hd__ebufn_2
X_04953_ _04965_/CLK line[3] vssd1 vssd1 vccd1 vccd1 _04954_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_65_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07672_ _07672_/A _07699_/Y vssd1 vssd1 vccd1 vccd1 _13832_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[25\].VALID\[8\].TOBUF OVHB\[25\].VALID\[8\].FF/Q OVHB\[25\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04931_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_37_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05742__D line[122] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09411_ _09411_/A _09414_/Y vssd1 vssd1 vccd1 vccd1 _13891_/Z sky130_fd_sc_hd__ebufn_2
X_06623_ _06645_/CLK line[13] vssd1 vssd1 vccd1 vccd1 _06624_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_92_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09342_ _09342_/CLK _09343_/X vssd1 vssd1 vccd1 vccd1 _09340_/CLK sky130_fd_sc_hd__dlclkp_1
X_06554_ _06554_/A _06579_/Y vssd1 vssd1 vccd1 vccd1 _13834_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_61_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05505_ _05525_/CLK line[14] vssd1 vssd1 vccd1 vccd1 _05506_/A sky130_fd_sc_hd__dfxtp_1
X_09273_ _13916_/X wr vssd1 vssd1 vccd1 vccd1 _09273_/X sky130_fd_sc_hd__and2_1
XANTENNA__12575__D line[46] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06485_ _06505_/CLK line[78] vssd1 vssd1 vccd1 vccd1 _06486_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_193_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07669__D line[107] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08224_ _13932_/X vssd1 vssd1 vccd1 vccd1 _08224_/Y sky130_fd_sc_hd__inv_2
XANTENNA__06573__D line[104] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05436_ _05436_/A _05459_/Y vssd1 vssd1 vccd1 vccd1 _13836_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_165_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08155_ _08185_/CLK line[64] vssd1 vssd1 vccd1 vccd1 _08156_/A sky130_fd_sc_hd__dfxtp_1
X_05367_ _05385_/CLK line[79] vssd1 vssd1 vccd1 vccd1 _05368_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10673__A _13924_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09884__D line[81] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07106_ _07106_/A _07139_/Y vssd1 vssd1 vccd1 vccd1 _13826_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09239__A _13916_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08086_ _08086_/A _08119_/Y vssd1 vssd1 vccd1 vccd1 _13686_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_146_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05298_ _05298_/A _05319_/Y vssd1 vssd1 vccd1 vccd1 _13698_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_134_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XDATA\[14\].CLKBUF\[4\] clk vssd1 vssd1 vccd1 vccd1 _06507_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__10823__D line[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07037_ _07065_/CLK line[74] vssd1 vssd1 vccd1 vccd1 _07038_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_134_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[1\].VOBUF OVHB\[1\].V/Q OVHB\[1\].INV/Y vssd1 vssd1 vccd1 vccd1 _04912_/B1
+ sky130_fd_sc_hd__ebufn_2
XANTENNA__05917__D line[74] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08988_ _08990_/CLK line[56] vssd1 vssd1 vccd1 vccd1 _08989_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_57_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XOVHB\[15\].VALID\[7\].FF OVHB\[15\].V/CLK A[14] vssd1 vssd1 vccd1 vccd1 OVHB\[15\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_180_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07939_ _07939_/A _07944_/Y vssd1 vssd1 vccd1 vccd1 _13819_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_56_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10950_ _10950_/CLK line[57] vssd1 vssd1 vccd1 vccd1 _10951_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06748__D line[56] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_OVHB\[19\].VALID\[13\].FF_D A[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09124__D line[118] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09609_ _09609_/A _09624_/Y vssd1 vssd1 vccd1 vccd1 _13809_/Z sky130_fd_sc_hd__ebufn_2
X_10881_ _10881_/A _10884_/Y vssd1 vssd1 vccd1 vccd1 _13681_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10848__A _13925_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12620_ _12630_/CLK line[52] vssd1 vssd1 vccd1 vccd1 _12621_/A sky130_fd_sc_hd__dfxtp_1
XPHY_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12551_ _12551_/A _12564_/Y vssd1 vssd1 vccd1 vccd1 _13671_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11502_ _11510_/CLK line[53] vssd1 vssd1 vccd1 vccd1 _11503_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_169_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06483__D line[77] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12482_ _12490_/CLK line[117] vssd1 vssd1 vccd1 vccd1 _12483_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[31\].VALID\[7\].TOBUF OVHB\[31\].VALID\[7\].FF/Q OVHB\[31\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/A2 sky130_fd_sc_hd__ebufn_2
X_11433_ _11433_/A _11444_/Y vssd1 vssd1 vccd1 vccd1 _13673_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05099__D line[70] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XOVHB\[9\].VALID\[0\].TOBUF OVHB\[9\].VALID\[0\].FF/Q OVHB\[9\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04924_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[29\].VALID\[12\].FF_D A[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11364_ _11370_/CLK line[118] vssd1 vssd1 vccd1 vccd1 _11365_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[19\].VALID\[11\].FF OVHB\[19\].V/CLK A[18] vssd1 vssd1 vccd1 vccd1 OVHB\[19\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_13103_ _13103_/A _13124_/Y vssd1 vssd1 vccd1 vccd1 _13663_/Z sky130_fd_sc_hd__ebufn_2
X_10315_ _10315_/A _10324_/Y vssd1 vssd1 vccd1 vccd1 _13675_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_98_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13894__A _13899_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11295_ _11295_/A _11304_/Y vssd1 vssd1 vccd1 vccd1 _13815_/Z sky130_fd_sc_hd__ebufn_2
X_13034_ _13050_/CLK line[113] vssd1 vssd1 vccd1 vccd1 _13035_/A sky130_fd_sc_hd__dfxtp_1
X_10246_ _10250_/CLK line[119] vssd1 vssd1 vccd1 vccd1 _10247_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[10\].VALID\[0\].FF_D A[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XDATA\[13\].CLKBUF\[1\] clk vssd1 vssd1 vccd1 vccd1 _06122_/CLK sky130_fd_sc_hd__clkbuf_4
X_10177_ _10177_/A _10184_/Y vssd1 vssd1 vccd1 vccd1 _13817_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_94_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11564__D line[81] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06658__D line[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13936_ _13938_/B _13938_/A _13938_/C _13938_/D vssd1 vssd1 vccd1 vccd1 _13936_/X
+ sky130_fd_sc_hd__and4b_4
XANTENNA__09034__D line[91] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13867_ _13867_/A _13894_/Y vssd1 vssd1 vccd1 vccd1 _13867_/Z sky130_fd_sc_hd__ebufn_2
X_12818_ _12840_/CLK line[29] vssd1 vssd1 vccd1 vccd1 _12819_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08873__D line[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[13\].VALID\[9\].FF OVHB\[13\].V/CLK A[16] vssd1 vssd1 vccd1 vccd1 OVHB\[13\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_50_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13798_ _13820_/CLK line[93] vssd1 vssd1 vccd1 vccd1 _13799_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_188_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12749_ _12749_/A _12774_/Y vssd1 vssd1 vccd1 vccd1 _13869_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_175_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06270_ _06270_/A _06299_/Y vssd1 vssd1 vccd1 vccd1 _13830_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13788__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05221_ _05245_/CLK line[12] vssd1 vssd1 vccd1 vccd1 _05222_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_128_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05152_ _05152_/A _05179_/Y vssd1 vssd1 vccd1 vccd1 _13832_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_128_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11739__D line[33] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[1\].VALID\[7\].FF_D A[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09960_ _09970_/CLK line[116] vssd1 vssd1 vccd1 vccd1 _09961_/A sky130_fd_sc_hd__dfxtp_1
X_05083_ _05105_/CLK line[77] vssd1 vssd1 vccd1 vccd1 _05084_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09209__D line[43] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08911_ _08911_/A _08924_/Y vssd1 vssd1 vccd1 vccd1 _13671_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08113__D line[40] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09891_ _09891_/A _09904_/Y vssd1 vssd1 vccd1 vccd1 _13811_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[18\].VALID\[13\].TOBUF OVHB\[18\].VALID\[13\].FF/Q OVHB\[18\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04916_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_111_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08842_ _08850_/CLK line[117] vssd1 vssd1 vccd1 vccd1 _08843_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12213__A _13934_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08773_ _08773_/A _08784_/Y vssd1 vssd1 vccd1 vccd1 _13813_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_85_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05985_ _06015_/CLK line[96] vssd1 vssd1 vccd1 vccd1 _05986_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_38_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07724_ _07730_/CLK line[118] vssd1 vssd1 vccd1 vccd1 _07725_/A sky130_fd_sc_hd__dfxtp_1
X_04936_ _04936_/A _04969_/Y vssd1 vssd1 vccd1 vccd1 _13616_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05472__D line[127] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07655_ _07655_/A _07664_/Y vssd1 vssd1 vccd1 vccd1 _13815_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_26_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06606_ _06610_/CLK line[119] vssd1 vssd1 vccd1 vccd1 _06607_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_53_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07586_ _07590_/CLK line[55] vssd1 vssd1 vccd1 vccd1 _07587_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_43_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09325_ _09325_/A _09344_/Y vssd1 vssd1 vccd1 vccd1 _13805_/Z sky130_fd_sc_hd__ebufn_2
X_06537_ _06537_/A _06544_/Y vssd1 vssd1 vccd1 vccd1 _13817_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[15\].V_RESET_B rst_n vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07399__D line[97] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09256_ _09270_/CLK line[50] vssd1 vssd1 vccd1 vccd1 _09257_/A sky130_fd_sc_hd__dfxtp_1
X_06468_ _06470_/CLK line[56] vssd1 vssd1 vccd1 vccd1 _06469_/A sky130_fd_sc_hd__dfxtp_1
X_08207_ _08207_/A _08224_/Y vssd1 vssd1 vccd1 vccd1 _13807_/Z sky130_fd_sc_hd__ebufn_2
X_05419_ _05419_/A _05424_/Y vssd1 vssd1 vccd1 vccd1 _13819_/Z sky130_fd_sc_hd__ebufn_2
X_09187_ _09187_/A _09204_/Y vssd1 vssd1 vccd1 vccd1 _13667_/Z sky130_fd_sc_hd__ebufn_2
X_06399_ _06399_/A _06404_/Y vssd1 vssd1 vccd1 vccd1 _13679_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[11\].VALID\[12\].TOBUF OVHB\[11\].VALID\[12\].FF/Q OVHB\[11\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04929_/B2 sky130_fd_sc_hd__ebufn_2
X_08138_ _08150_/CLK line[51] vssd1 vssd1 vccd1 vccd1 _08139_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_134_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10553__D line[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08069_ _08069_/A _08084_/Y vssd1 vssd1 vccd1 vccd1 _13669_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_108_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05647__D line[79] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[23\].VALID\[0\].FF_D A[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10100_ _10110_/CLK line[52] vssd1 vssd1 vccd1 vccd1 _10101_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08023__D line[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[8\].CGAND _13898_/Y wr vssd1 vssd1 vccd1 vccd1 OVHB\[8\].CGAND/X sky130_fd_sc_hd__and2_4
X_11080_ _11090_/CLK line[116] vssd1 vssd1 vccd1 vccd1 _11081_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_122_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13864__D line[123] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10031_ _10031_/A _10044_/Y vssd1 vssd1 vccd1 vccd1 _13671_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_0_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07862__D line[53] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_OVHB\[0\].CGAND_A _13931_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[8\].VALID\[0\].FF OVHB\[8\].V/CLK A[7] vssd1 vssd1 vccd1 vccd1 OVHB\[8\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[16\].VALID\[4\].FF_D A[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[19\].CLKBUF\[0\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11982_ _12000_/CLK line[31] vssd1 vssd1 vccd1 vccd1 _11983_/A sky130_fd_sc_hd__dfxtp_1
X_13721_ _13721_/A _13754_/Y vssd1 vssd1 vccd1 vccd1 _13721_/Z sky130_fd_sc_hd__ebufn_2
X_10933_ _10933_/A _10954_/Y vssd1 vssd1 vccd1 vccd1 _13733_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[7\].VALID\[5\].TOBUF OVHB\[7\].VALID\[5\].FF/Q OVHB\[7\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04927_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_205_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09789__D line[38] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10864_ _10880_/CLK line[17] vssd1 vssd1 vccd1 vccd1 _10865_/A sky130_fd_sc_hd__dfxtp_1
X_13652_ _13680_/CLK line[26] vssd1 vssd1 vccd1 vccd1 _13653_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08048__A _13932_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12603_ _12603_/A _12634_/Y vssd1 vssd1 vccd1 vccd1 _13723_/Z sky130_fd_sc_hd__ebufn_2
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10728__D line[83] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10795_ _10795_/A _10814_/Y vssd1 vssd1 vccd1 vccd1 _13875_/Z sky130_fd_sc_hd__ebufn_2
X_13583_ _13583_/A _13614_/Y vssd1 vssd1 vccd1 vccd1 _13863_/Z sky130_fd_sc_hd__ebufn_2
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13104__D line[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12534_ _12560_/CLK line[27] vssd1 vssd1 vccd1 vccd1 _12535_/A sky130_fd_sc_hd__dfxtp_1
XPHY_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12943__D line[72] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12465_ _12465_/A _12494_/Y vssd1 vssd1 vccd1 vccd1 _13865_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_185_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11416_ _11440_/CLK line[28] vssd1 vssd1 vccd1 vccd1 _11417_/A sky130_fd_sc_hd__dfxtp_1
X_12396_ _12420_/CLK line[92] vssd1 vssd1 vccd1 vccd1 _12397_/A sky130_fd_sc_hd__dfxtp_1
X_11347_ _11347_/A _11374_/Y vssd1 vssd1 vccd1 vccd1 _13867_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_113_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11278_ _11300_/CLK line[93] vssd1 vssd1 vccd1 vccd1 _11279_/A sky130_fd_sc_hd__dfxtp_1
X_13017_ _13017_/CLK _13018_/X vssd1 vssd1 vccd1 vccd1 _13015_/CLK sky130_fd_sc_hd__dlclkp_1
X_10229_ _10229_/A _10254_/Y vssd1 vssd1 vccd1 vccd1 _13869_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07772__D line[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11294__D line[86] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06388__D line[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05770_ _05770_/CLK line[121] vssd1 vssd1 vccd1 vccd1 _05771_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_208_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13919_ A[4] vssd1 vssd1 vccd1 vccd1 _13927_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA__09699__D line[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07440_ _07450_/CLK line[116] vssd1 vssd1 vccd1 vccd1 _07441_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_35_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XOVHB\[31\].VALID\[12\].TOBUF OVHB\[31\].VALID\[12\].FF/Q OVHB\[31\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04929_/B2 sky130_fd_sc_hd__ebufn_2
X_07371_ _07371_/A _07384_/Y vssd1 vssd1 vccd1 vccd1 _13811_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[6\].VALID\[2\].FF OVHB\[6\].V/CLK A[9] vssd1 vssd1 vccd1 vccd1 OVHB\[6\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_09110_ _09130_/CLK line[126] vssd1 vssd1 vccd1 vccd1 _09111_/A sky130_fd_sc_hd__dfxtp_1
X_06322_ _06330_/CLK line[117] vssd1 vssd1 vccd1 vccd1 _06323_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_148_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07012__D line[63] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09041_ _09041_/A _09064_/Y vssd1 vssd1 vccd1 vccd1 _13801_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12853__D line[45] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06253_ _06253_/A _06264_/Y vssd1 vssd1 vccd1 vccd1 _13813_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[14\].VALID\[0\].TOBUF OVHB\[14\].VALID\[0\].FF/Q OVHB\[14\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04924_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__07947__D line[106] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05204_ _05210_/CLK line[118] vssd1 vssd1 vccd1 vccd1 _05205_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06851__D line[103] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06184_ _06190_/CLK line[54] vssd1 vssd1 vccd1 vccd1 _06185_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11469__D line[38] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05135_ _05135_/A _05144_/Y vssd1 vssd1 vccd1 vccd1 _13815_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_116_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09943_ _09943_/A _09974_/Y vssd1 vssd1 vccd1 vccd1 _13863_/Z sky130_fd_sc_hd__ebufn_2
X_05066_ _05070_/CLK line[55] vssd1 vssd1 vccd1 vccd1 _05067_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08778__D line[88] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09874_ _09900_/CLK line[91] vssd1 vssd1 vccd1 vccd1 _09875_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_OVHB\[29\].VALID\[4\].FF_D A[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08825_ _08825_/A _08854_/Y vssd1 vssd1 vccd1 vccd1 _13865_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12878__A _13937_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08756_ _08780_/CLK line[92] vssd1 vssd1 vccd1 vccd1 _08757_/A sky130_fd_sc_hd__dfxtp_1
X_05968_ _05980_/CLK line[83] vssd1 vssd1 vccd1 vccd1 _05969_/A sky130_fd_sc_hd__dfxtp_1
X_04919_ A_h[8] _04919_/B2 A_h[8] _04919_/B2 vssd1 vssd1 vccd1 vccd1 _04919_/X sky130_fd_sc_hd__a2bb2o_2
XFILLER_54_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07707_ _07707_/A _07734_/Y vssd1 vssd1 vccd1 vccd1 _13867_/Z sky130_fd_sc_hd__ebufn_2
X_08687_ _08687_/A _08714_/Y vssd1 vssd1 vccd1 vccd1 _13727_/Z sky130_fd_sc_hd__ebufn_2
X_05899_ _05899_/A _05914_/Y vssd1 vssd1 vccd1 vccd1 _13739_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_199_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07638_ _07660_/CLK line[93] vssd1 vssd1 vccd1 vccd1 _07639_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09402__D line[117] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07569_ _07569_/A _07594_/Y vssd1 vssd1 vccd1 vccd1 _13729_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_110_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09308_ _13916_/X wr vssd1 vssd1 vccd1 vccd1 _09308_/X sky130_fd_sc_hd__and2_1
X_10580_ _10600_/CLK line[30] vssd1 vssd1 vccd1 vccd1 _10581_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_194_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09239_ _13916_/X vssd1 vssd1 vccd1 vccd1 _09239_/Y sky130_fd_sc_hd__inv_2
XFILLER_126_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12250_ _12280_/CLK line[16] vssd1 vssd1 vccd1 vccd1 _12251_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06761__D line[76] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11379__D line[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11201_ _11201_/A _11234_/Y vssd1 vssd1 vccd1 vccd1 _13721_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[4\].VALID\[4\].FF OVHB\[4\].V/CLK A[11] vssd1 vssd1 vccd1 vccd1 OVHB\[4\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10283__D line[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12181_ _12181_/A _12214_/Y vssd1 vssd1 vccd1 vccd1 _13861_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.M\[3\].MUX\[0\]_A2 _13819_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05377__D line[69] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11132_ _11160_/CLK line[26] vssd1 vssd1 vccd1 vccd1 _11133_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_107_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13594__D line[113] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11063_ _11063_/A _11094_/Y vssd1 vssd1 vccd1 vccd1 _13863_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_135_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08688__D line[61] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10014_ _10040_/CLK line[27] vssd1 vssd1 vccd1 vccd1 _10015_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_DEC.DEC0.AND3_B A[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06001__D line[98] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11965_ _11965_/CLK line[9] vssd1 vssd1 vccd1 vccd1 _11966_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_205_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11842__D line[95] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13704_ _13704_/A _13719_/Y vssd1 vssd1 vccd1 vccd1 _13704_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06936__D line[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10916_ _10916_/A _10919_/Y vssd1 vssd1 vccd1 vccd1 _13716_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_204_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09312__D line[90] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11896_ _11896_/A _11899_/Y vssd1 vssd1 vccd1 vccd1 _13856_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05840__D line[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13635_ _13645_/CLK line[4] vssd1 vssd1 vccd1 vccd1 _13636_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10458__D line[88] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10847_ _10847_/CLK _10848_/X vssd1 vssd1 vccd1 vccd1 _10845_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA_DATA\[17\].CLKBUF\[2\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13566_ _13566_/A _13579_/Y vssd1 vssd1 vccd1 vccd1 _13846_/Z sky130_fd_sc_hd__ebufn_2
X_10778_ _13924_/X wr vssd1 vssd1 vccd1 vccd1 _10778_/X sky130_fd_sc_hd__and2_1
XFILLER_12_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13769__D line[65] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12517_ _12525_/CLK line[5] vssd1 vssd1 vccd1 vccd1 _12518_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_118_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13497_ _13505_/CLK line[69] vssd1 vssd1 vccd1 vccd1 _13498_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_157_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12448_ _12448_/A _12459_/Y vssd1 vssd1 vccd1 vccd1 _13848_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10193__D line[109] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12379_ _12385_/CLK line[70] vssd1 vssd1 vccd1 vccd1 _12380_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05287__D line[42] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XDATA\[4\].CLKBUF\[5\] clk vssd1 vssd1 vccd1 vccd1 _12422_/CLK sky130_fd_sc_hd__clkbuf_4
X_06940_ _06960_/CLK line[30] vssd1 vssd1 vccd1 vccd1 _06941_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_86_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06871_ _06871_/A _06894_/Y vssd1 vssd1 vccd1 vccd1 _13871_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[2\].VALID\[6\].FF OVHB\[2\].V/CLK A[13] vssd1 vssd1 vccd1 vccd1 OVHB\[2\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_67_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13009__D line[102] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__04925__A2_N _04925_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08610_ _08640_/CLK line[16] vssd1 vssd1 vccd1 vccd1 _08611_/A sky130_fd_sc_hd__dfxtp_1
X_05822_ _05840_/CLK line[31] vssd1 vssd1 vccd1 vccd1 _05823_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_67_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09590_ _09620_/CLK line[80] vssd1 vssd1 vccd1 vccd1 _09591_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_55_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[12\].VALID\[5\].TOBUF OVHB\[12\].VALID\[5\].FF/Q OVHB\[12\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04927_/B2 sky130_fd_sc_hd__ebufn_2
X_08541_ _08541_/A _08574_/Y vssd1 vssd1 vccd1 vccd1 _13861_/Z sky130_fd_sc_hd__ebufn_2
X_05753_ _05753_/A _05774_/Y vssd1 vssd1 vccd1 vccd1 _13873_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_211_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08472_ _08500_/CLK line[90] vssd1 vssd1 vccd1 vccd1 _08473_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_23_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05684_ _05700_/CLK line[81] vssd1 vssd1 vccd1 vccd1 _05685_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05750__D line[126] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07423_ _07423_/A _07454_/Y vssd1 vssd1 vccd1 vccd1 _13863_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_196_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10368__D line[61] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07354_ _07380_/CLK line[91] vssd1 vssd1 vccd1 vccd1 _07355_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_31_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06305_ _06305_/A _06334_/Y vssd1 vssd1 vccd1 vccd1 _13865_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12583__D line[35] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07285_ _07285_/A _07314_/Y vssd1 vssd1 vccd1 vccd1 _13725_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_109_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07677__D line[111] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09024_ _09024_/A _09029_/Y vssd1 vssd1 vccd1 vccd1 _13784_/Z sky130_fd_sc_hd__ebufn_2
X_06236_ _06260_/CLK line[92] vssd1 vssd1 vccd1 vccd1 _06237_/A sky130_fd_sc_hd__dfxtp_1
X_06167_ _06167_/A _06194_/Y vssd1 vssd1 vccd1 vccd1 _13727_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09892__D line[85] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05118_ _05140_/CLK line[93] vssd1 vssd1 vccd1 vccd1 _05119_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_49_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06098_ _06120_/CLK line[29] vssd1 vssd1 vccd1 vccd1 _06099_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10831__D line[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05049_ _05049_/A _05074_/Y vssd1 vssd1 vccd1 vccd1 _13729_/Z sky130_fd_sc_hd__ebufn_2
X_09926_ _09926_/A _09939_/Y vssd1 vssd1 vccd1 vccd1 _13846_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[30\].VALID\[0\].FF OVHB\[30\].V/CLK A[7] vssd1 vssd1 vccd1 vccd1 OVHB\[30\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__05925__D line[78] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[12\].VALID\[7\].FF_D A[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08301__D line[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09857_ _09865_/CLK line[69] vssd1 vssd1 vccd1 vccd1 _09858_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[3\].CLKBUF\[2\] clk vssd1 vssd1 vccd1 vccd1 _12037_/CLK sky130_fd_sc_hd__clkbuf_4
X_08808_ _08808_/A _08819_/Y vssd1 vssd1 vccd1 vccd1 _13848_/Z sky130_fd_sc_hd__ebufn_2
X_09788_ _09788_/A _09799_/Y vssd1 vssd1 vccd1 vccd1 _13708_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_45_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08739_ _08745_/CLK line[70] vssd1 vssd1 vccd1 vccd1 _08740_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12758__D line[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ _11750_/A _11759_/Y vssd1 vssd1 vccd1 vccd1 _13710_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[0\].VALID\[8\].FF OVHB\[0\].V/CLK A[15] vssd1 vssd1 vccd1 vccd1 OVHB\[0\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10701_ _10705_/CLK line[71] vssd1 vssd1 vccd1 vccd1 _10702_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11681_ _11685_/CLK line[7] vssd1 vssd1 vccd1 vccd1 _11682_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13420_ _13420_/A _13439_/Y vssd1 vssd1 vccd1 vccd1 _13700_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10632_ _10632_/A _10639_/Y vssd1 vssd1 vccd1 vccd1 _13712_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13351_ _13365_/CLK line[2] vssd1 vssd1 vccd1 vccd1 _13352_/A sky130_fd_sc_hd__dfxtp_1
X_10563_ _10565_/CLK line[8] vssd1 vssd1 vccd1 vccd1 _10564_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_139_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12302_ _12302_/A _12319_/Y vssd1 vssd1 vccd1 vccd1 _13702_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06491__D line[66] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10494_ _10494_/A _10499_/Y vssd1 vssd1 vccd1 vccd1 _13854_/Z sky130_fd_sc_hd__ebufn_2
X_13282_ _13282_/A _13299_/Y vssd1 vssd1 vccd1 vccd1 _13842_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_6_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12233_ _12245_/CLK line[3] vssd1 vssd1 vccd1 vccd1 _12234_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_123_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12164_ _12164_/A _12179_/Y vssd1 vssd1 vccd1 vccd1 _13844_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_122_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XDATA\[23\].CLKBUF\[6\] clk vssd1 vssd1 vccd1 vccd1 _09377_/CLK sky130_fd_sc_hd__clkbuf_4
XOVHB\[29\].VALID\[1\].FF OVHB\[29\].V/CLK A[8] vssd1 vssd1 vccd1 vccd1 OVHB\[29\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_11115_ _11125_/CLK line[4] vssd1 vssd1 vccd1 vccd1 _11116_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_111_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12095_ _12105_/CLK line[68] vssd1 vssd1 vccd1 vccd1 _12096_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_122_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MUX.M\[2\].MUX\[1\]_A0 _13665_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11046_ _11046_/A _11059_/Y vssd1 vssd1 vccd1 vccd1 _13846_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_39_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__04924__B1 A_h[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11572__D line[85] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12997_ _13015_/CLK line[111] vssd1 vssd1 vccd1 vccd1 _12998_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06666__D line[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11948_ _11948_/A _11969_/Y vssd1 vssd1 vccd1 vccd1 _13628_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_45_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09042__D line[95] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11879_ _11895_/CLK line[97] vssd1 vssd1 vccd1 vccd1 _11880_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09977__D line[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06963__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13618_ _13618_/A _13649_/Y vssd1 vssd1 vccd1 vccd1 _13618_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08881__D line[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13499__D line[70] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[28\].VALID\[11\].TOBUF OVHB\[28\].VALID\[11\].FF/Q OVHB\[28\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04915_/B2 sky130_fd_sc_hd__ebufn_2
X_13549_ _13575_/CLK line[107] vssd1 vssd1 vccd1 vccd1 _13550_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_173_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XOVHB\[1\].VALID\[14\].TOBUF OVHB\[1\].VALID\[14\].FF/Q OVHB\[1\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07070_ _07100_/CLK line[80] vssd1 vssd1 vccd1 vccd1 _07071_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_146_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06021_ _06021_/A _06054_/Y vssd1 vssd1 vccd1 vccd1 _13861_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[15\].CLKBUF\[4\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[25\].VALID\[7\].FF_D A[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11747__D line[37] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07972_ _07972_/A _07979_/Y vssd1 vssd1 vccd1 vccd1 _13852_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09217__D line[47] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09711_ _09725_/CLK line[2] vssd1 vssd1 vccd1 vccd1 _09712_/A sky130_fd_sc_hd__dfxtp_1
X_06923_ _06925_/CLK line[8] vssd1 vssd1 vccd1 vccd1 _06924_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_95_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XDATA\[22\].CLKBUF\[3\] clk vssd1 vssd1 vccd1 vccd1 _08992_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_68_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09642_ _09642_/A _09659_/Y vssd1 vssd1 vccd1 vccd1 _13842_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_67_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06854_ _06854_/A _06859_/Y vssd1 vssd1 vccd1 vccd1 _13854_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_27_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XOVHB\[27\].VALID\[3\].FF OVHB\[27\].V/CLK A[10] vssd1 vssd1 vccd1 vccd1 OVHB\[27\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_05805_ _05805_/CLK line[9] vssd1 vssd1 vccd1 vccd1 _05806_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__04915__B1 A_h[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06785_ _06785_/CLK line[73] vssd1 vssd1 vccd1 vccd1 _06786_/A sky130_fd_sc_hd__dfxtp_1
X_09573_ _09585_/CLK line[67] vssd1 vssd1 vccd1 vccd1 _09574_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_209_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11482__D line[58] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XOVHB\[21\].VALID\[10\].TOBUF OVHB\[21\].VALID\[10\].FF/Q OVHB\[21\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04932_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_36_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08524_ _08524_/A _08539_/Y vssd1 vssd1 vccd1 vccd1 _13844_/Z sky130_fd_sc_hd__ebufn_2
X_05736_ _05736_/A _05739_/Y vssd1 vssd1 vccd1 vccd1 _13856_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[8\].CLKBUF\[4\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05480__D line[116] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10098__D line[51] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05667_ _05667_/CLK _05668_/X vssd1 vssd1 vccd1 vccd1 _05665_/CLK sky130_fd_sc_hd__dlclkp_1
X_08455_ _08465_/CLK line[68] vssd1 vssd1 vccd1 vccd1 _08456_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07406_ _07406_/A _07419_/Y vssd1 vssd1 vccd1 vccd1 _13846_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08791__D line[108] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08386_ _08386_/A _08399_/Y vssd1 vssd1 vccd1 vccd1 _13706_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05598_ _13901_/X wr vssd1 vssd1 vccd1 vccd1 _05598_/X sky130_fd_sc_hd__and2_1
XPHY_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07337_ _07345_/CLK line[69] vssd1 vssd1 vccd1 vccd1 _07338_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_183_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07268_ _07268_/A _07279_/Y vssd1 vssd1 vccd1 vccd1 _13708_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_191_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06219_ _06225_/CLK line[70] vssd1 vssd1 vccd1 vccd1 _06220_/A sky130_fd_sc_hd__dfxtp_1
X_09007_ _09025_/CLK line[79] vssd1 vssd1 vccd1 vccd1 _09008_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_152_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07199_ _07205_/CLK line[6] vssd1 vssd1 vccd1 vccd1 _07200_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_151_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11657__D line[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[6\].VALID\[12\].FF_D A[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10561__D line[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05655__D line[68] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08031__D line[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09909_ _09935_/CLK line[107] vssd1 vssd1 vccd1 vccd1 _09910_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_59_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13872__D line[127] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12920_ _12920_/A _12949_/Y vssd1 vssd1 vccd1 vccd1 _13760_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08966__D line[60] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07870__D line[57] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12851_ _12875_/CLK line[44] vssd1 vssd1 vccd1 vccd1 _12852_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12488__D line[120] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11802_ _11802_/A _11829_/Y vssd1 vssd1 vccd1 vccd1 _13762_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_199_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XDATA\[21\].CLKBUF\[0\] clk vssd1 vssd1 vccd1 vccd1 _08607_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_27_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[6\].VALID\[2\].FF_D A[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12782_ _12782_/A _12809_/Y vssd1 vssd1 vccd1 vccd1 _13622_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05390__D line[80] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[19\].VALID\[5\].TOBUF OVHB\[19\].VALID\[5\].FF/Q OVHB\[19\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04927_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_92_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11733_ _11755_/CLK line[45] vssd1 vssd1 vccd1 vccd1 _11734_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XDATA\[11\].CLKBUF\[6\] clk vssd1 vssd1 vccd1 vccd1 _05737_/CLK sky130_fd_sc_hd__clkbuf_4
XPHY_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[25\].VALID\[5\].FF OVHB\[25\].V/CLK A[12] vssd1 vssd1 vccd1 vccd1 OVHB\[25\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_11664_ _11664_/A _11689_/Y vssd1 vssd1 vccd1 vccd1 _13624_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13403_ _13898_/Y wr vssd1 vssd1 vccd1 vccd1 _13403_/X sky130_fd_sc_hd__and2_1
XPHY_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10736__D line[87] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10615_ _10635_/CLK line[46] vssd1 vssd1 vccd1 vccd1 _10616_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13897__A A[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13112__D line[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11595_ _11615_/CLK line[110] vssd1 vssd1 vccd1 vccd1 _11596_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08206__D line[82] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13334_ _13938_/X vssd1 vssd1 vccd1 vccd1 _13334_/Y sky130_fd_sc_hd__inv_2
X_10546_ _10546_/A _10569_/Y vssd1 vssd1 vccd1 vccd1 _13626_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_41_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13265_ _13295_/CLK line[96] vssd1 vssd1 vccd1 vccd1 _13266_/A sky130_fd_sc_hd__dfxtp_1
X_10477_ _10495_/CLK line[111] vssd1 vssd1 vccd1 vccd1 _10478_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_6_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08503__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12216_ _12216_/A _12249_/Y vssd1 vssd1 vccd1 vccd1 _13616_/Z sky130_fd_sc_hd__ebufn_2
X_13196_ _13196_/A _13229_/Y vssd1 vssd1 vccd1 vccd1 _13756_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10471__D line[108] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12147_ _12175_/CLK line[106] vssd1 vssd1 vccd1 vccd1 _12148_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05565__D line[32] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12078_ _12078_/A _12109_/Y vssd1 vssd1 vccd1 vccd1 _13758_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_2_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11029_ _11055_/CLK line[107] vssd1 vssd1 vccd1 vccd1 _11030_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07780__D line[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12398__D line[93] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06396__D line[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06570_ _06570_/A _06579_/Y vssd1 vssd1 vccd1 vccd1 _13850_/Z sky130_fd_sc_hd__ebufn_2
X_05521_ _05525_/CLK line[7] vssd1 vssd1 vccd1 vccd1 _05522_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_178_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08240_ _08240_/A _08259_/Y vssd1 vssd1 vccd1 vccd1 _13840_/Z sky130_fd_sc_hd__ebufn_2
X_05452_ _05452_/A _05459_/Y vssd1 vssd1 vccd1 vccd1 _13852_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_193_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08171_ _08185_/CLK line[66] vssd1 vssd1 vccd1 vccd1 _08172_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10646__D line[60] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05383_ _05385_/CLK line[72] vssd1 vssd1 vccd1 vccd1 _05384_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[0\].VALID\[1\].TOBUF OVHB\[0\].VALID\[1\].FF/Q OVHB\[0\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04926_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__13022__D line[122] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07122_ _07122_/A _07139_/Y vssd1 vssd1 vccd1 vccd1 _13842_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_186_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XDATA\[10\].CLKBUF\[3\] clk vssd1 vssd1 vccd1 vccd1 _05352_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__07020__D line[52] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[25\].VALID\[4\].TOBUF OVHB\[25\].VALID\[4\].FF/Q OVHB\[25\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04925_/B2 sky130_fd_sc_hd__ebufn_2
X_07053_ _07065_/CLK line[67] vssd1 vssd1 vccd1 vccd1 _07054_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12861__D line[34] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07955__D line[110] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06004_ _06004_/A _06019_/Y vssd1 vssd1 vccd1 vccd1 _13844_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[23\].VALID\[7\].FF OVHB\[23\].V/CLK A[14] vssd1 vssd1 vccd1 vccd1 OVHB\[23\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_142_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07955_ _07975_/CLK line[110] vssd1 vssd1 vccd1 vccd1 _07956_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[13\].CLKBUF\[6\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06906_ _06906_/A _06929_/Y vssd1 vssd1 vccd1 vccd1 _13626_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07886_ _07886_/A _07909_/Y vssd1 vssd1 vccd1 vccd1 _13766_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_56_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09625_ _09655_/CLK line[96] vssd1 vssd1 vccd1 vccd1 _09626_/A sky130_fd_sc_hd__dfxtp_1
X_06837_ _06855_/CLK line[111] vssd1 vssd1 vccd1 vccd1 _06838_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12101__D line[71] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09556_ _09556_/A _09589_/Y vssd1 vssd1 vccd1 vccd1 _13756_/Z sky130_fd_sc_hd__ebufn_2
X_06768_ _06768_/A _06789_/Y vssd1 vssd1 vccd1 vccd1 _13768_/Z sky130_fd_sc_hd__ebufn_2
XPHY_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08507_ _08535_/CLK line[106] vssd1 vssd1 vccd1 vccd1 _08508_/A sky130_fd_sc_hd__dfxtp_1
XPHY_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05719_ _05735_/CLK line[97] vssd1 vssd1 vccd1 vccd1 _05720_/A sky130_fd_sc_hd__dfxtp_1
XPHY_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06699_ _06715_/CLK line[33] vssd1 vssd1 vccd1 vccd1 _06700_/A sky130_fd_sc_hd__dfxtp_1
X_09487_ _09515_/CLK line[42] vssd1 vssd1 vccd1 vccd1 _09488_/A sky130_fd_sc_hd__dfxtp_1
XPHY_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08438_ _08438_/A _08469_/Y vssd1 vssd1 vccd1 vccd1 _13758_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09410__D line[121] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XDECH.DEC0.AND0 A_h[3] A_h[4] vssd1 vssd1 vccd1 vccd1 _13982_/D sky130_fd_sc_hd__nor2_2
XPHY_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08369_ _08395_/CLK line[43] vssd1 vssd1 vccd1 vccd1 _08370_/A sky130_fd_sc_hd__dfxtp_1
X_10400_ _10400_/A _10429_/Y vssd1 vssd1 vccd1 vccd1 _13760_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[6\].CLKBUF\[6\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11380_ _11380_/A _11409_/Y vssd1 vssd1 vccd1 vccd1 _13620_/Z sky130_fd_sc_hd__ebufn_2
X_10331_ _10355_/CLK line[44] vssd1 vssd1 vccd1 vccd1 _10332_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_164_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10262_ _10262_/A _10289_/Y vssd1 vssd1 vccd1 vccd1 _13622_/Z sky130_fd_sc_hd__ebufn_2
X_13050_ _13050_/CLK line[121] vssd1 vssd1 vccd1 vccd1 _13051_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06124__A _13903_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11387__D line[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12001_ _12001_/A _12004_/Y vssd1 vssd1 vccd1 vccd1 _13681_/Z sky130_fd_sc_hd__ebufn_2
X_10193_ _10215_/CLK line[109] vssd1 vssd1 vccd1 vccd1 _10194_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05385__D line[73] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08696__D line[50] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[21\].VALID\[9\].FF OVHB\[21\].V/CLK A[16] vssd1 vssd1 vccd1 vccd1 OVHB\[21\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_13952_ A_h[2] vssd1 vssd1 vccd1 vccd1 _13960_/C sky130_fd_sc_hd__clkbuf_2
XOVHB\[31\].VALID\[3\].TOBUF OVHB\[31\].VALID\[3\].FF/Q OVHB\[31\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04919_/B2 sky130_fd_sc_hd__ebufn_2
X_12903_ _12903_/A _12914_/Y vssd1 vssd1 vccd1 vccd1 _13743_/Z sky130_fd_sc_hd__ebufn_2
X_13883_ _13883_/A _13894_/Y vssd1 vssd1 vccd1 vccd1 _13883_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_34_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08993__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12011__D line[44] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12834_ _12840_/CLK line[22] vssd1 vssd1 vccd1 vccd1 _12835_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_74_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07105__D line[96] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12765_ _12765_/A _12774_/Y vssd1 vssd1 vccd1 vccd1 _13885_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11850__D line[84] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06944__D line[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11716_ _11720_/CLK line[23] vssd1 vssd1 vccd1 vccd1 _11717_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09320__D line[94] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12696_ _12700_/CLK line[87] vssd1 vssd1 vccd1 vccd1 _12697_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11647_ _11647_/A _11654_/Y vssd1 vssd1 vccd1 vccd1 _13887_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06018__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11578_ _11580_/CLK line[88] vssd1 vssd1 vccd1 vccd1 _11579_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13777__D line[69] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13317_ _13317_/A _13334_/Y vssd1 vssd1 vccd1 vccd1 _13877_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_183_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10529_ _10529_/A _10534_/Y vssd1 vssd1 vccd1 vccd1 _13889_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_115_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13248_ _13260_/CLK line[83] vssd1 vssd1 vccd1 vccd1 _13249_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09043__TE_B _09064_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13179_ _13179_/A _13194_/Y vssd1 vssd1 vccd1 vccd1 _13739_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05295__D line[46] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_04952_ _04952_/A _04969_/Y vssd1 vssd1 vccd1 vccd1 _13632_/Z sky130_fd_sc_hd__ebufn_2
X_07740_ _07740_/A _07769_/Y vssd1 vssd1 vccd1 vccd1 _13620_/Z sky130_fd_sc_hd__ebufn_2
X_07671_ _07695_/CLK line[108] vssd1 vssd1 vccd1 vccd1 _07672_/A sky130_fd_sc_hd__dfxtp_1
X_09410_ _09410_/CLK line[121] vssd1 vssd1 vccd1 vccd1 _09411_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_25_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06622_ _06622_/A _06649_/Y vssd1 vssd1 vccd1 vccd1 _13622_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[23\].VALID\[9\].TOBUF OVHB\[23\].VALID\[9\].FF/Q OVHB\[23\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04914_/B2 sky130_fd_sc_hd__ebufn_2
X_09341_ _09341_/A _09344_/Y vssd1 vssd1 vccd1 vccd1 _13821_/Z sky130_fd_sc_hd__ebufn_2
X_06553_ _06575_/CLK line[109] vssd1 vssd1 vccd1 vccd1 _06554_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11760__D line[48] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05504_ _05504_/A _05529_/Y vssd1 vssd1 vccd1 vccd1 _13624_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[14\].V_RESET_B rst_n vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06484_ _06484_/A _06509_/Y vssd1 vssd1 vccd1 vccd1 _13764_/Z sky130_fd_sc_hd__ebufn_2
X_09272_ _09272_/CLK _09273_/X vssd1 vssd1 vccd1 vccd1 _09270_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_20_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10376__D line[50] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05435_ _05455_/CLK line[110] vssd1 vssd1 vccd1 vccd1 _05436_/A sky130_fd_sc_hd__dfxtp_1
X_08223_ _13932_/X wr vssd1 vssd1 vccd1 vccd1 _08223_/X sky130_fd_sc_hd__and2_1
XFILLER_166_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10954__A _13925_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05366_ _05366_/A _05389_/Y vssd1 vssd1 vccd1 vccd1 _13766_/Z sky130_fd_sc_hd__ebufn_2
X_08154_ _13932_/X vssd1 vssd1 vccd1 vccd1 _08154_/Y sky130_fd_sc_hd__inv_2
XANTENNA__10673__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13687__D line[42] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07105_ _07135_/CLK line[96] vssd1 vssd1 vccd1 vccd1 _07106_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12591__D line[39] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08085_ _08115_/CLK line[32] vssd1 vssd1 vccd1 vccd1 _08086_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_146_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05297_ _05315_/CLK line[47] vssd1 vssd1 vccd1 vccd1 _05298_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07685__D line[100] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07036_ _07036_/A _07069_/Y vssd1 vssd1 vccd1 vccd1 _13756_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_164_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_DATA\[27\].CLKBUF\[0\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11000__D line[94] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08987_ _08987_/A _08994_/Y vssd1 vssd1 vccd1 vccd1 _13747_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11935__D line[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07938_ _07940_/CLK line[88] vssd1 vssd1 vccd1 vccd1 _07939_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05933__D line[67] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_OVHB\[2\].VALID\[5\].FF_D A[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07869_ _07869_/A _07874_/Y vssd1 vssd1 vccd1 vccd1 _13749_/Z sky130_fd_sc_hd__ebufn_2
X_09608_ _09620_/CLK line[83] vssd1 vssd1 vccd1 vccd1 _09609_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_113_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10880_ _10880_/CLK line[25] vssd1 vssd1 vccd1 vccd1 _10881_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_43_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10848__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09539_ _09539_/A _09554_/Y vssd1 vssd1 vccd1 vccd1 _13739_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12766__D line[119] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XOVHB\[4\].CGAND _13935_/X wr vssd1 vssd1 vccd1 vccd1 OVHB\[4\].CGAND/X sky130_fd_sc_hd__and2_4
XPHY_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12550_ _12560_/CLK line[20] vssd1 vssd1 vccd1 vccd1 _12551_/A sky130_fd_sc_hd__dfxtp_1
XPHY_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11501_ _11501_/A _11514_/Y vssd1 vssd1 vccd1 vccd1 _13741_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12481_ _12481_/A _12494_/Y vssd1 vssd1 vccd1 vccd1 _13881_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11432_ _11440_/CLK line[21] vssd1 vssd1 vccd1 vccd1 _11433_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_MUX.M\[3\].MUX\[3\]_A0 _13655_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11363_ _11363_/A _11374_/Y vssd1 vssd1 vccd1 vccd1 _13883_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[7\].VALID\[1\].TOBUF OVHB\[7\].VALID\[1\].FF/Q OVHB\[7\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04926_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__07595__D line[64] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13102_ _13120_/CLK line[31] vssd1 vssd1 vccd1 vccd1 _13103_/A sky130_fd_sc_hd__dfxtp_1
X_10314_ _10320_/CLK line[22] vssd1 vssd1 vccd1 vccd1 _10315_/A sky130_fd_sc_hd__dfxtp_1
X_11294_ _11300_/CLK line[86] vssd1 vssd1 vccd1 vccd1 _11295_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_152_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13033_ _13033_/A _13054_/Y vssd1 vssd1 vccd1 vccd1 _13873_/Z sky130_fd_sc_hd__ebufn_2
X_10245_ _10245_/A _10254_/Y vssd1 vssd1 vccd1 vccd1 _13885_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06789__A _13905_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10176_ _10180_/CLK line[87] vssd1 vssd1 vccd1 vccd1 _10177_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_94_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13935_ _13938_/A _13938_/B _13938_/C _13938_/D vssd1 vssd1 vccd1 vccd1 _13935_/X
+ sky130_fd_sc_hd__and4bb_4
XFILLER_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_OVHB\[13\].VALID\[14\].FF_D A[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13866_ _13890_/CLK line[124] vssd1 vssd1 vccd1 vccd1 _13867_/A sky130_fd_sc_hd__dfxtp_1
X_12817_ _12817_/A _12844_/Y vssd1 vssd1 vccd1 vccd1 _13657_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12676__D line[92] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11580__D line[89] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13797_ _13797_/A _13824_/Y vssd1 vssd1 vccd1 vccd1 _13797_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06674__D line[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[16\].V_D TIE/HI vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12748_ _12770_/CLK line[125] vssd1 vssd1 vccd1 vccd1 _12749_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09050__D line[84] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[17\].VALID\[2\].FF_D A[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12679_ _12679_/A _12704_/Y vssd1 vssd1 vccd1 vccd1 _13799_/Z sky130_fd_sc_hd__ebufn_2
XPHY_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09985__D line[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05220_ _05220_/A _05249_/Y vssd1 vssd1 vccd1 vccd1 _13620_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_156_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[23\].VALID\[13\].FF_D A[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[14\].VALID\[14\].TOBUF OVHB\[14\].VALID\[14\].FF/Q OVHB\[14\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/B2 sky130_fd_sc_hd__ebufn_2
X_05151_ _05175_/CLK line[108] vssd1 vssd1 vccd1 vccd1 _05152_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10924__D line[59] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13300__D line[112] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05082_ _05082_/A _05109_/Y vssd1 vssd1 vccd1 vccd1 _13762_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_143_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08910_ _08920_/CLK line[20] vssd1 vssd1 vccd1 vccd1 _08911_/A sky130_fd_sc_hd__dfxtp_1
X_09890_ _09900_/CLK line[84] vssd1 vssd1 vccd1 vccd1 _09891_/A sky130_fd_sc_hd__dfxtp_1
X_08841_ _08841_/A _08854_/Y vssd1 vssd1 vccd1 vccd1 _13881_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12213__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11755__D line[41] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08772_ _08780_/CLK line[85] vssd1 vssd1 vccd1 vccd1 _08773_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06849__D line[102] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05984_ _13902_/X vssd1 vssd1 vccd1 vccd1 _05984_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09225__D line[36] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05108__A _13931_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07723_ _07723_/A _07734_/Y vssd1 vssd1 vccd1 vccd1 _13883_/Z sky130_fd_sc_hd__ebufn_2
X_04935_ _04965_/CLK line[0] vssd1 vssd1 vccd1 vccd1 _04936_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_53_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07654_ _07660_/CLK line[86] vssd1 vssd1 vccd1 vccd1 _07655_/A sky130_fd_sc_hd__dfxtp_1
X_06605_ _06605_/A _06614_/Y vssd1 vssd1 vccd1 vccd1 _13885_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[8\].VALID\[9\].FF_D A[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11490__D line[62] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07585_ _07585_/A _07594_/Y vssd1 vssd1 vccd1 vccd1 _13745_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_179_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09324_ _09340_/CLK line[81] vssd1 vssd1 vccd1 vccd1 _09325_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_43_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06584__D line[123] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06536_ _06540_/CLK line[87] vssd1 vssd1 vccd1 vccd1 _06537_/A sky130_fd_sc_hd__dfxtp_1
X_09255_ _09255_/A _09274_/Y vssd1 vssd1 vccd1 vccd1 _13735_/Z sky130_fd_sc_hd__ebufn_2
X_06467_ _06467_/A _06474_/Y vssd1 vssd1 vccd1 vccd1 _13747_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[1\].CLKBUF\[7\] clk vssd1 vssd1 vccd1 vccd1 _08292_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_21_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08206_ _08220_/CLK line[82] vssd1 vssd1 vccd1 vccd1 _08207_/A sky130_fd_sc_hd__dfxtp_1
X_05418_ _05420_/CLK line[88] vssd1 vssd1 vccd1 vccd1 _05419_/A sky130_fd_sc_hd__dfxtp_1
X_09186_ _09200_/CLK line[18] vssd1 vssd1 vccd1 vccd1 _09187_/A sky130_fd_sc_hd__dfxtp_1
X_06398_ _06400_/CLK line[24] vssd1 vssd1 vccd1 vccd1 _06399_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_5_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08154__A _13932_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05349_ _05349_/A _05354_/Y vssd1 vssd1 vccd1 vccd1 _13749_/Z sky130_fd_sc_hd__ebufn_2
X_08137_ _08137_/A _08154_/Y vssd1 vssd1 vccd1 vccd1 _13737_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_107_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[15\].VALID\[10\].FF_D A[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08068_ _08080_/CLK line[19] vssd1 vssd1 vccd1 vccd1 _08069_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_108_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07019_ _07019_/A _07034_/Y vssd1 vssd1 vccd1 vccd1 _13739_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_108_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_MUX.SEL0BUF\[2\]_A A[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10030_ _10040_/CLK line[20] vssd1 vssd1 vccd1 vccd1 _10031_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11665__D line[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_OVHB\[16\].CG_CLK clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[0\].CGAND_B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06759__D line[75] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09135__D line[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05663__D line[72] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XDATA\[31\].CLKBUF\[5\] clk vssd1 vssd1 vccd1 vccd1 _11862_/CLK sky130_fd_sc_hd__clkbuf_4
X_11981_ _11981_/A _12004_/Y vssd1 vssd1 vccd1 vccd1 _13661_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_29_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13880__D line[116] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[25\].CLKBUF\[2\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[4\].CGAND_A _13935_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13720_ _13750_/CLK line[48] vssd1 vssd1 vccd1 vccd1 _13721_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08974__D line[49] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10932_ _10950_/CLK line[63] vssd1 vssd1 vccd1 vccd1 _10933_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08329__A _13913_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[5\].VALID\[6\].TOBUF OVHB\[5\].VALID\[6\].FF/Q OVHB\[5\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04923_/A2 sky130_fd_sc_hd__ebufn_2
XFILLER_16_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13651_ _13651_/A _13684_/Y vssd1 vssd1 vccd1 vccd1 _13651_/Z sky130_fd_sc_hd__ebufn_2
X_10863_ _10863_/A _10884_/Y vssd1 vssd1 vccd1 vccd1 _13663_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08048__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12602_ _12630_/CLK line[58] vssd1 vssd1 vccd1 vccd1 _12603_/A sky130_fd_sc_hd__dfxtp_1
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13582_ _13610_/CLK line[122] vssd1 vssd1 vccd1 vccd1 _13583_/A sky130_fd_sc_hd__dfxtp_1
X_10794_ _10810_/CLK line[113] vssd1 vssd1 vccd1 vccd1 _10795_/A sky130_fd_sc_hd__dfxtp_1
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12533_ _12533_/A _12564_/Y vssd1 vssd1 vccd1 vccd1 _13653_/Z sky130_fd_sc_hd__ebufn_2
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12464_ _12490_/CLK line[123] vssd1 vssd1 vccd1 vccd1 _12465_/A sky130_fd_sc_hd__dfxtp_1
X_11415_ _11415_/A _11444_/Y vssd1 vssd1 vccd1 vccd1 _13655_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_126_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13120__D line[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12395_ _12395_/A _12424_/Y vssd1 vssd1 vccd1 vccd1 _13795_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05838__D line[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDATA\[0\].CLKBUF\[4\] clk vssd1 vssd1 vccd1 vccd1 _05107_/CLK sky130_fd_sc_hd__clkbuf_4
X_11346_ _11370_/CLK line[124] vssd1 vssd1 vccd1 vccd1 _11347_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08214__D line[86] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11277_ _11277_/A _11304_/Y vssd1 vssd1 vccd1 vccd1 _13797_/Z sky130_fd_sc_hd__ebufn_2
X_13016_ _13016_/A _13019_/Y vssd1 vssd1 vccd1 vccd1 _13856_/Z sky130_fd_sc_hd__ebufn_2
X_10228_ _10250_/CLK line[125] vssd1 vssd1 vccd1 vccd1 _10229_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_140_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10159_ _10159_/A _10184_/Y vssd1 vssd1 vccd1 vccd1 _13799_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05573__D line[45] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09623__A _13920_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13790__D line[80] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13918_ A[3] vssd1 vssd1 vccd1 vccd1 _13927_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_50_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13849_ _13855_/CLK line[102] vssd1 vssd1 vccd1 vccd1 _13850_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12984__A _13937_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDATA\[30\].CLKBUF\[2\] clk vssd1 vssd1 vccd1 vccd1 _11477_/CLK sky130_fd_sc_hd__clkbuf_4
X_07370_ _07380_/CLK line[84] vssd1 vssd1 vccd1 vccd1 _07371_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_50_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06321_ _06321_/A _06334_/Y vssd1 vssd1 vccd1 vccd1 _13881_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05598__A _13901_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09040_ _09060_/CLK line[94] vssd1 vssd1 vccd1 vccd1 _09041_/A sky130_fd_sc_hd__dfxtp_1
X_06252_ _06260_/CLK line[85] vssd1 vssd1 vccd1 vccd1 _06253_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_176_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05203_ _05203_/A _05214_/Y vssd1 vssd1 vccd1 vccd1 _13883_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10654__D line[49] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06183_ _06183_/A _06194_/Y vssd1 vssd1 vccd1 vccd1 _13743_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[12\].VALID\[1\].TOBUF OVHB\[12\].VALID\[1\].FF/Q OVHB\[12\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04926_/B2 sky130_fd_sc_hd__ebufn_2
XOVHB\[9\].VALID\[7\].FF OVHB\[9\].V/CLK A[14] vssd1 vssd1 vccd1 vccd1 OVHB\[9\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10009__A _13922_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13030__D line[126] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05748__D line[125] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05134_ _05140_/CLK line[86] vssd1 vssd1 vccd1 vccd1 _05135_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08124__D line[59] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMUX.SEL1BUF\[1\] A[1] vssd1 vssd1 vccd1 vccd1 MUX.SEL1BUF\[1\]/X sky130_fd_sc_hd__clkbuf_2
X_09942_ _09970_/CLK line[122] vssd1 vssd1 vccd1 vccd1 _09943_/A sky130_fd_sc_hd__dfxtp_1
X_05065_ _05065_/A _05074_/Y vssd1 vssd1 vccd1 vccd1 _13745_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_131_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07963__D line[99] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09873_ _09873_/A _09904_/Y vssd1 vssd1 vccd1 vccd1 _13793_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_100_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08824_ _08850_/CLK line[123] vssd1 vssd1 vccd1 vccd1 _08825_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12878__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08755_ _08755_/A _08784_/Y vssd1 vssd1 vccd1 vccd1 _13795_/Z sky130_fd_sc_hd__ebufn_2
X_05967_ _05967_/A _05984_/Y vssd1 vssd1 vccd1 vccd1 _13807_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_72_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07706_ _07730_/CLK line[124] vssd1 vssd1 vccd1 vccd1 _07707_/A sky130_fd_sc_hd__dfxtp_1
X_04918_ A_h[11] vssd1 vssd1 vccd1 vccd1 _04918_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08686_ _08710_/CLK line[60] vssd1 vssd1 vccd1 vccd1 _08687_/A sky130_fd_sc_hd__dfxtp_1
X_05898_ _05910_/CLK line[51] vssd1 vssd1 vccd1 vccd1 _05899_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10829__D line[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07637_ _07637_/A _07664_/Y vssd1 vssd1 vccd1 vccd1 _13797_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13205__D line[78] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07568_ _07590_/CLK line[61] vssd1 vssd1 vccd1 vccd1 _07569_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07203__D line[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09307_ _09307_/CLK _09308_/X vssd1 vssd1 vccd1 vccd1 _09305_/CLK sky130_fd_sc_hd__dlclkp_1
X_06519_ _06519_/A _06544_/Y vssd1 vssd1 vccd1 vccd1 _13799_/Z sky130_fd_sc_hd__ebufn_2
X_07499_ _07499_/A _07524_/Y vssd1 vssd1 vccd1 vccd1 _13659_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11303__A _13933_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09238_ _13916_/X wr vssd1 vssd1 vccd1 vccd1 _09238_/X sky130_fd_sc_hd__and2_1
X_09169_ _13916_/X vssd1 vssd1 vccd1 vccd1 _09169_/Y sky130_fd_sc_hd__inv_2
XFILLER_182_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11200_ _11230_/CLK line[48] vssd1 vssd1 vccd1 vccd1 _11201_/A sky130_fd_sc_hd__dfxtp_1
X_12180_ _12210_/CLK line[112] vssd1 vssd1 vccd1 vccd1 _12181_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_MUX.M\[3\].MUX\[0\]_A3 _13889_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11131_ _11131_/A _11164_/Y vssd1 vssd1 vccd1 vccd1 _13651_/Z sky130_fd_sc_hd__ebufn_2
X_11062_ _11090_/CLK line[122] vssd1 vssd1 vccd1 vccd1 _11063_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[7\].VALID\[9\].FF OVHB\[7\].V/CLK A[16] vssd1 vssd1 vccd1 vccd1 OVHB\[7\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11395__D line[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10013_ _10013_/A _10044_/Y vssd1 vssd1 vccd1 vccd1 _13653_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_49_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06489__D line[65] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[20\].VALID\[1\].FF_D A[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11964_ _11964_/A _11969_/Y vssd1 vssd1 vccd1 vccd1 _13644_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_151_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13703_ _13715_/CLK line[35] vssd1 vssd1 vccd1 vccd1 _13704_/A sky130_fd_sc_hd__dfxtp_1
X_10915_ _10915_/CLK line[41] vssd1 vssd1 vccd1 vccd1 _10916_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_204_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11895_ _11895_/CLK line[105] vssd1 vssd1 vccd1 vccd1 _11896_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[13\].VALID\[5\].FF_D A[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13634_ _13634_/A _13649_/Y vssd1 vssd1 vccd1 vccd1 _13634_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[8\].VALID\[11\].TOBUF OVHB\[8\].VALID\[11\].FF/Q OVHB\[8\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04915_/B2 sky130_fd_sc_hd__ebufn_2
X_10846_ _10846_/A _10849_/Y vssd1 vssd1 vccd1 vccd1 _13646_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07113__D line[109] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_DATA\[23\].CLKBUF\[4\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12954__D line[91] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13565_ _13575_/CLK line[100] vssd1 vssd1 vccd1 vccd1 _13566_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_157_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10777_ _10777_/CLK _10778_/X vssd1 vssd1 vccd1 vccd1 _10775_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__06952__D line[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12516_ _12516_/A _12529_/Y vssd1 vssd1 vccd1 vccd1 _13636_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_12_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13496_ _13496_/A _13509_/Y vssd1 vssd1 vccd1 vccd1 _13776_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_9_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12447_ _12455_/CLK line[101] vssd1 vssd1 vccd1 vccd1 _12448_/A sky130_fd_sc_hd__dfxtp_1
X_12378_ _12378_/A _12389_/Y vssd1 vssd1 vccd1 vccd1 _13778_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13785__D line[73] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11329_ _11335_/CLK line[102] vssd1 vssd1 vccd1 vccd1 _11330_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08879__D line[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07138__A _13909_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06870_ _06890_/CLK line[126] vssd1 vssd1 vccd1 vccd1 _06871_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_94_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[1\].VALID\[10\].TOBUF OVHB\[1\].VALID\[10\].FF/Q OVHB\[1\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04932_/B2 sky130_fd_sc_hd__ebufn_2
X_05821_ _05821_/A _05844_/Y vssd1 vssd1 vccd1 vccd1 _13661_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10499__A _13923_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08540_ _08570_/CLK line[112] vssd1 vssd1 vccd1 vccd1 _08541_/A sky130_fd_sc_hd__dfxtp_1
X_05752_ _05770_/CLK line[127] vssd1 vssd1 vccd1 vccd1 _05753_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[10\].VALID\[6\].TOBUF OVHB\[10\].VALID\[6\].FF/Q OVHB\[10\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04923_/A2 sky130_fd_sc_hd__ebufn_2
XFILLER_208_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09503__D line[35] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08471_ _08471_/A _08504_/Y vssd1 vssd1 vccd1 vccd1 _13791_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_211_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05683_ _05683_/A _05704_/Y vssd1 vssd1 vccd1 vccd1 _13803_/Z sky130_fd_sc_hd__ebufn_2
X_07422_ _07450_/CLK line[122] vssd1 vssd1 vccd1 vccd1 _07423_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[8\].V OVHB\[8\].V/CLK TIE/HI rst_n vssd1 vssd1 vccd1 vccd1 OVHB\[8\].V/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_195_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07353_ _07353_/A _07384_/Y vssd1 vssd1 vccd1 vccd1 _13793_/Z sky130_fd_sc_hd__ebufn_2
X_06304_ _06330_/CLK line[123] vssd1 vssd1 vccd1 vccd1 _06305_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06862__D line[122] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07284_ _07310_/CLK line[59] vssd1 vssd1 vccd1 vccd1 _07285_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_191_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09023_ _09025_/CLK line[72] vssd1 vssd1 vccd1 vccd1 _09024_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10384__D line[54] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06235_ _06235_/A _06264_/Y vssd1 vssd1 vccd1 vccd1 _13795_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05478__D line[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06166_ _06190_/CLK line[60] vssd1 vssd1 vccd1 vccd1 _06167_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13695__D line[46] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[23\].VALID\[14\].FF OVHB\[23\].V/CLK A[21] vssd1 vssd1 vccd1 vccd1 OVHB\[23\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_05117_ _05117_/A _05144_/Y vssd1 vssd1 vccd1 vccd1 _13797_/Z sky130_fd_sc_hd__ebufn_2
X_06097_ _06097_/A _06124_/Y vssd1 vssd1 vccd1 vccd1 _13657_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08789__D line[107] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07693__D line[104] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05048_ _05070_/CLK line[61] vssd1 vssd1 vccd1 vccd1 _05049_/A sky130_fd_sc_hd__dfxtp_1
X_09925_ _09935_/CLK line[100] vssd1 vssd1 vccd1 vccd1 _09926_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_172_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11793__A _13927_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09856_ _09856_/A _09869_/Y vssd1 vssd1 vccd1 vccd1 _13776_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_112_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XOVHB\[31\].V OVHB\[31\].V/CLK TIE/HI rst_n vssd1 vssd1 vccd1 vccd1 OVHB\[31\].V/Q
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06102__D line[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08807_ _08815_/CLK line[101] vssd1 vssd1 vccd1 vccd1 _08808_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[16\].VALID\[1\].FF OVHB\[16\].V/CLK A[8] vssd1 vssd1 vccd1 vccd1 OVHB\[16\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_46_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09787_ _09795_/CLK line[37] vssd1 vssd1 vccd1 vccd1 _09788_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_45_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11943__D line[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06999_ _13909_/Y vssd1 vssd1 vccd1 vccd1 _06999_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08738_ _08738_/A _08749_/Y vssd1 vssd1 vccd1 vccd1 _13778_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[26\].VALID\[5\].FF_D A[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05941__D line[71] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10559__D line[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08669_ _08675_/CLK line[38] vssd1 vssd1 vccd1 vccd1 _08670_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_14_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10700_ _10700_/A _10709_/Y vssd1 vssd1 vccd1 vccd1 _13780_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08029__D line[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ _11680_/A _11689_/Y vssd1 vssd1 vccd1 vccd1 _13640_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10631_ _10635_/CLK line[39] vssd1 vssd1 vccd1 vccd1 _10632_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07868__D line[56] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[19\].VALID\[9\].FF_D A[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13350_ _13350_/A _13369_/Y vssd1 vssd1 vccd1 vccd1 _13630_/Z sky130_fd_sc_hd__ebufn_2
X_10562_ _10562_/A _10569_/Y vssd1 vssd1 vccd1 vccd1 _13642_/Z sky130_fd_sc_hd__ebufn_2
X_12301_ _12315_/CLK line[34] vssd1 vssd1 vccd1 vccd1 _12302_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11968__A _13934_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10294__D line[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13281_ _13295_/CLK line[98] vssd1 vssd1 vccd1 vccd1 _13282_/A sky130_fd_sc_hd__dfxtp_1
X_10493_ _10495_/CLK line[104] vssd1 vssd1 vccd1 vccd1 _10494_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_182_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12232_ _12232_/A _12249_/Y vssd1 vssd1 vccd1 vccd1 _13632_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_6_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_OVHB\[31\].CG_CLK clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12163_ _12175_/CLK line[99] vssd1 vssd1 vccd1 vccd1 _12164_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[19\].VALID\[1\].TOBUF OVHB\[19\].VALID\[1\].FF/Q OVHB\[19\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04926_/B2 sky130_fd_sc_hd__ebufn_2
X_11114_ _11114_/A _11129_/Y vssd1 vssd1 vccd1 vccd1 _13634_/Z sky130_fd_sc_hd__ebufn_2
X_12094_ _12094_/A _12109_/Y vssd1 vssd1 vccd1 vccd1 _13774_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.M\[2\].MUX\[1\]_A1 _13735_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11045_ _11055_/CLK line[100] vssd1 vssd1 vccd1 vccd1 _11046_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[22\].V OVHB\[22\].V/CLK TIE/HI rst_n vssd1 vssd1 vccd1 vccd1 OVHB\[22\].V/Q
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_39_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__04924__B2 _04924_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05851__D line[44] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12996_ _12996_/A _13019_/Y vssd1 vssd1 vccd1 vccd1 _13836_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[24\].VALID\[12\].TOBUF OVHB\[24\].VALID\[12\].FF/Q OVHB\[24\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04929_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__10469__D line[107] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11947_ _11965_/CLK line[15] vssd1 vssd1 vccd1 vccd1 _11948_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_17_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11878_ _11878_/A _11899_/Y vssd1 vssd1 vccd1 vccd1 _13838_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[14\].VALID\[3\].FF OVHB\[14\].V/CLK A[10] vssd1 vssd1 vccd1 vccd1 OVHB\[14\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_13617_ _13645_/CLK line[10] vssd1 vssd1 vccd1 vccd1 _13618_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12684__D line[81] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10829_ _10845_/CLK line[1] vssd1 vssd1 vccd1 vccd1 _10830_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07778__D line[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12039__A _13934_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[31\].VALID\[7\].FF OVHB\[31\].V/CLK A[14] vssd1 vssd1 vccd1 vccd1 OVHB\[31\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_13548_ _13548_/A _13579_/Y vssd1 vssd1 vccd1 vccd1 _13828_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[7\].VALID\[0\].FF_D A[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13479_ _13505_/CLK line[75] vssd1 vssd1 vccd1 vccd1 _13480_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09993__D line[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06020_ _06050_/CLK line[112] vssd1 vssd1 vccd1 vccd1 _06021_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_133_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_DATA\[21\].CLKBUF\[6\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10932__D line[63] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08402__D line[58] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07971_ _07975_/CLK line[103] vssd1 vssd1 vccd1 vccd1 _07972_/A sky130_fd_sc_hd__dfxtp_1
X_09710_ _09710_/A _09729_/Y vssd1 vssd1 vccd1 vccd1 _13630_/Z sky130_fd_sc_hd__ebufn_2
X_06922_ _06922_/A _06929_/Y vssd1 vssd1 vccd1 vccd1 _13642_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_101_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07018__D line[51] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[13\].V OVHB\[13\].V/CLK TIE/HI rst_n vssd1 vssd1 vccd1 vccd1 OVHB\[13\].V/Q
+ sky130_fd_sc_hd__dfrtp_1
X_09641_ _09655_/CLK line[98] vssd1 vssd1 vccd1 vccd1 _09642_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12859__D line[33] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06853_ _06855_/CLK line[104] vssd1 vssd1 vccd1 vccd1 _06854_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_27_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05804_ _05804_/A _05809_/Y vssd1 vssd1 vccd1 vccd1 _13644_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_27_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09572_ _09572_/A _09589_/Y vssd1 vssd1 vccd1 vccd1 _13772_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[25\].VALID\[0\].TOBUF OVHB\[25\].VALID\[0\].FF/Q OVHB\[25\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04924_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__04915__B2 _04915_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06784_ _06784_/A _06789_/Y vssd1 vssd1 vccd1 vccd1 _13784_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09233__D line[40] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08523_ _08535_/CLK line[99] vssd1 vssd1 vccd1 vccd1 _08524_/A sky130_fd_sc_hd__dfxtp_1
X_05735_ _05735_/CLK line[105] vssd1 vssd1 vccd1 vccd1 _05736_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_36_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13333__A _13938_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08454_ _08454_/A _08469_/Y vssd1 vssd1 vccd1 vccd1 _13774_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05666_ _05666_/A _05669_/Y vssd1 vssd1 vccd1 vccd1 _13786_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07405_ _07415_/CLK line[100] vssd1 vssd1 vccd1 vccd1 _07406_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_168_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08385_ _08395_/CLK line[36] vssd1 vssd1 vccd1 vccd1 _08386_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05597_ _05597_/CLK _05598_/X vssd1 vssd1 vccd1 vccd1 _05595_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_211_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06592__D line[127] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07336_ _07336_/A _07349_/Y vssd1 vssd1 vccd1 vccd1 _13776_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_176_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07267_ _07275_/CLK line[37] vssd1 vssd1 vccd1 vccd1 _07268_/A sky130_fd_sc_hd__dfxtp_1
X_09006_ _09006_/A _09029_/Y vssd1 vssd1 vccd1 vccd1 _13766_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[12\].VALID\[5\].FF OVHB\[12\].V/CLK A[12] vssd1 vssd1 vccd1 vccd1 OVHB\[12\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_06218_ _06218_/A _06229_/Y vssd1 vssd1 vccd1 vccd1 _13778_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_136_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07198_ _07198_/A _07209_/Y vssd1 vssd1 vccd1 vccd1 _13638_/Z sky130_fd_sc_hd__ebufn_2
X_06149_ _06155_/CLK line[38] vssd1 vssd1 vccd1 vccd1 _06150_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_117_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09408__D line[120] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13508__A _13898_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09908_ _09908_/A _09939_/Y vssd1 vssd1 vccd1 vccd1 _13828_/Z sky130_fd_sc_hd__ebufn_2
X_09839_ _09865_/CLK line[75] vssd1 vssd1 vccd1 vccd1 _09840_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_58_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11673__D line[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06767__D line[79] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12850_ _12850_/A _12879_/Y vssd1 vssd1 vccd1 vccd1 _13690_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09143__D line[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11801_ _11825_/CLK line[76] vssd1 vssd1 vccd1 vccd1 _11802_/A sky130_fd_sc_hd__dfxtp_1
X_12781_ _12805_/CLK line[12] vssd1 vssd1 vccd1 vccd1 _12782_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08982__D line[53] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11732_ _11732_/A _11759_/Y vssd1 vssd1 vccd1 vccd1 _13692_/Z sky130_fd_sc_hd__ebufn_2
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[17\].VALID\[6\].TOBUF OVHB\[17\].VALID\[6\].FF/Q OVHB\[17\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04923_/A2 sky130_fd_sc_hd__ebufn_2
XPHY_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11663_ _11685_/CLK line[13] vssd1 vssd1 vccd1 vccd1 _11664_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13402_ _13402_/CLK _13403_/X vssd1 vssd1 vccd1 vccd1 _13400_/CLK sky130_fd_sc_hd__dlclkp_1
XPHY_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10614_ _10614_/A _10639_/Y vssd1 vssd1 vccd1 vccd1 _13694_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11594_ _11594_/A _11619_/Y vssd1 vssd1 vccd1 vccd1 _13834_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13333_ _13938_/X wr vssd1 vssd1 vccd1 vccd1 _13333_/X sky130_fd_sc_hd__and2_1
X_10545_ _10565_/CLK line[14] vssd1 vssd1 vccd1 vccd1 _10546_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12009__D line[43] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__04924__A2_N _04924_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09168__A _13916_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06007__D line[101] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13264_ _13938_/X vssd1 vssd1 vccd1 vccd1 _13264_/Y sky130_fd_sc_hd__inv_2
X_10476_ _10476_/A _10499_/Y vssd1 vssd1 vccd1 vccd1 _13836_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11848__D line[83] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12215_ _12245_/CLK line[0] vssd1 vssd1 vccd1 vccd1 _12216_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_108_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13195_ _13225_/CLK line[64] vssd1 vssd1 vccd1 vccd1 _13196_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[0\].VALID\[13\].FF_D A[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09318__D line[93] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12146_ _12146_/A _12179_/Y vssd1 vssd1 vccd1 vccd1 _13826_/Z sky130_fd_sc_hd__ebufn_2
X_12077_ _12105_/CLK line[74] vssd1 vssd1 vccd1 vccd1 _12078_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[10\].VALID\[7\].FF OVHB\[10\].V/CLK A[14] vssd1 vssd1 vccd1 vccd1 OVHB\[10\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_49_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11028_ _11028_/A _11059_/Y vssd1 vssd1 vccd1 vccd1 _13828_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_2_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05581__D line[34] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10199__D line[97] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12979_ _12979_/A _12984_/Y vssd1 vssd1 vccd1 vccd1 _13819_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_18_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05520_ _05520_/A _05529_/Y vssd1 vssd1 vccd1 vccd1 _13640_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08892__D line[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[13\].V_RESET_B rst_n vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05451_ _05455_/CLK line[103] vssd1 vssd1 vccd1 vccd1 _05452_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_20_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08170_ _08170_/A _08189_/Y vssd1 vssd1 vccd1 vccd1 _13770_/Z sky130_fd_sc_hd__ebufn_2
X_05382_ _05382_/A _05389_/Y vssd1 vssd1 vccd1 vccd1 _13782_/Z sky130_fd_sc_hd__ebufn_2
X_07121_ _07135_/CLK line[98] vssd1 vssd1 vccd1 vccd1 _07122_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_146_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07052_ _07052_/A _07069_/Y vssd1 vssd1 vccd1 vccd1 _13772_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[23\].VALID\[5\].TOBUF OVHB\[23\].VALID\[5\].FF/Q OVHB\[23\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04927_/B2 sky130_fd_sc_hd__ebufn_2
X_06003_ _06015_/CLK line[99] vssd1 vssd1 vccd1 vccd1 _06004_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10662__D line[53] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05756__D line[114] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08132__D line[63] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07954_ _07954_/A _07979_/Y vssd1 vssd1 vccd1 vccd1 _13834_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_68_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07971__D line[103] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06905_ _06925_/CLK line[14] vssd1 vssd1 vccd1 vccd1 _06906_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12589__D line[38] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07885_ _07905_/CLK line[78] vssd1 vssd1 vccd1 vccd1 _07886_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[22\].VALID\[8\].FF_D A[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09624_ _13920_/Y vssd1 vssd1 vccd1 vccd1 _09624_/Y sky130_fd_sc_hd__inv_2
X_06836_ _06836_/A _06859_/Y vssd1 vssd1 vccd1 vccd1 _13836_/Z sky130_fd_sc_hd__ebufn_2
X_09555_ _09585_/CLK line[64] vssd1 vssd1 vccd1 vccd1 _09556_/A sky130_fd_sc_hd__dfxtp_1
X_06767_ _06785_/CLK line[79] vssd1 vssd1 vccd1 vccd1 _06768_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09898__D line[88] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08506_ _08506_/A _08539_/Y vssd1 vssd1 vccd1 vccd1 _13826_/Z sky130_fd_sc_hd__ebufn_2
XPHY_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05718_ _05718_/A _05739_/Y vssd1 vssd1 vccd1 vccd1 _13838_/Z sky130_fd_sc_hd__ebufn_2
XPHY_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09486_ _09486_/A _09519_/Y vssd1 vssd1 vccd1 vccd1 _13686_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06698_ _06698_/A _06719_/Y vssd1 vssd1 vccd1 vccd1 _13698_/Z sky130_fd_sc_hd__ebufn_2
XPHY_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10837__D line[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08437_ _08465_/CLK line[74] vssd1 vssd1 vccd1 vccd1 _08438_/A sky130_fd_sc_hd__dfxtp_1
X_05649_ _05665_/CLK line[65] vssd1 vssd1 vccd1 vccd1 _05650_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13213__D line[67] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08307__D line[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08368_ _08368_/A _08399_/Y vssd1 vssd1 vccd1 vccd1 _13688_/Z sky130_fd_sc_hd__ebufn_2
XDECH.DEC0.AND1 A_h[4] A_h[3] vssd1 vssd1 vccd1 vccd1 _13949_/D sky130_fd_sc_hd__and2b_2
XFILLER_137_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07319_ _07345_/CLK line[75] vssd1 vssd1 vccd1 vccd1 _07320_/A sky130_fd_sc_hd__dfxtp_1
X_08299_ _08325_/CLK line[11] vssd1 vssd1 vccd1 vccd1 _08300_/A sky130_fd_sc_hd__dfxtp_1
X_10330_ _10330_/A _10359_/Y vssd1 vssd1 vccd1 vccd1 _13690_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10572__D line[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10261_ _10285_/CLK line[12] vssd1 vssd1 vccd1 vccd1 _10262_/A sky130_fd_sc_hd__dfxtp_1
X_12000_ _12000_/CLK line[25] vssd1 vssd1 vccd1 vccd1 _12001_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[0\].CGAND _13931_/Y wr vssd1 vssd1 vccd1 vccd1 OVHB\[0\].CGAND/X sky130_fd_sc_hd__and2_4
XFILLER_133_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10192_ _10192_/A _10219_/Y vssd1 vssd1 vccd1 vccd1 _13832_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07881__D line[76] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12499__D line[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13951_ A_h[1] vssd1 vssd1 vccd1 vccd1 _13960_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_86_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06497__D line[69] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12902_ _12910_/CLK line[53] vssd1 vssd1 vccd1 vccd1 _12903_/A sky130_fd_sc_hd__dfxtp_1
X_13882_ _13890_/CLK line[117] vssd1 vssd1 vccd1 vccd1 _13883_/A sky130_fd_sc_hd__dfxtp_1
X_12833_ _12833_/A _12844_/Y vssd1 vssd1 vccd1 vccd1 _13673_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_34_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12764_ _12770_/CLK line[118] vssd1 vssd1 vccd1 vccd1 _12765_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11715_ _11715_/A _11724_/Y vssd1 vssd1 vccd1 vccd1 _13675_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_70_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10747__D line[106] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12695_ _12695_/A _12704_/Y vssd1 vssd1 vccd1 vccd1 _13815_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[3\].VALID\[3\].FF_D A[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11646_ _11650_/CLK line[119] vssd1 vssd1 vccd1 vccd1 _11647_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07121__D line[98] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12962__D line[95] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11577_ _11577_/A _11584_/Y vssd1 vssd1 vccd1 vccd1 _13817_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06960__D line[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13316_ _13330_/CLK line[114] vssd1 vssd1 vccd1 vccd1 _13317_/A sky130_fd_sc_hd__dfxtp_1
X_10528_ _10530_/CLK line[120] vssd1 vssd1 vccd1 vccd1 _10529_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11578__D line[88] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13247_ _13247_/A _13264_/Y vssd1 vssd1 vccd1 vccd1 _13807_/Z sky130_fd_sc_hd__ebufn_2
X_10459_ _10459_/A _10464_/Y vssd1 vssd1 vccd1 vccd1 _13819_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09048__D line[83] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13178_ _13190_/CLK line[51] vssd1 vssd1 vccd1 vccd1 _13179_/A sky130_fd_sc_hd__dfxtp_1
X_12129_ _12129_/A _12144_/Y vssd1 vssd1 vccd1 vccd1 _13809_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_04951_ _04965_/CLK line[2] vssd1 vssd1 vccd1 vccd1 _04952_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[3\].VALID\[0\].FF OVHB\[3\].V/CLK A[7] vssd1 vssd1 vccd1 vccd1 OVHB\[3\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_37_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_DATA\[14\].CLKBUF\[0\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12202__D line[117] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07670_ _07670_/A _07699_/Y vssd1 vssd1 vccd1 vccd1 _13830_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[14\].VALID\[10\].TOBUF OVHB\[14\].VALID\[10\].FF/Q OVHB\[14\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04932_/B2 sky130_fd_sc_hd__ebufn_2
X_06621_ _06645_/CLK line[12] vssd1 vssd1 vccd1 vccd1 _06622_/A sky130_fd_sc_hd__dfxtp_1
X_09340_ _09340_/CLK line[89] vssd1 vssd1 vccd1 vccd1 _09341_/A sky130_fd_sc_hd__dfxtp_1
X_06552_ _06552_/A _06579_/Y vssd1 vssd1 vccd1 vccd1 _13832_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09511__D line[39] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05503_ _05525_/CLK line[13] vssd1 vssd1 vccd1 vccd1 _05504_/A sky130_fd_sc_hd__dfxtp_1
X_09271_ _09271_/A _09274_/Y vssd1 vssd1 vccd1 vccd1 _13751_/Z sky130_fd_sc_hd__ebufn_2
X_06483_ _06505_/CLK line[77] vssd1 vssd1 vccd1 vccd1 _06484_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_20_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08222_ _08222_/CLK _08223_/X vssd1 vssd1 vccd1 vccd1 _08220_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_138_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05434_ _05434_/A _05459_/Y vssd1 vssd1 vccd1 vccd1 _13834_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_119_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XOVHB\[28\].VALID\[14\].FF OVHB\[28\].V/CLK A[21] vssd1 vssd1 vccd1 vccd1 OVHB\[28\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_08153_ _13932_/X wr vssd1 vssd1 vccd1 vccd1 _08153_/X sky130_fd_sc_hd__and2_1
X_05365_ _05385_/CLK line[78] vssd1 vssd1 vccd1 vccd1 _05366_/A sky130_fd_sc_hd__dfxtp_1
X_07104_ _13909_/Y vssd1 vssd1 vccd1 vccd1 _07104_/Y sky130_fd_sc_hd__inv_2
XANTENNA__06870__D line[126] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08084_ _13932_/X vssd1 vssd1 vccd1 vccd1 _08084_/Y sky130_fd_sc_hd__inv_2
XANTENNA_DATA\[7\].CLKBUF\[0\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05296_ _05296_/A _05319_/Y vssd1 vssd1 vccd1 vccd1 _13696_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11488__D line[61] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07035_ _07065_/CLK line[64] vssd1 vssd1 vccd1 vccd1 _07036_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_161_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05486__D line[119] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[18\].VALID\[0\].FF_D A[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08797__D line[111] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08986_ _08990_/CLK line[55] vssd1 vssd1 vccd1 vccd1 _08987_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[7\].VALID\[13\].FF_D A[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07937_ _07937_/A _07944_/Y vssd1 vssd1 vccd1 vccd1 _13817_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_28_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12112__D line[90] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07868_ _07870_/CLK line[56] vssd1 vssd1 vccd1 vccd1 _07869_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06110__D line[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09607_ _09607_/A _09624_/Y vssd1 vssd1 vccd1 vccd1 _13807_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_28_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06819_ _06819_/A _06824_/Y vssd1 vssd1 vccd1 vccd1 _13819_/Z sky130_fd_sc_hd__ebufn_2
X_07799_ _07799_/A _07804_/Y vssd1 vssd1 vccd1 vccd1 _13679_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11951__D line[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09538_ _09550_/CLK line[51] vssd1 vssd1 vccd1 vccd1 _09539_/A sky130_fd_sc_hd__dfxtp_1
XPHY_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09421__D line[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[1\].VALID\[2\].FF OVHB\[1\].V/CLK A[9] vssd1 vssd1 vccd1 vccd1 OVHB\[1\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09469_ _09469_/A _09484_/Y vssd1 vssd1 vccd1 vccd1 _13669_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11500_ _11510_/CLK line[52] vssd1 vssd1 vccd1 vccd1 _11501_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_157_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08037__D line[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12480_ _12490_/CLK line[116] vssd1 vssd1 vccd1 vccd1 _12481_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13878__D line[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11431_ _11431_/A _11444_/Y vssd1 vssd1 vccd1 vccd1 _13671_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_22_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_MUX.M\[3\].MUX\[3\]_A1 _13725_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[9\].VALID\[7\].FF_D A[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11362_ _11370_/CLK line[117] vssd1 vssd1 vccd1 vccd1 _11363_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_164_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13101_ _13101_/A _13124_/Y vssd1 vssd1 vccd1 vccd1 _13661_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_137_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10313_ _10313_/A _10324_/Y vssd1 vssd1 vccd1 vccd1 _13673_/Z sky130_fd_sc_hd__ebufn_2
X_11293_ _11293_/A _11304_/Y vssd1 vssd1 vccd1 vccd1 _13813_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[5\].VALID\[2\].TOBUF OVHB\[5\].VALID\[2\].FF/Q OVHB\[5\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04930_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__05396__D line[92] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13032_ _13050_/CLK line[127] vssd1 vssd1 vccd1 vccd1 _13033_/A sky130_fd_sc_hd__dfxtp_1
X_10244_ _10250_/CLK line[118] vssd1 vssd1 vccd1 vccd1 _10245_/A sky130_fd_sc_hd__dfxtp_1
X_10175_ _10175_/A _10184_/Y vssd1 vssd1 vccd1 vccd1 _13815_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08500__D line[89] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13118__D line[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13934_ _13938_/C _13938_/B _13938_/A _13938_/D vssd1 vssd1 vccd1 vccd1 _13934_/X
+ sky130_fd_sc_hd__and4b_4
XFILLER_47_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[5\].CG_CLK clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06020__D line[112] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13865_ _13865_/A _13894_/Y vssd1 vssd1 vccd1 vccd1 _13865_/Z sky130_fd_sc_hd__ebufn_2
X_12816_ _12840_/CLK line[28] vssd1 vssd1 vccd1 vccd1 _12817_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_15_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13796_ _13820_/CLK line[92] vssd1 vssd1 vccd1 vccd1 _13797_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05214__A _13931_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10477__D line[111] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12747_ _12747_/A _12774_/Y vssd1 vssd1 vccd1 vccd1 _13867_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_63_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12678_ _12700_/CLK line[93] vssd1 vssd1 vccd1 vccd1 _12679_/A sky130_fd_sc_hd__dfxtp_1
XPHY_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12692__D line[85] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11629_ _11629_/A _11654_/Y vssd1 vssd1 vccd1 vccd1 _13869_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_8_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07786__D line[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05150_ _05150_/A _05179_/Y vssd1 vssd1 vccd1 vccd1 _13830_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_190_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05081_ _05105_/CLK line[76] vssd1 vssd1 vccd1 vccd1 _05082_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11101__D line[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10940__D line[52] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08840_ _08850_/CLK line[116] vssd1 vssd1 vccd1 vccd1 _08841_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_85_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08410__D line[62] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[0\].VALID\[14\].FF OVHB\[0\].V/CLK A[21] vssd1 vssd1 vccd1 vccd1 OVHB\[0\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_97_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08771_ _08771_/A _08784_/Y vssd1 vssd1 vccd1 vccd1 _13811_/Z sky130_fd_sc_hd__ebufn_2
X_05983_ _13902_/X wr vssd1 vssd1 vccd1 vccd1 _05983_/X sky130_fd_sc_hd__and2_1
XFILLER_66_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13028__D line[125] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07722_ _07730_/CLK line[117] vssd1 vssd1 vccd1 vccd1 _07723_/A sky130_fd_sc_hd__dfxtp_1
X_04934_ _04934_/A _04934_/B _04934_/C _04934_/D vssd1 vssd1 vccd1 vccd1 hit sky130_fd_sc_hd__nor4_2
XFILLER_38_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05108__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07026__D line[55] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12867__D line[37] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07653_ _07653_/A _07664_/Y vssd1 vssd1 vccd1 vccd1 _13813_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_65_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06604_ _06610_/CLK line[118] vssd1 vssd1 vccd1 vccd1 _06605_/A sky130_fd_sc_hd__dfxtp_1
X_07584_ _07590_/CLK line[54] vssd1 vssd1 vccd1 vccd1 _07585_/A sky130_fd_sc_hd__dfxtp_1
X_09323_ _09323_/A _09344_/Y vssd1 vssd1 vccd1 vccd1 _13803_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_34_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06535_ _06535_/A _06544_/Y vssd1 vssd1 vccd1 vccd1 _13815_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[12\].CLKBUF\[2\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09254_ _09270_/CLK line[49] vssd1 vssd1 vccd1 vccd1 _09255_/A sky130_fd_sc_hd__dfxtp_1
X_06466_ _06470_/CLK line[55] vssd1 vssd1 vccd1 vccd1 _06467_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_166_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08205_ _08205_/A _08224_/Y vssd1 vssd1 vccd1 vccd1 _13805_/Z sky130_fd_sc_hd__ebufn_2
X_05417_ _05417_/A _05424_/Y vssd1 vssd1 vccd1 vccd1 _13817_/Z sky130_fd_sc_hd__ebufn_2
X_09185_ _09185_/A _09204_/Y vssd1 vssd1 vccd1 vccd1 _13665_/Z sky130_fd_sc_hd__ebufn_2
X_06397_ _06397_/A _06404_/Y vssd1 vssd1 vccd1 vccd1 _13677_/Z sky130_fd_sc_hd__ebufn_2
X_08136_ _08150_/CLK line[50] vssd1 vssd1 vccd1 vccd1 _08137_/A sky130_fd_sc_hd__dfxtp_1
X_05348_ _05350_/CLK line[56] vssd1 vssd1 vccd1 vccd1 _05349_/A sky130_fd_sc_hd__dfxtp_1
X_08067_ _08067_/A _08084_/Y vssd1 vssd1 vccd1 vccd1 _13667_/Z sky130_fd_sc_hd__ebufn_2
X_05279_ _05279_/A _05284_/Y vssd1 vssd1 vccd1 vccd1 _13679_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_162_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07018_ _07030_/CLK line[51] vssd1 vssd1 vccd1 vccd1 _07019_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_68_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10850__D line[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_DATA\[5\].CLKBUF\[2\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08969_ _08969_/A _08994_/Y vssd1 vssd1 vccd1 vccd1 _13729_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_124_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11980_ _12000_/CLK line[30] vssd1 vssd1 vccd1 vccd1 _11981_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_124_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10931_ _10931_/A _10954_/Y vssd1 vssd1 vccd1 vccd1 _13731_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[31\].CLKBUF\[4\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[4\].CGAND_B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[24\].VALID\[12\].FF OVHB\[24\].V/CLK A[19] vssd1 vssd1 vccd1 vccd1 OVHB\[24\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12777__D line[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[23\].CGAND_A _13916_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11681__D line[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06775__D line[68] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10862_ _10880_/CLK line[31] vssd1 vssd1 vccd1 vccd1 _10863_/A sky130_fd_sc_hd__dfxtp_1
X_13650_ _13680_/CLK line[16] vssd1 vssd1 vccd1 vccd1 _13651_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_140_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09151__D line[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[3\].VALID\[7\].TOBUF OVHB\[3\].VALID\[7\].FF/Q OVHB\[3\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/A2 sky130_fd_sc_hd__ebufn_2
XFILLER_71_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12601_ _12601_/A _12634_/Y vssd1 vssd1 vccd1 vccd1 _13721_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[8\].CGAND_A _13898_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13581_ _13581_/A _13614_/Y vssd1 vssd1 vccd1 vccd1 _13861_/Z sky130_fd_sc_hd__ebufn_2
X_10793_ _10793_/A _10814_/Y vssd1 vssd1 vccd1 vccd1 _13873_/Z sky130_fd_sc_hd__ebufn_2
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12532_ _12560_/CLK line[26] vssd1 vssd1 vccd1 vccd1 _12533_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08990__D line[57] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12463_ _12463_/A _12494_/Y vssd1 vssd1 vccd1 vccd1 _13863_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_200_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11414_ _11440_/CLK line[27] vssd1 vssd1 vccd1 vccd1 _11415_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09057__TE_B _09064_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12394_ _12420_/CLK line[91] vssd1 vssd1 vccd1 vccd1 _12395_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12017__D line[47] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11345_ _11345_/A _11374_/Y vssd1 vssd1 vccd1 vccd1 _13865_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_153_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06015__D line[105] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11276_ _11300_/CLK line[92] vssd1 vssd1 vccd1 vccd1 _11277_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_180_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11856__D line[87] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[14\].VALID\[14\].FF OVHB\[14\].V/CLK A[21] vssd1 vssd1 vccd1 vccd1 OVHB\[14\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_13015_ _13015_/CLK line[105] vssd1 vssd1 vccd1 vccd1 _13016_/A sky130_fd_sc_hd__dfxtp_1
X_10227_ _10227_/A _10254_/Y vssd1 vssd1 vccd1 vccd1 _13867_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09326__D line[82] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09904__A _13921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10158_ _10180_/CLK line[93] vssd1 vssd1 vccd1 vccd1 _10159_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09623__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10089_ _10089_/A _10114_/Y vssd1 vssd1 vccd1 vccd1 _13729_/Z sky130_fd_sc_hd__ebufn_2
X_13917_ A[2] vssd1 vssd1 vccd1 vccd1 _13927_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_208_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11591__D line[108] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06685__D line[32] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13848_ _13848_/A _13859_/Y vssd1 vssd1 vccd1 vccd1 _13848_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_16_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13779_ _13785_/CLK line[70] vssd1 vssd1 vccd1 vccd1 _13780_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MUX.M\[0\].MUX\[0\]_A0 _13616_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06320_ _06330_/CLK line[116] vssd1 vssd1 vccd1 vccd1 _06321_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05879__A _13902_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05598__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06251_ _06251_/A _06264_/Y vssd1 vssd1 vccd1 vccd1 _13811_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[29\].CLKBUF\[0\] clk vssd1 vssd1 vccd1 vccd1 _10847_/CLK sky130_fd_sc_hd__clkbuf_4
X_05202_ _05210_/CLK line[117] vssd1 vssd1 vccd1 vccd1 _05203_/A sky130_fd_sc_hd__dfxtp_1
X_06182_ _06190_/CLK line[53] vssd1 vssd1 vccd1 vccd1 _06183_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_116_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[10\].VALID\[2\].TOBUF OVHB\[10\].VALID\[2\].FF/Q OVHB\[10\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04930_/B2 sky130_fd_sc_hd__ebufn_2
XDATA\[19\].CLKBUF\[6\] clk vssd1 vssd1 vccd1 vccd1 _07977_/CLK sky130_fd_sc_hd__clkbuf_4
X_05133_ _05133_/A _05144_/Y vssd1 vssd1 vccd1 vccd1 _13813_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[14\].VALID\[3\].FF_D A[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XOVHB\[24\].VALID\[1\].FF OVHB\[24\].V/CLK A[8] vssd1 vssd1 vccd1 vccd1 OVHB\[24\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_09941_ _09941_/A _09974_/Y vssd1 vssd1 vccd1 vccd1 _13861_/Z sky130_fd_sc_hd__ebufn_2
X_05064_ _05070_/CLK line[54] vssd1 vssd1 vccd1 vccd1 _05065_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11766__D line[60] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10670__D line[57] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09872_ _09900_/CLK line[90] vssd1 vssd1 vccd1 vccd1 _09873_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_97_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05764__D line[118] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08140__D line[52] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08823_ _08823_/A _08854_/Y vssd1 vssd1 vccd1 vccd1 _13863_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_57_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08754_ _08780_/CLK line[91] vssd1 vssd1 vccd1 vccd1 _08755_/A sky130_fd_sc_hd__dfxtp_1
X_05966_ _05980_/CLK line[82] vssd1 vssd1 vccd1 vccd1 _05967_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_72_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07705_ _07705_/A _07734_/Y vssd1 vssd1 vccd1 vccd1 _13865_/Z sky130_fd_sc_hd__ebufn_2
X_04917_ _04917_/A _04917_/B _04917_/C _04917_/D vssd1 vssd1 vccd1 vccd1 _04934_/A
+ sky130_fd_sc_hd__or4_2
X_08685_ _08685_/A _08714_/Y vssd1 vssd1 vccd1 vccd1 _13725_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_72_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05897_ _05897_/A _05914_/Y vssd1 vssd1 vccd1 vccd1 _13737_/Z sky130_fd_sc_hd__ebufn_2
X_07636_ _07660_/CLK line[92] vssd1 vssd1 vccd1 vccd1 _07637_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_53_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07567_ _07567_/A _07594_/Y vssd1 vssd1 vccd1 vccd1 _13727_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11006__D line[82] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09306_ _09306_/A _09309_/Y vssd1 vssd1 vccd1 vccd1 _13786_/Z sky130_fd_sc_hd__ebufn_2
X_06518_ _06540_/CLK line[93] vssd1 vssd1 vccd1 vccd1 _06519_/A sky130_fd_sc_hd__dfxtp_1
X_07498_ _07520_/CLK line[29] vssd1 vssd1 vccd1 vccd1 _07499_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10845__D line[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09237_ _09237_/CLK _09238_/X vssd1 vssd1 vccd1 vccd1 _09235_/CLK sky130_fd_sc_hd__dlclkp_1
X_06449_ _06449_/A _06474_/Y vssd1 vssd1 vccd1 vccd1 _13729_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11303__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13221__D line[71] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05939__D line[70] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08315__D line[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09168_ _13916_/X wr vssd1 vssd1 vccd1 vccd1 _09168_/X sky130_fd_sc_hd__and2_1
XANTENNA_DATA\[10\].CLKBUF\[4\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08119_ _13932_/X vssd1 vssd1 vccd1 vccd1 _08119_/Y sky130_fd_sc_hd__inv_2
X_09099_ _13915_/X vssd1 vssd1 vccd1 vccd1 _09099_/Y sky130_fd_sc_hd__inv_2
XFILLER_162_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11130_ _11160_/CLK line[16] vssd1 vssd1 vccd1 vccd1 _11131_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_79_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10580__D line[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11061_ _11061_/A _11094_/Y vssd1 vssd1 vccd1 vccd1 _13861_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[18\].CLKBUF\[3\] clk vssd1 vssd1 vccd1 vccd1 _07592_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_49_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05674__D line[91] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[15\].V_D TIE/HI vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10012_ _10040_/CLK line[26] vssd1 vssd1 vccd1 vccd1 _10013_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_88_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08050__D line[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[4\].VALID\[12\].TOBUF OVHB\[4\].VALID\[12\].FF/Q OVHB\[4\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04929_/B2 sky130_fd_sc_hd__ebufn_2
XOVHB\[22\].VALID\[3\].FF OVHB\[22\].V/CLK A[10] vssd1 vssd1 vccd1 vccd1 OVHB\[22\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_151_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07244__A _13910_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11963_ _11965_/CLK line[8] vssd1 vssd1 vccd1 vccd1 _11964_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_189_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13702_ _13702_/A _13719_/Y vssd1 vssd1 vccd1 vccd1 _13702_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[3\].CLKBUF\[4\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10914_ _10914_/A _10919_/Y vssd1 vssd1 vccd1 vccd1 _13714_/Z sky130_fd_sc_hd__ebufn_2
X_11894_ _11894_/A _11899_/Y vssd1 vssd1 vccd1 vccd1 _13854_/Z sky130_fd_sc_hd__ebufn_2
X_10845_ _10845_/CLK line[9] vssd1 vssd1 vccd1 vccd1 _10846_/A sky130_fd_sc_hd__dfxtp_1
X_13633_ _13645_/CLK line[3] vssd1 vssd1 vccd1 vccd1 _13634_/A sky130_fd_sc_hd__dfxtp_1
X_10776_ _10776_/A _10779_/Y vssd1 vssd1 vccd1 vccd1 _13856_/Z sky130_fd_sc_hd__ebufn_2
X_13564_ _13564_/A _13579_/Y vssd1 vssd1 vccd1 vccd1 _13844_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10755__D line[110] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12515_ _12525_/CLK line[4] vssd1 vssd1 vccd1 vccd1 _12516_/A sky130_fd_sc_hd__dfxtp_1
X_13495_ _13505_/CLK line[68] vssd1 vssd1 vccd1 vccd1 _13496_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_12_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13131__D line[44] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[27\].VALID\[3\].FF_D A[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05849__D line[43] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12446_ _12446_/A _12459_/Y vssd1 vssd1 vccd1 vccd1 _13846_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08225__D line[96] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12970__D line[84] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12377_ _12385_/CLK line[69] vssd1 vssd1 vccd1 vccd1 _12378_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_125_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_OVHB\[24\].VALID\[14\].FF_D A[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11328_ _11328_/A _11339_/Y vssd1 vssd1 vccd1 vccd1 _13848_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07419__A _13910_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07138__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11259_ _11265_/CLK line[70] vssd1 vssd1 vccd1 vccd1 _11260_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[20\].VALID\[10\].FF OVHB\[20\].V/CLK A[17] vssd1 vssd1 vccd1 vccd1 OVHB\[20\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__09056__D line[87] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05820_ _05840_/CLK line[30] vssd1 vssd1 vccd1 vccd1 _05821_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_67_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XDATA\[17\].CLKBUF\[0\] clk vssd1 vssd1 vccd1 vccd1 _07207_/CLK sky130_fd_sc_hd__clkbuf_4
X_05751_ _05751_/A _05774_/Y vssd1 vssd1 vccd1 vccd1 _13871_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13306__D line[124] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12210__D line[121] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08470_ _08500_/CLK line[80] vssd1 vssd1 vccd1 vccd1 _08471_/A sky130_fd_sc_hd__dfxtp_1
X_05682_ _05700_/CLK line[95] vssd1 vssd1 vccd1 vccd1 _05683_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07304__D line[54] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07421_ _07421_/A _07454_/Y vssd1 vssd1 vccd1 vccd1 _13861_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_35_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XOVHB\[20\].VALID\[5\].FF OVHB\[20\].V/CLK A[12] vssd1 vssd1 vccd1 vccd1 OVHB\[20\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_07352_ _07380_/CLK line[90] vssd1 vssd1 vccd1 vccd1 _07353_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_188_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06303_ _06303_/A _06334_/Y vssd1 vssd1 vccd1 vccd1 _13863_/Z sky130_fd_sc_hd__ebufn_2
X_07283_ _07283_/A _07314_/Y vssd1 vssd1 vccd1 vccd1 _13723_/Z sky130_fd_sc_hd__ebufn_2
X_09022_ _09022_/A _09029_/Y vssd1 vssd1 vccd1 vccd1 _13782_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[10\].VALID\[12\].FF OVHB\[10\].V/CLK A[19] vssd1 vssd1 vccd1 vccd1 OVHB\[10\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_06234_ _06260_/CLK line[91] vssd1 vssd1 vccd1 vccd1 _06235_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_136_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08713__A _13914_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12880__D line[48] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06165_ _06165_/A _06194_/Y vssd1 vssd1 vccd1 vccd1 _13725_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_116_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05116_ _05140_/CLK line[92] vssd1 vssd1 vccd1 vccd1 _05117_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_172_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06096_ _06120_/CLK line[28] vssd1 vssd1 vccd1 vccd1 _06097_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11496__D line[50] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[16\].VALID\[11\].FF_D A[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05047_ _05047_/A _05074_/Y vssd1 vssd1 vccd1 vccd1 _13727_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_120_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09924_ _09924_/A _09939_/Y vssd1 vssd1 vccd1 vccd1 _13844_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_86_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11793__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09855_ _09865_/CLK line[68] vssd1 vssd1 vccd1 vccd1 _09856_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_100_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08806_ _08806_/A _08819_/Y vssd1 vssd1 vccd1 vccd1 _13846_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_65_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06998_ _13909_/Y wr vssd1 vssd1 vccd1 vccd1 _06998_/X sky130_fd_sc_hd__and2_1
X_09786_ _09786_/A _09799_/Y vssd1 vssd1 vccd1 vccd1 _13706_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_27_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08737_ _08745_/CLK line[69] vssd1 vssd1 vccd1 vccd1 _08738_/A sky130_fd_sc_hd__dfxtp_1
X_05949_ _13902_/X vssd1 vssd1 vccd1 vccd1 _05949_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12120__D line[94] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[27\].VALID\[14\].TOBUF OVHB\[27\].VALID\[14\].FF/Q OVHB\[27\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/B2 sky130_fd_sc_hd__ebufn_2
X_08668_ _08668_/A _08679_/Y vssd1 vssd1 vccd1 vccd1 _13708_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07214__D line[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XOVHB\[19\].VALID\[6\].FF OVHB\[19\].V/CLK A[13] vssd1 vssd1 vccd1 vccd1 OVHB\[19\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[26\].VALID\[10\].FF_D A[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07619_ _07625_/CLK line[70] vssd1 vssd1 vccd1 vccd1 _07620_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08599_ _08605_/CLK line[6] vssd1 vssd1 vccd1 vccd1 _08600_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[28\].CLKBUF\[7\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10630_ _10630_/A _10639_/Y vssd1 vssd1 vccd1 vccd1 _13710_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10561_ _10565_/CLK line[7] vssd1 vssd1 vccd1 vccd1 _10562_/A sky130_fd_sc_hd__dfxtp_1
X_12300_ _12300_/A _12319_/Y vssd1 vssd1 vccd1 vccd1 _13700_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08045__D line[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13280_ _13280_/A _13299_/Y vssd1 vssd1 vccd1 vccd1 _13840_/Z sky130_fd_sc_hd__ebufn_2
X_10492_ _10492_/A _10499_/Y vssd1 vssd1 vccd1 vccd1 _13852_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11968__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13886__D line[119] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12231_ _12245_/CLK line[2] vssd1 vssd1 vccd1 vccd1 _12232_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_108_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12162_ _12162_/A _12179_/Y vssd1 vssd1 vccd1 vccd1 _13842_/Z sky130_fd_sc_hd__ebufn_2
X_11113_ _11125_/CLK line[3] vssd1 vssd1 vccd1 vccd1 _11114_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[17\].VALID\[2\].TOBUF OVHB\[17\].VALID\[2\].FF/Q OVHB\[17\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04930_/B2 sky130_fd_sc_hd__ebufn_2
X_12093_ _12105_/CLK line[67] vssd1 vssd1 vccd1 vccd1 _12094_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_1_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MUX.M\[2\].MUX\[1\]_A2 _13805_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[20\].VALID\[13\].TOBUF OVHB\[20\].VALID\[13\].FF/Q OVHB\[20\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04916_/B2 sky130_fd_sc_hd__ebufn_2
X_11044_ _11044_/A _11059_/Y vssd1 vssd1 vccd1 vccd1 _13844_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_49_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09604__D line[81] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12995_ _13015_/CLK line[110] vssd1 vssd1 vccd1 vccd1 _12996_/A sky130_fd_sc_hd__dfxtp_1
X_11946_ _11946_/A _11969_/Y vssd1 vssd1 vccd1 vccd1 _13626_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_55_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_OVHB\[12\].V_RESET_B rst_n vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11877_ _11895_/CLK line[111] vssd1 vssd1 vccd1 vccd1 _11878_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_60_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13616_ _13616_/A _13649_/Y vssd1 vssd1 vccd1 vccd1 _13616_/Z sky130_fd_sc_hd__ebufn_2
X_10828_ _10828_/A _10849_/Y vssd1 vssd1 vccd1 vccd1 _13628_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_186_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10485__D line[100] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13547_ _13575_/CLK line[106] vssd1 vssd1 vccd1 vccd1 _13548_/A sky130_fd_sc_hd__dfxtp_1
X_10759_ _10775_/CLK line[97] vssd1 vssd1 vccd1 vccd1 _10760_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[1\].CLKBUF\[6\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05579__D line[33] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[10\].VALID\[6\].FF_D A[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13478_ _13478_/A _13509_/Y vssd1 vssd1 vccd1 vccd1 _13758_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[17\].VALID\[8\].FF OVHB\[17\].V/CLK A[15] vssd1 vssd1 vccd1 vccd1 OVHB\[17\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13796__D line[92] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12429_ _12455_/CLK line[107] vssd1 vssd1 vccd1 vccd1 _12430_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07794__D line[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XOVHB\[5\].VALID\[14\].FF OVHB\[5\].V/CLK A[21] vssd1 vssd1 vccd1 vccd1 OVHB\[5\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_126_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06053__A _13902_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07970_ _07970_/A _07979_/Y vssd1 vssd1 vccd1 vccd1 _13850_/Z sky130_fd_sc_hd__ebufn_2
X_06921_ _06925_/CLK line[7] vssd1 vssd1 vccd1 vccd1 _06922_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06203__D line[77] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[19\].INV _13956_/X vssd1 vssd1 vccd1 vccd1 OVHB\[19\].INV/Y sky130_fd_sc_hd__inv_2
XFILLER_67_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09640_ _09640_/A _09659_/Y vssd1 vssd1 vccd1 vccd1 _13840_/Z sky130_fd_sc_hd__ebufn_2
X_06852_ _06852_/A _06859_/Y vssd1 vssd1 vccd1 vccd1 _13852_/Z sky130_fd_sc_hd__ebufn_2
X_05803_ _05805_/CLK line[8] vssd1 vssd1 vccd1 vccd1 _05804_/A sky130_fd_sc_hd__dfxtp_1
X_09571_ _09585_/CLK line[66] vssd1 vssd1 vccd1 vccd1 _09572_/A sky130_fd_sc_hd__dfxtp_1
X_06783_ _06785_/CLK line[72] vssd1 vssd1 vccd1 vccd1 _06784_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13036__D line[114] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08522_ _08522_/A _08539_/Y vssd1 vssd1 vccd1 vccd1 _13842_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13614__A _13898_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05734_ _05734_/A _05739_/Y vssd1 vssd1 vccd1 vccd1 _13854_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[23\].VALID\[1\].TOBUF OVHB\[23\].VALID\[1\].FF/Q OVHB\[23\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04926_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_23_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08453_ _08465_/CLK line[67] vssd1 vssd1 vccd1 vccd1 _08454_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12875__D line[41] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05665_ _05665_/CLK line[73] vssd1 vssd1 vccd1 vccd1 _05666_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13333__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07404_ _07404_/A _07419_/Y vssd1 vssd1 vccd1 vccd1 _13844_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07969__D line[102] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08384_ _08384_/A _08399_/Y vssd1 vssd1 vccd1 vccd1 _13704_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_149_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05596_ _05596_/A _05599_/Y vssd1 vssd1 vccd1 vccd1 _13716_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06228__A _13903_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07335_ _07345_/CLK line[68] vssd1 vssd1 vccd1 vccd1 _07336_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10395__D line[64] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07266_ _07266_/A _07279_/Y vssd1 vssd1 vccd1 vccd1 _13706_/Z sky130_fd_sc_hd__ebufn_2
X_09005_ _09025_/CLK line[78] vssd1 vssd1 vccd1 vccd1 _09006_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_191_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06217_ _06225_/CLK line[69] vssd1 vssd1 vccd1 vccd1 _06218_/A sky130_fd_sc_hd__dfxtp_1
X_07197_ _07205_/CLK line[5] vssd1 vssd1 vccd1 vccd1 _07198_/A sky130_fd_sc_hd__dfxtp_1
X_06148_ _06148_/A _06159_/Y vssd1 vssd1 vccd1 vccd1 _13708_/Z sky130_fd_sc_hd__ebufn_2
X_06079_ _06085_/CLK line[6] vssd1 vssd1 vccd1 vccd1 _06080_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_132_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[29\].VALID\[12\].FF OVHB\[29\].V/CLK A[19] vssd1 vssd1 vccd1 vccd1 OVHB\[29\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__09274__A _13916_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09907_ _09935_/CLK line[106] vssd1 vssd1 vccd1 vccd1 _09908_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13508__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09838_ _09838_/A _09869_/Y vssd1 vssd1 vccd1 vccd1 _13758_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_59_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05952__D line[90] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[30\].VALID\[2\].FF_D A[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09769_ _09795_/CLK line[43] vssd1 vssd1 vccd1 vccd1 _09770_/A sky130_fd_sc_hd__dfxtp_1
X_11800_ _11800_/A _11829_/Y vssd1 vssd1 vccd1 vccd1 _13760_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[30\].CG clk OVHB\[30\].CGAND/X vssd1 vssd1 vccd1 vccd1 OVHB\[30\].V/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_15_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12780_ _12780_/A _12809_/Y vssd1 vssd1 vccd1 vccd1 _13620_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12785__D line[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11731_ _11755_/CLK line[44] vssd1 vssd1 vccd1 vccd1 _11732_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07879__D line[75] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06783__D line[72] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[15\].VALID\[7\].TOBUF OVHB\[15\].VALID\[7\].FF/Q OVHB\[15\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/A2 sky130_fd_sc_hd__ebufn_2
XPHY_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11662_ _11662_/A _11689_/Y vssd1 vssd1 vccd1 vccd1 _13622_/Z sky130_fd_sc_hd__ebufn_2
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[23\].VALID\[6\].FF_D A[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XMUX.M\[0\].MUX\[1\] _13630_/Z _13700_/Z _13770_/Z _13840_/Z MUX.SEL0BUF\[0\]/X MUX.SEL1BUF\[0\]/X
+ vssd1 vssd1 vccd1 vccd1 Do[1] sky130_fd_sc_hd__mux4_1
XPHY_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13401_ _13401_/A _13404_/Y vssd1 vssd1 vccd1 vccd1 _13681_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10613_ _10635_/CLK line[45] vssd1 vssd1 vccd1 vccd1 _10614_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10883__A _13925_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11593_ _11615_/CLK line[109] vssd1 vssd1 vccd1 vccd1 _11594_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[2\].CG clk OVHB\[2\].CGAND/X vssd1 vssd1 vccd1 vccd1 OVHB\[2\].V/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_195_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09449__A _13920_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10544_ _10544_/A _10569_/Y vssd1 vssd1 vccd1 vccd1 _13624_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13332_ _13332_/CLK _13333_/X vssd1 vssd1 vccd1 vccd1 _13330_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_41_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[19\].VALID\[14\].FF OVHB\[19\].V/CLK A[21] vssd1 vssd1 vccd1 vccd1 OVHB\[19\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_10475_ _10495_/CLK line[110] vssd1 vssd1 vccd1 vccd1 _10476_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09168__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13263_ _13938_/X wr vssd1 vssd1 vccd1 vccd1 _13263_/X sky130_fd_sc_hd__and2_1
XFILLER_182_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12214_ _13934_/X vssd1 vssd1 vccd1 vccd1 _12214_/Y sky130_fd_sc_hd__inv_2
X_13194_ _13938_/X vssd1 vssd1 vccd1 vccd1 _13194_/Y sky130_fd_sc_hd__inv_2
XDATA\[9\].CLKBUF\[7\] clk vssd1 vssd1 vccd1 vccd1 _13892_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA_DATA\[22\].CLKBUF\[0\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12145_ _12175_/CLK line[96] vssd1 vssd1 vccd1 vccd1 _12146_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12025__D line[36] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07119__D line[97] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12076_ _12076_/A _12109_/Y vssd1 vssd1 vccd1 vccd1 _13756_/Z sky130_fd_sc_hd__ebufn_2
X_11027_ _11055_/CLK line[106] vssd1 vssd1 vccd1 vccd1 _11028_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06958__D line[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09334__D line[86] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_MUX.M\[1\].MUX\[2\]_A0 _13618_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12978_ _12980_/CLK line[88] vssd1 vssd1 vccd1 vccd1 _12979_/A sky130_fd_sc_hd__dfxtp_1
X_11929_ _11929_/A _11934_/Y vssd1 vssd1 vccd1 vccd1 _13889_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06693__D line[45] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05450_ _05450_/A _05459_/Y vssd1 vssd1 vccd1 vccd1 _13850_/Z sky130_fd_sc_hd__ebufn_2
X_05381_ _05385_/CLK line[71] vssd1 vssd1 vccd1 vccd1 _05382_/A sky130_fd_sc_hd__dfxtp_1
X_07120_ _07120_/A _07139_/Y vssd1 vssd1 vccd1 vccd1 _13840_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_173_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07051_ _07065_/CLK line[66] vssd1 vssd1 vccd1 vccd1 _07052_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_127_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09509__D line[38] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06002_ _06002_/A _06019_/Y vssd1 vssd1 vccd1 vccd1 _13842_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__04941__D line[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[21\].VALID\[6\].TOBUF OVHB\[21\].VALID\[6\].FF/Q OVHB\[21\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04923_/A2 sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[4\].VALID\[1\].FF_D A[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07953_ _07975_/CLK line[109] vssd1 vssd1 vccd1 vccd1 _07954_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11774__D line[49] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDATA\[8\].CLKBUF\[4\] clk vssd1 vssd1 vccd1 vccd1 _13507_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__06868__D line[125] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06904_ _06904_/A _06929_/Y vssd1 vssd1 vccd1 vccd1 _13624_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11129__A _13933_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07884_ _07884_/A _07909_/Y vssd1 vssd1 vccd1 vccd1 _13764_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09244__D line[59] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09623_ _13920_/Y wr vssd1 vssd1 vccd1 vccd1 _09623_/X sky130_fd_sc_hd__and2_1
X_06835_ _06855_/CLK line[110] vssd1 vssd1 vccd1 vccd1 _06836_/A sky130_fd_sc_hd__dfxtp_1
X_06766_ _06766_/A _06789_/Y vssd1 vssd1 vccd1 vccd1 _13766_/Z sky130_fd_sc_hd__ebufn_2
X_09554_ _13920_/Y vssd1 vssd1 vccd1 vccd1 _09554_/Y sky130_fd_sc_hd__inv_2
X_08505_ _08535_/CLK line[96] vssd1 vssd1 vccd1 vccd1 _08506_/A sky130_fd_sc_hd__dfxtp_1
X_05717_ _05735_/CLK line[111] vssd1 vssd1 vccd1 vccd1 _05718_/A sky130_fd_sc_hd__dfxtp_1
XPHY_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06697_ _06715_/CLK line[47] vssd1 vssd1 vccd1 vccd1 _06698_/A sky130_fd_sc_hd__dfxtp_1
X_09485_ _09515_/CLK line[32] vssd1 vssd1 vccd1 vccd1 _09486_/A sky130_fd_sc_hd__dfxtp_1
XPHY_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08436_ _08436_/A _08469_/Y vssd1 vssd1 vccd1 vccd1 _13756_/Z sky130_fd_sc_hd__ebufn_2
X_05648_ _05648_/A _05669_/Y vssd1 vssd1 vccd1 vccd1 _13768_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_12_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[1\].VALID\[12\].FF OVHB\[1\].V/CLK A[19] vssd1 vssd1 vccd1 vccd1 OVHB\[1\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_196_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08367_ _08395_/CLK line[42] vssd1 vssd1 vccd1 vccd1 _08368_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_168_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05579_ _05595_/CLK line[33] vssd1 vssd1 vccd1 vccd1 _05580_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XDECH.DEC0.AND2 A_h[3] A_h[4] vssd1 vssd1 vccd1 vccd1 _13960_/D sky130_fd_sc_hd__and2b_2
XANTENNA__11014__D line[86] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07318_ _07318_/A _07349_/Y vssd1 vssd1 vccd1 vccd1 _13758_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06108__D line[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08298_ _08298_/A _08329_/Y vssd1 vssd1 vccd1 vccd1 _13618_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_109_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11949__D line[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07249_ _07275_/CLK line[43] vssd1 vssd1 vccd1 vccd1 _07250_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_137_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09419__D line[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10260_ _10260_/A _10289_/Y vssd1 vssd1 vccd1 vccd1 _13620_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08323__D line[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10191_ _10215_/CLK line[108] vssd1 vssd1 vccd1 vccd1 _10192_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12423__A _13935_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XOVHB\[8\].VALID\[3\].FF OVHB\[8\].V/CLK A[10] vssd1 vssd1 vccd1 vccd1 OVHB\[8\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_13950_ A_h[0] vssd1 vssd1 vccd1 vccd1 _13960_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__05682__D line[95] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12901_ _12901_/A _12914_/Y vssd1 vssd1 vccd1 vccd1 _13741_/Z sky130_fd_sc_hd__ebufn_2
X_13881_ _13881_/A _13894_/Y vssd1 vssd1 vccd1 vccd1 _13881_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[17\].VALID\[12\].TOBUF OVHB\[17\].VALID\[12\].FF/Q OVHB\[17\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04929_/B2 sky130_fd_sc_hd__ebufn_2
X_12832_ _12840_/CLK line[21] vssd1 vssd1 vccd1 vccd1 _12833_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_46_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XDATA\[7\].CLKBUF\[1\] clk vssd1 vssd1 vccd1 vccd1 _13122_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_61_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12763_ _12763_/A _12774_/Y vssd1 vssd1 vccd1 vccd1 _13883_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11714_ _11720_/CLK line[22] vssd1 vssd1 vccd1 vccd1 _11715_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12694_ _12700_/CLK line[86] vssd1 vssd1 vccd1 vccd1 _12695_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11645_ _11645_/A _11654_/Y vssd1 vssd1 vccd1 vccd1 _13885_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11576_ _11580_/CLK line[87] vssd1 vssd1 vccd1 vccd1 _11577_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08083__A _13932_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[25\].VALID\[10\].FF OVHB\[25\].V/CLK A[17] vssd1 vssd1 vccd1 vccd1 OVHB\[25\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10763__D line[99] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13315_ _13315_/A _13334_/Y vssd1 vssd1 vccd1 vccd1 _13875_/Z sky130_fd_sc_hd__ebufn_2
X_10527_ _10527_/A _10534_/Y vssd1 vssd1 vccd1 vccd1 _13887_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_183_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05857__D line[47] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08233__D line[109] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10458_ _10460_/CLK line[88] vssd1 vssd1 vccd1 vccd1 _10459_/A sky130_fd_sc_hd__dfxtp_1
X_13246_ _13260_/CLK line[82] vssd1 vssd1 vccd1 vccd1 _13247_/A sky130_fd_sc_hd__dfxtp_1
X_10389_ _10389_/A _10394_/Y vssd1 vssd1 vccd1 vccd1 _13749_/Z sky130_fd_sc_hd__ebufn_2
X_13177_ _13177_/A _13194_/Y vssd1 vssd1 vccd1 vccd1 _13737_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[10\].VALID\[11\].TOBUF OVHB\[10\].VALID\[11\].FF/Q OVHB\[10\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04915_/B2 sky130_fd_sc_hd__ebufn_2
X_12128_ _12140_/CLK line[83] vssd1 vssd1 vccd1 vccd1 _12129_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_96_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XDATA\[27\].CLKBUF\[5\] clk vssd1 vssd1 vccd1 vccd1 _10462_/CLK sky130_fd_sc_hd__clkbuf_4
XMUX.M\[3\].MUX\[6\] _13661_/Z _13731_/Z _13801_/Z _13871_/Z MUX.SEL0BUF\[3\]/X MUX.SEL1BUF\[3\]/X
+ vssd1 vssd1 vccd1 vccd1 Do[30] sky130_fd_sc_hd__mux4_1
X_04950_ _04950_/A _04969_/Y vssd1 vssd1 vccd1 vccd1 _13630_/Z sky130_fd_sc_hd__ebufn_2
X_12059_ _12059_/A _12074_/Y vssd1 vssd1 vccd1 vccd1 _13739_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_84_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_DATA\[20\].CLKBUF\[2\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09999__D line[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06620_ _06620_/A _06649_/Y vssd1 vssd1 vccd1 vccd1 _13620_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10003__D line[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08258__A _13932_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06551_ _06575_/CLK line[108] vssd1 vssd1 vccd1 vccd1 _06552_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10938__D line[51] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[6\].VALID\[5\].FF OVHB\[6\].V/CLK A[12] vssd1 vssd1 vccd1 vccd1 OVHB\[6\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XOVHB\[15\].VALID\[12\].FF OVHB\[15\].V/CLK A[19] vssd1 vssd1 vccd1 vccd1 OVHB\[15\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13314__D line[113] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05502_ _05502_/A _05529_/Y vssd1 vssd1 vccd1 vccd1 _13622_/Z sky130_fd_sc_hd__ebufn_2
X_09270_ _09270_/CLK line[57] vssd1 vssd1 vccd1 vccd1 _09271_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08408__D line[61] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06482_ _06482_/A _06509_/Y vssd1 vssd1 vccd1 vccd1 _13762_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_61_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08221_ _08221_/A _08224_/Y vssd1 vssd1 vccd1 vccd1 _13821_/Z sky130_fd_sc_hd__ebufn_2
X_05433_ _05455_/CLK line[109] vssd1 vssd1 vccd1 vccd1 _05434_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_20_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08152_ _08152_/CLK _08153_/X vssd1 vssd1 vccd1 vccd1 _08150_/CLK sky130_fd_sc_hd__dlclkp_1
X_05364_ _05364_/A _05389_/Y vssd1 vssd1 vccd1 vccd1 _13764_/Z sky130_fd_sc_hd__ebufn_2
X_07103_ _13909_/Y wr vssd1 vssd1 vccd1 vccd1 _07103_/X sky130_fd_sc_hd__and2_1
X_08083_ _13932_/X wr vssd1 vssd1 vccd1 vccd1 _08083_/X sky130_fd_sc_hd__and2_1
X_05295_ _05315_/CLK line[46] vssd1 vssd1 vccd1 vccd1 _05296_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_134_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07034_ _13909_/Y vssd1 vssd1 vccd1 vccd1 _07034_/Y sky130_fd_sc_hd__inv_2
XANTENNA__07982__D line[122] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08985_ _08985_/A _08994_/Y vssd1 vssd1 vccd1 vccd1 _13745_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_196_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06598__D line[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07936_ _07940_/CLK line[87] vssd1 vssd1 vccd1 vccd1 _07937_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_29_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07867_ _07867_/A _07874_/Y vssd1 vssd1 vccd1 vccd1 _13747_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_83_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09606_ _09620_/CLK line[82] vssd1 vssd1 vccd1 vccd1 _09607_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[26\].CLKBUF\[2\] clk vssd1 vssd1 vccd1 vccd1 _10077_/CLK sky130_fd_sc_hd__clkbuf_4
X_06818_ _06820_/CLK line[88] vssd1 vssd1 vccd1 vccd1 _06819_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_73_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07798_ _07800_/CLK line[24] vssd1 vssd1 vccd1 vccd1 _07799_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05007__D line[42] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09537_ _09537_/A _09554_/Y vssd1 vssd1 vccd1 vccd1 _13737_/Z sky130_fd_sc_hd__ebufn_2
X_06749_ _06749_/A _06754_/Y vssd1 vssd1 vccd1 vccd1 _13749_/Z sky130_fd_sc_hd__ebufn_2
XPHY_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09468_ _09480_/CLK line[19] vssd1 vssd1 vccd1 vccd1 _09469_/A sky130_fd_sc_hd__dfxtp_1
XPHY_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07222__D line[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08419_ _08419_/A _08434_/Y vssd1 vssd1 vccd1 vccd1 _13739_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09399_ _09399_/A _09414_/Y vssd1 vssd1 vccd1 vccd1 _13879_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XOVHB\[30\].VALID\[11\].TOBUF OVHB\[30\].VALID\[11\].FF/Q OVHB\[30\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04915_/B2 sky130_fd_sc_hd__ebufn_2
X_11430_ _11440_/CLK line[20] vssd1 vssd1 vccd1 vccd1 _11431_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11679__D line[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XOVHB\[4\].VALID\[7\].FF OVHB\[4\].V/CLK A[14] vssd1 vssd1 vccd1 vccd1 OVHB\[4\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_11361_ _11361_/A _11374_/Y vssd1 vssd1 vccd1 vccd1 _13881_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_125_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_MUX.M\[3\].MUX\[3\]_A2 _13795_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09149__D line[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13100_ _13120_/CLK line[30] vssd1 vssd1 vccd1 vccd1 _13101_/A sky130_fd_sc_hd__dfxtp_1
X_10312_ _10320_/CLK line[21] vssd1 vssd1 vccd1 vccd1 _10313_/A sky130_fd_sc_hd__dfxtp_1
X_11292_ _11300_/CLK line[85] vssd1 vssd1 vccd1 vccd1 _11293_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_180_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10243_ _10243_/A _10254_/Y vssd1 vssd1 vccd1 vccd1 _13883_/Z sky130_fd_sc_hd__ebufn_2
X_13031_ _13031_/A _13054_/Y vssd1 vssd1 vccd1 vccd1 _13871_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[3\].VALID\[3\].TOBUF OVHB\[3\].VALID\[3\].FF/Q OVHB\[3\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04919_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__08988__D line[56] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10174_ _10180_/CLK line[86] vssd1 vssd1 vccd1 vccd1 _10175_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[1\].VALID\[14\].FF_D A[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[28\].VALID\[6\].TOBUF OVHB\[28\].VALID\[6\].FF/Q OVHB\[28\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04923_/A2 sky130_fd_sc_hd__ebufn_2
XFILLER_154_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12303__D line[35] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[19\].CLKBUF\[3\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13933_ _13938_/C _13938_/A _13938_/B _13938_/D vssd1 vssd1 vccd1 vccd1 _13933_/X
+ sky130_fd_sc_hd__and4bb_4
XOVHB\[28\].VOBUF OVHB\[28\].V/Q OVHB\[28\].INV/Y vssd1 vssd1 vccd1 vccd1 _04912_/B1
+ sky130_fd_sc_hd__ebufn_2
XFILLER_47_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13864_ _13890_/CLK line[123] vssd1 vssd1 vccd1 vccd1 _13865_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09612__D line[85] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12815_ _12815_/A _12844_/Y vssd1 vssd1 vccd1 vccd1 _13655_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_34_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13795_ _13795_/A _13824_/Y vssd1 vssd1 vccd1 vccd1 _13795_/Z sky130_fd_sc_hd__ebufn_2
X_12746_ _12770_/CLK line[124] vssd1 vssd1 vccd1 vccd1 _12747_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_203_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12677_ _12677_/A _12704_/Y vssd1 vssd1 vccd1 vccd1 _13797_/Z sky130_fd_sc_hd__ebufn_2
XPHY_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06971__D line[44] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XDATA\[15\].CLKBUF\[5\] clk vssd1 vssd1 vccd1 vccd1 _06822_/CLK sky130_fd_sc_hd__clkbuf_4
X_11628_ _11650_/CLK line[125] vssd1 vssd1 vccd1 vccd1 _11629_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_8_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11589__D line[107] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10493__D line[104] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11559_ _11559_/A _11584_/Y vssd1 vssd1 vccd1 vccd1 _13799_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05587__D line[37] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[0\].VALID\[4\].FF_D A[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05080_ _05080_/A _05109_/Y vssd1 vssd1 vccd1 vccd1 _13760_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13159__A _13938_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08898__D line[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13229_ _13938_/X vssd1 vssd1 vccd1 vccd1 _13229_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XOVHB\[2\].VALID\[9\].FF OVHB\[2\].V/CLK A[16] vssd1 vssd1 vccd1 vccd1 OVHB\[2\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_08770_ _08780_/CLK line[84] vssd1 vssd1 vccd1 vccd1 _08771_/A sky130_fd_sc_hd__dfxtp_1
X_05982_ _05982_/CLK _05983_/X vssd1 vssd1 vccd1 vccd1 _05980_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_97_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_04933_ _04933_/A _04933_/B _04933_/C _04933_/D vssd1 vssd1 vccd1 vccd1 _04934_/D
+ sky130_fd_sc_hd__or4_2
XANTENNA__06211__D line[66] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07721_ _07721_/A _07734_/Y vssd1 vssd1 vccd1 vccd1 _13881_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_65_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07652_ _07660_/CLK line[85] vssd1 vssd1 vccd1 vccd1 _07653_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_80_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09522__D line[58] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06603_ _06603_/A _06614_/Y vssd1 vssd1 vccd1 vccd1 _13883_/Z sky130_fd_sc_hd__ebufn_2
X_07583_ _07583_/A _07594_/Y vssd1 vssd1 vccd1 vccd1 _13743_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10668__D line[56] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13044__D line[118] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09322_ _09340_/CLK line[95] vssd1 vssd1 vccd1 vccd1 _09323_/A sky130_fd_sc_hd__dfxtp_1
X_06534_ _06540_/CLK line[86] vssd1 vssd1 vccd1 vccd1 _06535_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08138__D line[51] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06465_ _06465_/A _06474_/Y vssd1 vssd1 vccd1 vccd1 _13745_/Z sky130_fd_sc_hd__ebufn_2
X_09253_ _09253_/A _09274_/Y vssd1 vssd1 vccd1 vccd1 _13733_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_194_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_OVHB\[3\].VALID\[10\].FF_D A[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05416_ _05420_/CLK line[87] vssd1 vssd1 vccd1 vccd1 _05417_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_166_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08204_ _08220_/CLK line[81] vssd1 vssd1 vccd1 vccd1 _08205_/A sky130_fd_sc_hd__dfxtp_1
X_09184_ _09200_/CLK line[17] vssd1 vssd1 vccd1 vccd1 _09185_/A sky130_fd_sc_hd__dfxtp_1
X_06396_ _06400_/CLK line[23] vssd1 vssd1 vccd1 vccd1 _06397_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_194_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08135_ _08135_/A _08154_/Y vssd1 vssd1 vccd1 vccd1 _13735_/Z sky130_fd_sc_hd__ebufn_2
X_05347_ _05347_/A _05354_/Y vssd1 vssd1 vccd1 vccd1 _13747_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_107_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05497__D line[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08066_ _08080_/CLK line[18] vssd1 vssd1 vccd1 vccd1 _08067_/A sky130_fd_sc_hd__dfxtp_1
X_05278_ _05280_/CLK line[24] vssd1 vssd1 vccd1 vccd1 _05279_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[14\].CLKBUF\[2\] clk vssd1 vssd1 vccd1 vccd1 _06437_/CLK sky130_fd_sc_hd__clkbuf_4
X_07017_ _07017_/A _07034_/Y vssd1 vssd1 vccd1 vccd1 _13737_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[30\].VALID\[3\].FF OVHB\[30\].V/CLK A[10] vssd1 vssd1 vccd1 vccd1 OVHB\[30\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_1_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08601__D line[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13219__D line[70] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[11\].VALID\[10\].FF OVHB\[11\].V/CLK A[17] vssd1 vssd1 vccd1 vccd1 OVHB\[11\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_08968_ _08990_/CLK line[61] vssd1 vssd1 vccd1 vccd1 _08969_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_103_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[15\].VALID\[1\].FF_D A[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07919_ _07919_/A _07944_/Y vssd1 vssd1 vccd1 vccd1 _13799_/Z sky130_fd_sc_hd__ebufn_2
X_08899_ _08899_/A _08924_/Y vssd1 vssd1 vccd1 vccd1 _13659_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_84_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10930_ _10950_/CLK line[62] vssd1 vssd1 vccd1 vccd1 _10931_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[23\].CGAND_B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05960__D line[94] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10578__D line[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10861_ _10861_/A _10884_/Y vssd1 vssd1 vccd1 vccd1 _13661_/Z sky130_fd_sc_hd__ebufn_2
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12600_ _12630_/CLK line[48] vssd1 vssd1 vccd1 vccd1 _12601_/A sky130_fd_sc_hd__dfxtp_1
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_OVHB\[8\].CGAND_B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[27\].CGAND_A _13923_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13580_ _13610_/CLK line[112] vssd1 vssd1 vccd1 vccd1 _13581_/A sky130_fd_sc_hd__dfxtp_1
X_10792_ _10810_/CLK line[127] vssd1 vssd1 vccd1 vccd1 _10793_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_25_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XOVHB\[1\].VALID\[8\].TOBUF OVHB\[1\].VALID\[8\].FF/Q OVHB\[1\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04931_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[25\].CG_CLK clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12531_ _12531_/A _12564_/Y vssd1 vssd1 vccd1 vccd1 _13651_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12793__D line[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07887__D line[79] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12462_ _12490_/CLK line[122] vssd1 vssd1 vccd1 vccd1 _12463_/A sky130_fd_sc_hd__dfxtp_1
X_11413_ _11413_/A _11444_/Y vssd1 vssd1 vccd1 vccd1 _13653_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11202__D line[58] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12393_ _12393_/A _12424_/Y vssd1 vssd1 vccd1 vccd1 _13793_/Z sky130_fd_sc_hd__ebufn_2
X_11344_ _11370_/CLK line[123] vssd1 vssd1 vccd1 vccd1 _11345_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[29\].VALID\[4\].FF OVHB\[29\].V/CLK A[11] vssd1 vssd1 vccd1 vccd1 OVHB\[29\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__05200__D line[116] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11275_ _11275_/A _11304_/Y vssd1 vssd1 vccd1 vccd1 _13795_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.M\[2\].MUX\[4\]_A0 _13671_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13014_ _13014_/A _13019_/Y vssd1 vssd1 vccd1 vccd1 _13854_/Z sky130_fd_sc_hd__ebufn_2
X_10226_ _10250_/CLK line[124] vssd1 vssd1 vccd1 vccd1 _10227_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08511__D line[108] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[6\].VALID\[8\].FF_D A[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13129__D line[43] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12033__D line[40] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10157_ _10157_/A _10184_/Y vssd1 vssd1 vccd1 vccd1 _13797_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_79_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[11\].VALID\[1\].FF OVHB\[11\].V/CLK A[8] vssd1 vssd1 vccd1 vccd1 OVHB\[11\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07127__D line[101] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10088_ _10110_/CLK line[61] vssd1 vssd1 vccd1 vccd1 _10089_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12968__D line[83] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13916_ _13916_/A _13916_/B _13916_/C _13916_/D vssd1 vssd1 vccd1 vccd1 _13916_/X
+ sky130_fd_sc_hd__and4_4
XFILLER_75_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13847_ _13855_/CLK line[101] vssd1 vssd1 vccd1 vccd1 _13848_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[17\].CLKBUF\[5\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13778_ _13778_/A _13789_/Y vssd1 vssd1 vccd1 vccd1 _13778_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_31_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MUX.M\[0\].MUX\[0\]_A1 _13686_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12729_ _12735_/CLK line[102] vssd1 vssd1 vccd1 vccd1 _12730_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06250_ _06260_/CLK line[84] vssd1 vssd1 vccd1 vccd1 _06251_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_176_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05201_ _05201_/A _05214_/Y vssd1 vssd1 vccd1 vccd1 _13881_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_209_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12208__D line[120] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06181_ _06181_/A _06194_/Y vssd1 vssd1 vccd1 vccd1 _13741_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_144_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05132_ _05140_/CLK line[85] vssd1 vssd1 vccd1 vccd1 _05133_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_143_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05110__D line[80] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09940_ _09970_/CLK line[112] vssd1 vssd1 vccd1 vccd1 _09941_/A sky130_fd_sc_hd__dfxtp_1
X_05063_ _05063_/A _05074_/Y vssd1 vssd1 vccd1 vccd1 _13743_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_132_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09871_ _09871_/A _09904_/Y vssd1 vssd1 vccd1 vccd1 _13791_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_124_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_OVHB\[28\].VALID\[1\].FF_D A[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08822_ _08850_/CLK line[122] vssd1 vssd1 vccd1 vccd1 _08823_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07037__D line[74] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[27\].VALID\[6\].FF OVHB\[27\].V/CLK A[13] vssd1 vssd1 vccd1 vccd1 OVHB\[27\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_57_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08753_ _08753_/A _08784_/Y vssd1 vssd1 vccd1 vccd1 _13793_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[8\].VALID\[14\].FF_D A[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[7\].VALID\[14\].TOBUF OVHB\[7\].VALID\[14\].FF/Q OVHB\[7\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/B2 sky130_fd_sc_hd__ebufn_2
X_05965_ _05965_/A _05984_/Y vssd1 vssd1 vccd1 vccd1 _13805_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11782__D line[53] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07704_ _07730_/CLK line[123] vssd1 vssd1 vccd1 vccd1 _07705_/A sky130_fd_sc_hd__dfxtp_1
X_04916_ A_h[18] _04916_/B2 A_h[18] _04916_/B2 vssd1 vssd1 vccd1 vccd1 _04917_/D sky130_fd_sc_hd__a2bb2oi_2
XANTENNA__06876__D line[114] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[6\].VALID\[12\].FF OVHB\[6\].V/CLK A[19] vssd1 vssd1 vccd1 vccd1 OVHB\[6\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_08684_ _08710_/CLK line[59] vssd1 vssd1 vccd1 vccd1 _08685_/A sky130_fd_sc_hd__dfxtp_1
X_05896_ _05910_/CLK line[50] vssd1 vssd1 vccd1 vccd1 _05897_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09252__D line[63] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07635_ _07635_/A _07664_/Y vssd1 vssd1 vccd1 vccd1 _13795_/Z sky130_fd_sc_hd__ebufn_2
X_07566_ _07590_/CLK line[60] vssd1 vssd1 vccd1 vccd1 _07567_/A sky130_fd_sc_hd__dfxtp_1
X_09305_ _09305_/CLK line[73] vssd1 vssd1 vccd1 vccd1 _09306_/A sky130_fd_sc_hd__dfxtp_1
X_06517_ _06517_/A _06544_/Y vssd1 vssd1 vccd1 vccd1 _13797_/Z sky130_fd_sc_hd__ebufn_2
X_07497_ _07497_/A _07524_/Y vssd1 vssd1 vccd1 vccd1 _13657_/Z sky130_fd_sc_hd__ebufn_2
X_09236_ _09236_/A _09239_/Y vssd1 vssd1 vccd1 vccd1 _13716_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_186_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06448_ _06470_/CLK line[61] vssd1 vssd1 vccd1 vccd1 _06449_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07500__D line[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12118__D line[93] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06379_ _06379_/A _06404_/Y vssd1 vssd1 vccd1 vccd1 _13659_/Z sky130_fd_sc_hd__ebufn_2
X_09167_ _09167_/CLK _09168_/X vssd1 vssd1 vccd1 vccd1 _09165_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__06116__D line[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08118_ _13932_/X wr vssd1 vssd1 vccd1 vccd1 _08118_/X sky130_fd_sc_hd__and2_1
XFILLER_174_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09098_ _13915_/X wr vssd1 vssd1 vccd1 vccd1 _09098_/X sky130_fd_sc_hd__and2_1
XOVHB\[27\].VALID\[10\].TOBUF OVHB\[27\].VALID\[10\].FF/Q OVHB\[27\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04932_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__11957__D line[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[0\].VALID\[13\].TOBUF OVHB\[0\].VALID\[13\].FF/Q OVHB\[0\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04916_/B2 sky130_fd_sc_hd__ebufn_2
X_08049_ _13932_/X vssd1 vssd1 vccd1 vccd1 _08049_/Y sky130_fd_sc_hd__inv_2
XFILLER_107_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09427__D line[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11060_ _11090_/CLK line[112] vssd1 vssd1 vccd1 vccd1 _11061_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10011_ _10011_/A _10044_/Y vssd1 vssd1 vccd1 vccd1 _13651_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_192_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11692__D line[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11962_ _11962_/A _11969_/Y vssd1 vssd1 vccd1 vccd1 _13642_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_151_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05690__D line[84] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13701_ _13715_/CLK line[34] vssd1 vssd1 vccd1 vccd1 _13702_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[11\].V_RESET_B rst_n vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10913_ _10915_/CLK line[40] vssd1 vssd1 vccd1 vccd1 _10914_/A sky130_fd_sc_hd__dfxtp_1
X_11893_ _11895_/CLK line[104] vssd1 vssd1 vccd1 vccd1 _11894_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_17_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13632_ _13632_/A _13649_/Y vssd1 vssd1 vccd1 vccd1 _13632_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[25\].VALID\[8\].FF OVHB\[25\].V/CLK A[15] vssd1 vssd1 vccd1 vccd1 OVHB\[25\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_10844_ _10844_/A _10849_/Y vssd1 vssd1 vccd1 vccd1 _13644_/Z sky130_fd_sc_hd__ebufn_2
X_13563_ _13575_/CLK line[99] vssd1 vssd1 vccd1 vccd1 _13564_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_158_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10775_ _10775_/CLK line[105] vssd1 vssd1 vccd1 vccd1 _10776_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_12_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12514_ _12514_/A _12529_/Y vssd1 vssd1 vccd1 vccd1 _13634_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_13_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13494_ _13494_/A _13509_/Y vssd1 vssd1 vccd1 vccd1 _13774_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_8_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12445_ _12455_/CLK line[100] vssd1 vssd1 vccd1 vccd1 _12446_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_138_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06026__D line[124] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12376_ _12376_/A _12389_/Y vssd1 vssd1 vccd1 vccd1 _13776_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_126_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11867__D line[106] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10771__D line[103] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11327_ _11335_/CLK line[101] vssd1 vssd1 vccd1 vccd1 _11328_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05865__D line[36] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08241__D line[98] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11258_ _11258_/A _11269_/Y vssd1 vssd1 vccd1 vccd1 _13778_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_192_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10209_ _10215_/CLK line[102] vssd1 vssd1 vccd1 vccd1 _10210_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_67_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11189_ _11195_/CLK line[38] vssd1 vssd1 vccd1 vccd1 _11190_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_39_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__04927__B1 A_h[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12698__D line[88] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05750_ _05770_/CLK line[126] vssd1 vssd1 vccd1 vccd1 _05751_/A sky130_fd_sc_hd__dfxtp_1
X_05681_ _05681_/A _05704_/Y vssd1 vssd1 vccd1 vccd1 _13801_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_35_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11107__D line[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07420_ _07450_/CLK line[112] vssd1 vssd1 vccd1 vccd1 _07421_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_211_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05105__D line[73] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09800__D line[48] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10946__D line[55] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07351_ _07351_/A _07384_/Y vssd1 vssd1 vccd1 vccd1 _13791_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_210_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13322__D line[117] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06302_ _06330_/CLK line[122] vssd1 vssd1 vccd1 vccd1 _06303_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08416__D line[50] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07282_ _07310_/CLK line[58] vssd1 vssd1 vccd1 vccd1 _07283_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[8\].VALID\[8\].TOBUF OVHB\[8\].VALID\[8\].FF/Q OVHB\[8\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04931_/B2 sky130_fd_sc_hd__ebufn_2
X_09021_ _09025_/CLK line[71] vssd1 vssd1 vccd1 vccd1 _09022_/A sky130_fd_sc_hd__dfxtp_1
X_06233_ _06233_/A _06264_/Y vssd1 vssd1 vccd1 vccd1 _13793_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_191_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_DATA\[15\].CLKBUF\[7\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08713__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06164_ _06190_/CLK line[59] vssd1 vssd1 vccd1 vccd1 _06165_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.SEL1BUF\[1\]_A A[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05115_ _05115_/A _05144_/Y vssd1 vssd1 vccd1 vccd1 _13795_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_105_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10681__D line[76] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06095_ _06095_/A _06124_/Y vssd1 vssd1 vccd1 vccd1 _13655_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05775__D line[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05046_ _05070_/CLK line[60] vssd1 vssd1 vccd1 vccd1 _05047_/A sky130_fd_sc_hd__dfxtp_1
X_09923_ _09935_/CLK line[99] vssd1 vssd1 vccd1 vccd1 _09924_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[11\].VALID\[4\].FF_D A[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09041__TE_B _09064_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09854_ _09854_/A _09869_/Y vssd1 vssd1 vccd1 vccd1 _13774_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__04969__A _13931_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07990__D line[126] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08805_ _08815_/CLK line[100] vssd1 vssd1 vccd1 vccd1 _08806_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_100_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09785_ _09795_/CLK line[36] vssd1 vssd1 vccd1 vccd1 _09786_/A sky130_fd_sc_hd__dfxtp_1
X_06997_ _06997_/CLK _06998_/X vssd1 vssd1 vccd1 vccd1 _06995_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_65_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08736_ _08736_/A _08749_/Y vssd1 vssd1 vccd1 vccd1 _13776_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_26_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05948_ _13902_/X wr vssd1 vssd1 vccd1 vccd1 _05948_/X sky130_fd_sc_hd__and2_1
XANTENNA_DATA\[8\].CLKBUF\[7\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08667_ _08675_/CLK line[37] vssd1 vssd1 vccd1 vccd1 _08668_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05879_ _13902_/X vssd1 vssd1 vccd1 vccd1 _05879_/Y sky130_fd_sc_hd__inv_2
XPHY_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07618_ _07618_/A _07629_/Y vssd1 vssd1 vccd1 vccd1 _13778_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_81_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08598_ _08598_/A _08609_/Y vssd1 vssd1 vccd1 vccd1 _13638_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05015__D line[46] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10856__D line[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07549_ _07555_/CLK line[38] vssd1 vssd1 vccd1 vccd1 _07550_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13232__D line[90] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10560_ _10560_/A _10569_/Y vssd1 vssd1 vccd1 vccd1 _13640_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_22_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07230__D line[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[30\].CLKBUF\[0\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09219_ _09235_/CLK line[33] vssd1 vssd1 vccd1 vccd1 _09220_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_10_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10491_ _10495_/CLK line[103] vssd1 vssd1 vccd1 vccd1 _10492_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[5\].CLKBUF\[6\] clk vssd1 vssd1 vccd1 vccd1 _12737_/CLK sky130_fd_sc_hd__clkbuf_4
X_12230_ _12230_/A _12249_/Y vssd1 vssd1 vccd1 vccd1 _13630_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_30_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12161_ _12175_/CLK line[98] vssd1 vssd1 vccd1 vccd1 _12162_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_123_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_OVHB\[10\].VALID\[12\].FF_D A[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09157__D line[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11112_ _11112_/A _11129_/Y vssd1 vssd1 vccd1 vccd1 _13632_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_1_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[2\].VALID\[10\].FF OVHB\[2\].V/CLK A[17] vssd1 vssd1 vccd1 vccd1 OVHB\[2\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_12092_ _12092_/A _12109_/Y vssd1 vssd1 vccd1 vccd1 _13772_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[15\].VALID\[3\].TOBUF OVHB\[15\].VALID\[3\].FF/Q OVHB\[15\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04919_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.M\[2\].MUX\[1\]_A3 _13875_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11043_ _11055_/CLK line[99] vssd1 vssd1 vccd1 vccd1 _11044_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_39_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13407__D line[42] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12311__D line[39] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12994_ _12994_/A _13019_/Y vssd1 vssd1 vccd1 vccd1 _13834_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07405__D line[100] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DEC.DEC0.AND1_B A[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11945_ _11965_/CLK line[14] vssd1 vssd1 vccd1 vccd1 _11946_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_189_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[20\].VALID\[11\].FF_D A[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11876_ _11876_/A _11899_/Y vssd1 vssd1 vccd1 vccd1 _13836_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09620__D line[89] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13615_ _13645_/CLK line[0] vssd1 vssd1 vccd1 vccd1 _13616_/A sky130_fd_sc_hd__dfxtp_1
X_10827_ _10845_/CLK line[15] vssd1 vssd1 vccd1 vccd1 _10828_/A sky130_fd_sc_hd__dfxtp_1
X_13546_ _13546_/A _13579_/Y vssd1 vssd1 vccd1 vccd1 _13826_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_13_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10758_ _10758_/A _10779_/Y vssd1 vssd1 vccd1 vccd1 _13838_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[31\].VALID\[0\].FF_D A[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07140__D line[112] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13477_ _13505_/CLK line[74] vssd1 vssd1 vccd1 vccd1 _13478_/A sky130_fd_sc_hd__dfxtp_1
X_10689_ _10705_/CLK line[65] vssd1 vssd1 vccd1 vccd1 _10690_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_145_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12428_ _12428_/A _12459_/Y vssd1 vssd1 vccd1 vccd1 _13828_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06334__A _13903_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11597__D line[111] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[30\].VALID\[10\].FF_D A[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12359_ _12385_/CLK line[75] vssd1 vssd1 vccd1 vccd1 _12360_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05595__D line[41] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06053__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_OVHB\[24\].VALID\[4\].FF_D A[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09067__D line[106] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDATA\[4\].CLKBUF\[3\] clk vssd1 vssd1 vccd1 vccd1 _12352_/CLK sky130_fd_sc_hd__clkbuf_4
X_06920_ _06920_/A _06929_/Y vssd1 vssd1 vccd1 vccd1 _13640_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_68_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06851_ _06855_/CLK line[103] vssd1 vssd1 vccd1 vccd1 _06852_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12221__D line[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05802_ _05802_/A _05809_/Y vssd1 vssd1 vccd1 vccd1 _13642_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[17\].VALID\[8\].FF_D A[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__04939__D line[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09570_ _09570_/A _09589_/Y vssd1 vssd1 vccd1 vccd1 _13770_/Z sky130_fd_sc_hd__ebufn_2
X_06782_ _06782_/A _06789_/Y vssd1 vssd1 vccd1 vccd1 _13782_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07315__D line[64] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08521_ _08535_/CLK line[98] vssd1 vssd1 vccd1 vccd1 _08522_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_82_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05733_ _05735_/CLK line[104] vssd1 vssd1 vccd1 vccd1 _05734_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_36_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[21\].VALID\[2\].TOBUF OVHB\[21\].VALID\[2\].FF/Q OVHB\[21\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04930_/B2 sky130_fd_sc_hd__ebufn_2
X_08452_ _08452_/A _08469_/Y vssd1 vssd1 vccd1 vccd1 _13772_/Z sky130_fd_sc_hd__ebufn_2
X_05664_ _05664_/A _05669_/Y vssd1 vssd1 vccd1 vccd1 _13784_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06509__A _13904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09530__D line[62] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07403_ _07415_/CLK line[99] vssd1 vssd1 vccd1 vccd1 _07404_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_50_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05595_ _05595_/CLK line[41] vssd1 vssd1 vccd1 vccd1 _05596_/A sky130_fd_sc_hd__dfxtp_1
X_08383_ _08395_/CLK line[35] vssd1 vssd1 vccd1 vccd1 _08384_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06228__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[29\].CLKBUF\[1\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07334_ _07334_/A _07349_/Y vssd1 vssd1 vccd1 vccd1 _13774_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08146__D line[55] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[14\].V_D TIE/HI vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07265_ _07275_/CLK line[36] vssd1 vssd1 vccd1 vccd1 _07266_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[24\].CLKBUF\[7\] clk vssd1 vssd1 vccd1 vccd1 _09692_/CLK sky130_fd_sc_hd__clkbuf_4
X_09004_ _09004_/A _09029_/Y vssd1 vssd1 vccd1 vccd1 _13764_/Z sky130_fd_sc_hd__ebufn_2
X_06216_ _06216_/A _06229_/Y vssd1 vssd1 vccd1 vccd1 _13776_/Z sky130_fd_sc_hd__ebufn_2
X_07196_ _07196_/A _07209_/Y vssd1 vssd1 vccd1 vccd1 _13636_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_3_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_OVHB\[29\].V_D TIE/HI vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XOVHB\[16\].VALID\[10\].FF OVHB\[16\].V/CLK A[17] vssd1 vssd1 vccd1 vccd1 OVHB\[16\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_06147_ _06155_/CLK line[37] vssd1 vssd1 vccd1 vccd1 _06148_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_145_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11300__D line[89] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06078_ _06078_/A _06089_/Y vssd1 vssd1 vccd1 vccd1 _13638_/Z sky130_fd_sc_hd__ebufn_2
X_05029_ _05035_/CLK line[38] vssd1 vssd1 vccd1 vccd1 _05030_/A sky130_fd_sc_hd__dfxtp_1
X_09906_ _09906_/A _09939_/Y vssd1 vssd1 vccd1 vccd1 _13826_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09705__D line[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09837_ _09865_/CLK line[74] vssd1 vssd1 vccd1 vccd1 _09838_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[3\].CLKBUF\[0\] clk vssd1 vssd1 vccd1 vccd1 _11967_/CLK sky130_fd_sc_hd__clkbuf_4
X_09768_ _09768_/A _09799_/Y vssd1 vssd1 vccd1 vccd1 _13688_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_92_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07803__A _13912_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08719_ _08745_/CLK line[75] vssd1 vssd1 vccd1 vccd1 _08720_/A sky130_fd_sc_hd__dfxtp_1
X_09699_ _09725_/CLK line[11] vssd1 vssd1 vccd1 vccd1 _09700_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11970__D line[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11730_ _11730_/A _11759_/Y vssd1 vssd1 vccd1 vccd1 _13690_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10586__D line[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11661_ _11685_/CLK line[12] vssd1 vssd1 vccd1 vccd1 _11662_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13400_ _13400_/CLK line[25] vssd1 vssd1 vccd1 vccd1 _13401_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[13\].VALID\[8\].TOBUF OVHB\[13\].VALID\[8\].FF/Q OVHB\[13\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04931_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__08056__D line[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10612_ _10612_/A _10639_/Y vssd1 vssd1 vccd1 vccd1 _13692_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11592_ _11592_/A _11619_/Y vssd1 vssd1 vccd1 vccd1 _13832_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10883__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MUX.M\[3\].MUX\[6\]_A0 _13661_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13331_ _13331_/A _13334_/Y vssd1 vssd1 vccd1 vccd1 _13891_/Z sky130_fd_sc_hd__ebufn_2
X_10543_ _10565_/CLK line[13] vssd1 vssd1 vccd1 vccd1 _10544_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07895__D line[68] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_DATA\[2\].CLKBUF\[0\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13262_ _13262_/CLK _13263_/X vssd1 vssd1 vccd1 vccd1 _13260_/CLK sky130_fd_sc_hd__dlclkp_1
X_10474_ _10474_/A _10499_/Y vssd1 vssd1 vccd1 vccd1 _13834_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_155_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12213_ _13934_/X wr vssd1 vssd1 vccd1 vccd1 _12213_/X sky130_fd_sc_hd__and2_1
XFILLER_6_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13193_ _13938_/X wr vssd1 vssd1 vccd1 vccd1 _13193_/X sky130_fd_sc_hd__and2_1
XFILLER_123_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11210__D line[62] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12144_ _13934_/X vssd1 vssd1 vccd1 vccd1 _12144_/Y sky130_fd_sc_hd__inv_2
XDATA\[23\].CLKBUF\[4\] clk vssd1 vssd1 vccd1 vccd1 _09307_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__06304__D line[123] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12075_ _12105_/CLK line[64] vssd1 vssd1 vccd1 vccd1 _12076_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_1_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11026_ _11026_/A _11059_/Y vssd1 vssd1 vccd1 vccd1 _13826_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13137__D line[47] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MUX.M\[1\].MUX\[2\]_A1 _13688_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07135__D line[105] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12976__D line[87] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12977_ _12977_/A _12984_/Y vssd1 vssd1 vccd1 vccd1 _13817_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_17_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11928_ _11930_/CLK line[120] vssd1 vssd1 vccd1 vccd1 _11929_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_32_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11859_ _11859_/A _11864_/Y vssd1 vssd1 vccd1 vccd1 _13819_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_60_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05380_ _05380_/A _05389_/Y vssd1 vssd1 vccd1 vccd1 _13780_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_186_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13529_ _13529_/A _13544_/Y vssd1 vssd1 vccd1 vccd1 _13809_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13600__D line[116] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07050_ _07050_/A _07069_/Y vssd1 vssd1 vccd1 vccd1 _13770_/Z sky130_fd_sc_hd__ebufn_2
X_06001_ _06015_/CLK line[98] vssd1 vssd1 vccd1 vccd1 _06002_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06999__A _13909_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07952_ _07952_/A _07979_/Y vssd1 vssd1 vccd1 vccd1 _13832_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[17\].VALID\[12\].FF_D A[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06903_ _06925_/CLK line[13] vssd1 vssd1 vccd1 vccd1 _06904_/A sky130_fd_sc_hd__dfxtp_1
X_07883_ _07905_/CLK line[77] vssd1 vssd1 vccd1 vccd1 _07884_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[22\].CLKBUF\[1\] clk vssd1 vssd1 vccd1 vccd1 _08922_/CLK sky130_fd_sc_hd__clkbuf_4
X_09622_ _09622_/CLK _09623_/X vssd1 vssd1 vccd1 vccd1 _09620_/CLK sky130_fd_sc_hd__dlclkp_1
X_06834_ _06834_/A _06859_/Y vssd1 vssd1 vccd1 vccd1 _13834_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_83_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07045__D line[78] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12886__D line[60] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09553_ _13920_/Y wr vssd1 vssd1 vccd1 vccd1 _09553_/X sky130_fd_sc_hd__and2_1
XDATA\[12\].CLKBUF\[7\] clk vssd1 vssd1 vccd1 vccd1 _06052_/CLK sky130_fd_sc_hd__clkbuf_4
X_06765_ _06785_/CLK line[78] vssd1 vssd1 vccd1 vccd1 _06766_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_83_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11790__D line[57] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08504_ _13913_/X vssd1 vssd1 vccd1 vccd1 _08504_/Y sky130_fd_sc_hd__inv_2
XANTENNA__06884__D line[118] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05716_ _05716_/A _05739_/Y vssd1 vssd1 vccd1 vccd1 _13836_/Z sky130_fd_sc_hd__ebufn_2
X_09484_ _13920_/Y vssd1 vssd1 vccd1 vccd1 _09484_/Y sky130_fd_sc_hd__inv_2
XPHY_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06696_ _06696_/A _06719_/Y vssd1 vssd1 vccd1 vccd1 _13696_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09260__D line[52] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05143__A _13931_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08435_ _08465_/CLK line[64] vssd1 vssd1 vccd1 vccd1 _08436_/A sky130_fd_sc_hd__dfxtp_1
X_05647_ _05665_/CLK line[79] vssd1 vssd1 vccd1 vccd1 _05648_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[27\].VALID\[11\].FF_D A[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08366_ _08366_/A _08399_/Y vssd1 vssd1 vccd1 vccd1 _13686_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05578_ _05578_/A _05599_/Y vssd1 vssd1 vccd1 vccd1 _13698_/Z sky130_fd_sc_hd__ebufn_2
XDECH.DEC0.AND3 A_h[4] A_h[3] vssd1 vssd1 vccd1 vccd1 _13971_/D sky130_fd_sc_hd__and2_2
X_07317_ _07345_/CLK line[74] vssd1 vssd1 vccd1 vccd1 _07318_/A sky130_fd_sc_hd__dfxtp_1
X_08297_ _08325_/CLK line[10] vssd1 vssd1 vccd1 vccd1 _08298_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_192_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13510__D line[80] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07248_ _07248_/A _07279_/Y vssd1 vssd1 vccd1 vccd1 _13688_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_118_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12126__D line[82] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_DATA\[27\].CLKBUF\[3\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07179_ _07205_/CLK line[11] vssd1 vssd1 vccd1 vccd1 _07180_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12704__A _13936_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10190_ _10190_/A _10219_/Y vssd1 vssd1 vccd1 vccd1 _13830_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_105_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11965__D line[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[13\].VALID\[13\].TOBUF OVHB\[13\].VALID\[13\].FF/Q OVHB\[13\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04916_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__12423__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09435__D line[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05318__A _13900_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12900_ _12910_/CLK line[52] vssd1 vssd1 vccd1 vccd1 _12901_/A sky130_fd_sc_hd__dfxtp_1
X_13880_ _13890_/CLK line[116] vssd1 vssd1 vccd1 vccd1 _13881_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_100_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12831_ _12831_/A _12844_/Y vssd1 vssd1 vccd1 vccd1 _13671_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_74_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06794__D line[91] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12762_ _12770_/CLK line[117] vssd1 vssd1 vccd1 vccd1 _12763_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_203_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09170__D line[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11713_ _11713_/A _11724_/Y vssd1 vssd1 vccd1 vccd1 _13673_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12693_ _12693_/A _12704_/Y vssd1 vssd1 vccd1 vccd1 _13813_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XDATA\[11\].CLKBUF\[4\] clk vssd1 vssd1 vccd1 vccd1 _05667_/CLK sky130_fd_sc_hd__clkbuf_4
XPHY_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[28\].VALID\[2\].TOBUF OVHB\[28\].VALID\[2\].FF/Q OVHB\[28\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04930_/B2 sky130_fd_sc_hd__ebufn_2
XPHY_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11644_ _11650_/CLK line[118] vssd1 vssd1 vccd1 vccd1 _11645_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_14_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08364__A _13913_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[18\].INV _13955_/X vssd1 vssd1 vccd1 vccd1 OVHB\[18\].INV/Y sky130_fd_sc_hd__inv_2
XPHY_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11575_ _11575_/A _11584_/Y vssd1 vssd1 vccd1 vccd1 _13815_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08083__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13314_ _13330_/CLK line[113] vssd1 vssd1 vccd1 vccd1 _13315_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_6_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10526_ _10530_/CLK line[119] vssd1 vssd1 vccd1 vccd1 _10527_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[24\].VOBUF OVHB\[24\].V/Q OVHB\[24\].INV/Y vssd1 vssd1 vccd1 vccd1 _04912_/B1
+ sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[20\].VALID\[7\].FF_D A[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13245_ _13245_/A _13264_/Y vssd1 vssd1 vccd1 vccd1 _13805_/Z sky130_fd_sc_hd__ebufn_2
X_10457_ _10457_/A _10464_/Y vssd1 vssd1 vccd1 vccd1 _13817_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_182_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06034__D line[113] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13176_ _13190_/CLK line[50] vssd1 vssd1 vccd1 vccd1 _13177_/A sky130_fd_sc_hd__dfxtp_1
X_10388_ _10390_/CLK line[56] vssd1 vssd1 vccd1 vccd1 _10389_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11875__D line[110] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12127_ _12127_/A _12144_/Y vssd1 vssd1 vccd1 vccd1 _13807_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[0\].CLKBUF\[2\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06969__D line[43] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09345__D line[96] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05873__D line[40] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12058_ _12070_/CLK line[51] vssd1 vssd1 vccd1 vccd1 _12059_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_77_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11009_ _11009_/A _11024_/Y vssd1 vssd1 vccd1 vccd1 _13809_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08539__A _13913_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08258__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06550_ _06550_/A _06579_/Y vssd1 vssd1 vccd1 vccd1 _13830_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_93_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05501_ _05525_/CLK line[12] vssd1 vssd1 vccd1 vccd1 _05502_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_178_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06481_ _06505_/CLK line[76] vssd1 vssd1 vccd1 vccd1 _06482_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11115__D line[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08220_ _08220_/CLK line[89] vssd1 vssd1 vccd1 vccd1 _08221_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06209__D line[65] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05432_ _05432_/A _05459_/Y vssd1 vssd1 vccd1 vccd1 _13832_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_60_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05363_ _05385_/CLK line[77] vssd1 vssd1 vccd1 vccd1 _05364_/A sky130_fd_sc_hd__dfxtp_1
X_08151_ _08151_/A _08154_/Y vssd1 vssd1 vccd1 vccd1 _13751_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13330__D line[121] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07102_ _07102_/CLK _07103_/X vssd1 vssd1 vccd1 vccd1 _07100_/CLK sky130_fd_sc_hd__dlclkp_1
XDATA\[10\].CLKBUF\[1\] clk vssd1 vssd1 vccd1 vccd1 _05282_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__08424__D line[54] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08082_ _08082_/CLK _08083_/X vssd1 vssd1 vccd1 vccd1 _08080_/CLK sky130_fd_sc_hd__dlclkp_1
X_05294_ _05294_/A _05319_/Y vssd1 vssd1 vccd1 vccd1 _13694_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_119_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07033_ _13909_/Y wr vssd1 vssd1 vccd1 vccd1 _07033_/X sky130_fd_sc_hd__and2_1
XFILLER_161_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[20\].CG clk OVHB\[20\].CGAND/X vssd1 vssd1 vccd1 vccd1 OVHB\[20\].V/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_142_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10044__A _13922_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08984_ _08990_/CLK line[54] vssd1 vssd1 vccd1 vccd1 _08985_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05783__D line[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09833__A _13921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07935_ _07935_/A _07944_/Y vssd1 vssd1 vccd1 vccd1 _13815_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_68_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[1\].VALID\[2\].FF_D A[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07866_ _07870_/CLK line[55] vssd1 vssd1 vccd1 vccd1 _07867_/A sky130_fd_sc_hd__dfxtp_1
X_09605_ _09605_/A _09624_/Y vssd1 vssd1 vccd1 vccd1 _13805_/Z sky130_fd_sc_hd__ebufn_2
X_06817_ _06817_/A _06824_/Y vssd1 vssd1 vccd1 vccd1 _13817_/Z sky130_fd_sc_hd__ebufn_2
X_07797_ _07797_/A _07804_/Y vssd1 vssd1 vccd1 vccd1 _13677_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13505__D line[73] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09536_ _09550_/CLK line[50] vssd1 vssd1 vccd1 vccd1 _09537_/A sky130_fd_sc_hd__dfxtp_1
X_06748_ _06750_/CLK line[56] vssd1 vssd1 vccd1 vccd1 _06749_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_71_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09467_ _09467_/A _09484_/Y vssd1 vssd1 vccd1 vccd1 _13667_/Z sky130_fd_sc_hd__ebufn_2
X_06679_ _06679_/A _06684_/Y vssd1 vssd1 vccd1 vccd1 _13679_/Z sky130_fd_sc_hd__ebufn_2
XPHY_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11025__D line[96] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08418_ _08430_/CLK line[51] vssd1 vssd1 vccd1 vccd1 _08419_/A sky130_fd_sc_hd__dfxtp_1
X_09398_ _09410_/CLK line[115] vssd1 vssd1 vccd1 vccd1 _09399_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05023__D line[35] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10864__D line[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08349_ _08349_/A _08364_/Y vssd1 vssd1 vccd1 vccd1 _13669_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05958__D line[93] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13240__D line[94] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10219__A _13922_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[7\].VALID\[10\].FF OVHB\[7\].V/CLK A[17] vssd1 vssd1 vccd1 vccd1 OVHB\[7\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_22_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08334__D line[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11360_ _11370_/CLK line[116] vssd1 vssd1 vccd1 vccd1 _11361_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_164_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_MUX.M\[3\].MUX\[3\]_A3 _13865_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10311_ _10311_/A _10324_/Y vssd1 vssd1 vccd1 vccd1 _13671_/Z sky130_fd_sc_hd__ebufn_2
X_11291_ _11291_/A _11304_/Y vssd1 vssd1 vccd1 vccd1 _13811_/Z sky130_fd_sc_hd__ebufn_2
X_13030_ _13050_/CLK line[126] vssd1 vssd1 vccd1 vccd1 _13031_/A sky130_fd_sc_hd__dfxtp_1
X_10242_ _10250_/CLK line[117] vssd1 vssd1 vccd1 vccd1 _10243_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_140_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XOVHB\[1\].VALID\[4\].TOBUF OVHB\[1\].VALID\[4\].FF/Q OVHB\[1\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04925_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_79_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10173_ _10173_/A _10184_/Y vssd1 vssd1 vccd1 vccd1 _13813_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09165__D line[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[26\].VALID\[7\].TOBUF OVHB\[26\].VALID\[7\].FF/Q OVHB\[26\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/A2 sky130_fd_sc_hd__ebufn_2
XFILLER_121_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_DATA\[25\].CLKBUF\[5\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10104__D line[54] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13932_ _13938_/C _13938_/B _13938_/A _13938_/D vssd1 vssd1 vccd1 vccd1 _13932_/X
+ sky130_fd_sc_hd__and4bb_4
XFILLER_19_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13863_ _13863_/A _13894_/Y vssd1 vssd1 vccd1 vccd1 _13863_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13415__D line[46] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12814_ _12840_/CLK line[27] vssd1 vssd1 vccd1 vccd1 _12815_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08509__D line[107] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13794_ _13820_/CLK line[91] vssd1 vssd1 vccd1 vccd1 _13795_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07413__D line[104] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12745_ _12745_/A _12774_/Y vssd1 vssd1 vccd1 vccd1 _13865_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_15_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11513__A _13926_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12676_ _12700_/CLK line[92] vssd1 vssd1 vccd1 vccd1 _12677_/A sky130_fd_sc_hd__dfxtp_1
XPHY_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11627_ _11627_/A _11654_/Y vssd1 vssd1 vccd1 vccd1 _13867_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_30_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11558_ _11580_/CLK line[93] vssd1 vssd1 vccd1 vccd1 _11559_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_7_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XOVHB\[18\].VALID\[2\].FF OVHB\[18\].V/CLK A[9] vssd1 vssd1 vccd1 vccd1 OVHB\[18\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_155_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10509_ _10509_/A _10534_/Y vssd1 vssd1 vccd1 vccd1 _13869_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_183_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11489_ _11489_/A _11514_/Y vssd1 vssd1 vccd1 vccd1 _13729_/Z sky130_fd_sc_hd__ebufn_2
X_13228_ _13938_/X wr vssd1 vssd1 vccd1 vccd1 _13228_/X sky130_fd_sc_hd__and2_1
XFILLER_112_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06699__D line[33] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13159_ _13938_/X vssd1 vssd1 vccd1 vccd1 _13159_/Y sky130_fd_sc_hd__inv_2
XFILLER_170_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09075__D line[110] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05981_ _05981_/A _05984_/Y vssd1 vssd1 vccd1 vccd1 _13821_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_38_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10014__D line[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07720_ _07730_/CLK line[116] vssd1 vssd1 vccd1 vccd1 _07721_/A sky130_fd_sc_hd__dfxtp_1
X_04932_ A_h[15] _04932_/B2 A_h[15] _04932_/B2 vssd1 vssd1 vccd1 vccd1 _04933_/D sky130_fd_sc_hd__a2bb2oi_2
XANTENNA__07173__A _13909_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07651_ _07651_/A _07664_/Y vssd1 vssd1 vccd1 vccd1 _13811_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_81_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06602_ _06610_/CLK line[117] vssd1 vssd1 vccd1 vccd1 _06603_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__04947__D line[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[7\].VALID\[6\].FF_D A[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07582_ _07590_/CLK line[53] vssd1 vssd1 vccd1 vccd1 _07583_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07323__D line[77] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09321_ _09321_/A _09344_/Y vssd1 vssd1 vccd1 vccd1 _13801_/Z sky130_fd_sc_hd__ebufn_2
X_06533_ _06533_/A _06544_/Y vssd1 vssd1 vccd1 vccd1 _13813_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_179_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09252_ _09270_/CLK line[63] vssd1 vssd1 vccd1 vccd1 _09253_/A sky130_fd_sc_hd__dfxtp_1
X_06464_ _06470_/CLK line[54] vssd1 vssd1 vccd1 vccd1 _06465_/A sky130_fd_sc_hd__dfxtp_1
X_08203_ _08203_/A _08224_/Y vssd1 vssd1 vccd1 vccd1 _13803_/Z sky130_fd_sc_hd__ebufn_2
X_05415_ _05415_/A _05424_/Y vssd1 vssd1 vccd1 vccd1 _13815_/Z sky130_fd_sc_hd__ebufn_2
X_09183_ _09183_/A _09204_/Y vssd1 vssd1 vccd1 vccd1 _13663_/Z sky130_fd_sc_hd__ebufn_2
X_06395_ _06395_/A _06404_/Y vssd1 vssd1 vccd1 vccd1 _13675_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[7\].VALID\[10\].TOBUF OVHB\[7\].VALID\[10\].FF/Q OVHB\[7\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04932_/B2 sky130_fd_sc_hd__ebufn_2
X_08134_ _08150_/CLK line[49] vssd1 vssd1 vccd1 vccd1 _08135_/A sky130_fd_sc_hd__dfxtp_1
X_05346_ _05350_/CLK line[55] vssd1 vssd1 vccd1 vccd1 _05347_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_162_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08065_ _08065_/A _08084_/Y vssd1 vssd1 vccd1 vccd1 _13665_/Z sky130_fd_sc_hd__ebufn_2
X_05277_ _05277_/A _05284_/Y vssd1 vssd1 vccd1 vccd1 _13677_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_146_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07348__A _13910_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07016_ _07030_/CLK line[50] vssd1 vssd1 vccd1 vccd1 _07017_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_103_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12404__D line[81] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[16\].VALID\[4\].FF OVHB\[16\].V/CLK A[11] vssd1 vssd1 vccd1 vccd1 OVHB\[16\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_08967_ _08967_/A _08994_/Y vssd1 vssd1 vccd1 vccd1 _13727_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_194_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07918_ _07940_/CLK line[93] vssd1 vssd1 vccd1 vccd1 _07919_/A sky130_fd_sc_hd__dfxtp_1
X_08898_ _08920_/CLK line[29] vssd1 vssd1 vccd1 vccd1 _08899_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09713__D line[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07849_ _07849_/A _07874_/Y vssd1 vssd1 vccd1 vccd1 _13729_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[10\].V_RESET_B rst_n vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10860_ _10880_/CLK line[30] vssd1 vssd1 vccd1 vccd1 _10861_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_71_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09519_ _13920_/Y vssd1 vssd1 vccd1 vccd1 _09519_/Y sky130_fd_sc_hd__inv_2
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10791_ _10791_/A _10814_/Y vssd1 vssd1 vccd1 vccd1 _13871_/Z sky130_fd_sc_hd__ebufn_2
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_OVHB\[27\].CGAND_B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12530_ _12560_/CLK line[16] vssd1 vssd1 vccd1 vccd1 _12531_/A sky130_fd_sc_hd__dfxtp_1
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10594__D line[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12461_ _12461_/A _12494_/Y vssd1 vssd1 vccd1 vccd1 _13861_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05688__D line[83] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11412_ _11440_/CLK line[26] vssd1 vssd1 vccd1 vccd1 _11413_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08064__D line[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12392_ _12420_/CLK line[90] vssd1 vssd1 vccd1 vccd1 _12393_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_193_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11343_ _11343_/A _11374_/Y vssd1 vssd1 vccd1 vccd1 _13863_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08999__D line[75] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11274_ _11300_/CLK line[91] vssd1 vssd1 vccd1 vccd1 _11275_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.M\[2\].MUX\[4\]_A1 _13741_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13013_ _13015_/CLK line[104] vssd1 vssd1 vccd1 vccd1 _13014_/A sky130_fd_sc_hd__dfxtp_1
X_10225_ _10225_/A _10254_/Y vssd1 vssd1 vccd1 vccd1 _13865_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_3_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06312__D line[127] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10156_ _10180_/CLK line[92] vssd1 vssd1 vccd1 vccd1 _10157_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_58_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10087_ _10087_/A _10114_/Y vssd1 vssd1 vccd1 vccd1 _13727_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10769__D line[102] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[29\].V_RESET_B rst_n vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13915_ _13916_/A _13916_/B _13916_/C _13916_/D vssd1 vssd1 vccd1 vccd1 _13915_/X
+ sky130_fd_sc_hd__and4b_4
XFILLER_208_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13145__D line[36] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08239__D line[97] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13846_ _13846_/A _13859_/Y vssd1 vssd1 vccd1 vccd1 _13846_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[14\].VALID\[6\].FF OVHB\[14\].V/CLK A[13] vssd1 vssd1 vccd1 vccd1 OVHB\[14\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[23\].CLKBUF\[7\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13777_ _13785_/CLK line[69] vssd1 vssd1 vccd1 vccd1 _13778_/A sky130_fd_sc_hd__dfxtp_1
X_10989_ _13925_/X vssd1 vssd1 vccd1 vccd1 _10989_/Y sky130_fd_sc_hd__inv_2
X_12728_ _12728_/A _12739_/Y vssd1 vssd1 vccd1 vccd1 _13848_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.M\[0\].MUX\[0\]_A2 _13756_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12659_ _12665_/CLK line[70] vssd1 vssd1 vccd1 vccd1 _12660_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05200_ _05210_/CLK line[116] vssd1 vssd1 vccd1 vccd1 _05201_/A sky130_fd_sc_hd__dfxtp_1
X_06180_ _06190_/CLK line[52] vssd1 vssd1 vccd1 vccd1 _06181_/A sky130_fd_sc_hd__dfxtp_1
X_05131_ _05131_/A _05144_/Y vssd1 vssd1 vccd1 vccd1 _13811_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_156_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12074__A _13934_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05062_ _05070_/CLK line[53] vssd1 vssd1 vccd1 vccd1 _05063_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08702__D line[53] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09870_ _09900_/CLK line[80] vssd1 vssd1 vccd1 vccd1 _09871_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_140_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08821_ _08821_/A _08854_/Y vssd1 vssd1 vccd1 vccd1 _13861_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_97_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XOVHB\[8\].VALID\[4\].TOBUF OVHB\[8\].VALID\[4\].FF/Q OVHB\[8\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04925_/B2 sky130_fd_sc_hd__ebufn_2
X_08752_ _08780_/CLK line[90] vssd1 vssd1 vccd1 vccd1 _08753_/A sky130_fd_sc_hd__dfxtp_1
X_05964_ _05980_/CLK line[81] vssd1 vssd1 vccd1 vccd1 _05965_/A sky130_fd_sc_hd__dfxtp_1
X_07703_ _07703_/A _07734_/Y vssd1 vssd1 vccd1 vccd1 _13863_/Z sky130_fd_sc_hd__ebufn_2
X_04915_ A_h[16] _04915_/B2 A_h[16] _04915_/B2 vssd1 vssd1 vccd1 vccd1 _04917_/C sky130_fd_sc_hd__a2bb2oi_2
XANTENNA__10679__D line[75] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08683_ _08683_/A _08714_/Y vssd1 vssd1 vccd1 vccd1 _13723_/Z sky130_fd_sc_hd__ebufn_2
X_05895_ _05895_/A _05914_/Y vssd1 vssd1 vccd1 vccd1 _13735_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13055__D line[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07634_ _07660_/CLK line[91] vssd1 vssd1 vccd1 vccd1 _07635_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07053__D line[67] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12894__D line[49] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07565_ _07565_/A _07594_/Y vssd1 vssd1 vccd1 vccd1 _13725_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12249__A _13935_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07988__D line[125] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09304_ _09304_/A _09309_/Y vssd1 vssd1 vccd1 vccd1 _13784_/Z sky130_fd_sc_hd__ebufn_2
X_06516_ _06540_/CLK line[92] vssd1 vssd1 vccd1 vccd1 _06517_/A sky130_fd_sc_hd__dfxtp_1
X_07496_ _07520_/CLK line[28] vssd1 vssd1 vccd1 vccd1 _07497_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_21_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XOVHB\[23\].VALID\[11\].TOBUF OVHB\[23\].VALID\[11\].FF/Q OVHB\[23\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04915_/B2 sky130_fd_sc_hd__ebufn_2
X_09235_ _09235_/CLK line[41] vssd1 vssd1 vccd1 vccd1 _09236_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_139_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06447_ _06447_/A _06474_/Y vssd1 vssd1 vccd1 vccd1 _13727_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[1\].CLKBUF\[5\] clk vssd1 vssd1 vccd1 vccd1 _08222_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_166_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[12\].VALID\[8\].FF OVHB\[12\].V/CLK A[15] vssd1 vssd1 vccd1 vccd1 OVHB\[12\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_166_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09166_ _09166_/A _09169_/Y vssd1 vssd1 vccd1 vccd1 _13646_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_166_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06378_ _06400_/CLK line[29] vssd1 vssd1 vccd1 vccd1 _06379_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05301__D line[34] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08117_ _08117_/CLK _08118_/X vssd1 vssd1 vccd1 vccd1 _08115_/CLK sky130_fd_sc_hd__dlclkp_1
X_05329_ _05329_/A _05354_/Y vssd1 vssd1 vccd1 vccd1 _13729_/Z sky130_fd_sc_hd__ebufn_2
X_09097_ _09097_/CLK _09098_/X vssd1 vssd1 vccd1 vccd1 _09095_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_79_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08048_ _13932_/X wr vssd1 vssd1 vccd1 vccd1 _08048_/X sky130_fd_sc_hd__and2_1
XANTENNA__08612__D line[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12134__D line[86] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07228__D line[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10010_ _10040_/CLK line[16] vssd1 vssd1 vccd1 vccd1 _10011_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09999_ _10005_/CLK line[6] vssd1 vssd1 vccd1 vccd1 _10000_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_130_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09443__D line[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XDATA\[31\].CLKBUF\[3\] clk vssd1 vssd1 vccd1 vccd1 _11792_/CLK sky130_fd_sc_hd__clkbuf_4
X_11961_ _11965_/CLK line[7] vssd1 vssd1 vccd1 vccd1 _11962_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_91_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13700_ _13700_/A _13719_/Y vssd1 vssd1 vccd1 vccd1 _13700_/Z sky130_fd_sc_hd__ebufn_2
X_10912_ _10912_/A _10919_/Y vssd1 vssd1 vccd1 vccd1 _13712_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13543__A _13898_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11892_ _11892_/A _11899_/Y vssd1 vssd1 vccd1 vccd1 _13852_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_44_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13631_ _13645_/CLK line[2] vssd1 vssd1 vccd1 vccd1 _13632_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[12\].VALID\[2\].FF_D A[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10843_ _10845_/CLK line[8] vssd1 vssd1 vccd1 vccd1 _10844_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_198_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13562_ _13562_/A _13579_/Y vssd1 vssd1 vccd1 vccd1 _13842_/Z sky130_fd_sc_hd__ebufn_2
X_10774_ _10774_/A _10779_/Y vssd1 vssd1 vccd1 vccd1 _13854_/Z sky130_fd_sc_hd__ebufn_2
X_12513_ _12525_/CLK line[3] vssd1 vssd1 vccd1 vccd1 _12514_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12309__D line[38] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13493_ _13505_/CLK line[67] vssd1 vssd1 vccd1 vccd1 _13494_/A sky130_fd_sc_hd__dfxtp_1
X_12444_ _12444_/A _12459_/Y vssd1 vssd1 vccd1 vccd1 _13844_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_145_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12375_ _12385_/CLK line[68] vssd1 vssd1 vccd1 vccd1 _12376_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[0\].CLKBUF\[2\] clk vssd1 vssd1 vccd1 vccd1 _05037_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__09618__D line[88] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11326_ _11326_/A _11339_/Y vssd1 vssd1 vccd1 vccd1 _13846_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_141_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13718__A _13899_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12044__D line[59] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11257_ _11265_/CLK line[69] vssd1 vssd1 vccd1 vccd1 _11258_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[25\].V OVHB\[25\].V/CLK TIE/HI rst_n vssd1 vssd1 vccd1 vccd1 OVHB\[25\].V/Q
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_95_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06042__D line[117] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10208_ _10208_/A _10219_/Y vssd1 vssd1 vccd1 vccd1 _13848_/Z sky130_fd_sc_hd__ebufn_2
X_11188_ _11188_/A _11199_/Y vssd1 vssd1 vccd1 vccd1 _13708_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11883__D line[99] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06977__D line[47] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10139_ _10145_/CLK line[70] vssd1 vssd1 vccd1 vccd1 _10140_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__04927__B2 _04927_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09353__D line[109] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[3\].VALID\[9\].FF_D A[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05680_ _05700_/CLK line[94] vssd1 vssd1 vccd1 vccd1 _05681_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_62_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13829_ _13855_/CLK line[107] vssd1 vssd1 vccd1 vccd1 _13830_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[30\].CLKBUF\[0\] clk vssd1 vssd1 vccd1 vccd1 _11407_/CLK sky130_fd_sc_hd__clkbuf_4
X_07350_ _07380_/CLK line[80] vssd1 vssd1 vccd1 vccd1 _07351_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07601__D line[76] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06301_ _06301_/A _06334_/Y vssd1 vssd1 vccd1 vccd1 _13861_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[20\].CLKBUF\[6\] clk vssd1 vssd1 vccd1 vccd1 _08537_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_149_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12219__D line[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07281_ _07281_/A _07314_/Y vssd1 vssd1 vccd1 vccd1 _13721_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11123__D line[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09020_ _09020_/A _09029_/Y vssd1 vssd1 vccd1 vccd1 _13780_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09378__A _13916_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06232_ _06260_/CLK line[90] vssd1 vssd1 vccd1 vccd1 _06233_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_191_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06217__D line[69] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XOVHB\[6\].VALID\[9\].TOBUF OVHB\[6\].VALID\[9\].FF/Q OVHB\[6\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04914_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[4\].VALID\[11\].FF_D A[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06163_ _06163_/A _06194_/Y vssd1 vssd1 vccd1 vccd1 _13723_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09528__D line[61] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05114_ _05140_/CLK line[91] vssd1 vssd1 vccd1 vccd1 _05115_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_116_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06094_ _06120_/CLK line[27] vssd1 vssd1 vccd1 vccd1 _06095_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_116_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05045_ _05045_/A _05074_/Y vssd1 vssd1 vccd1 vccd1 _13725_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_116_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09922_ _09922_/A _09939_/Y vssd1 vssd1 vccd1 vccd1 _13842_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[16\].V OVHB\[16\].V/CLK TIE/HI rst_n vssd1 vssd1 vccd1 vccd1 OVHB\[16\].V/Q
+ sky130_fd_sc_hd__dfrtp_1
X_09853_ _09865_/CLK line[67] vssd1 vssd1 vccd1 vccd1 _09854_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_112_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08804_ _08804_/A _08819_/Y vssd1 vssd1 vccd1 vccd1 _13844_/Z sky130_fd_sc_hd__ebufn_2
X_09784_ _09784_/A _09799_/Y vssd1 vssd1 vccd1 vccd1 _13704_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05791__D line[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06996_ _06996_/A _06999_/Y vssd1 vssd1 vccd1 vccd1 _13716_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_105_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08735_ _08745_/CLK line[68] vssd1 vssd1 vccd1 vccd1 _08736_/A sky130_fd_sc_hd__dfxtp_1
X_05947_ _05947_/CLK _05948_/X vssd1 vssd1 vccd1 vccd1 _05945_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_27_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_OVHB\[25\].VALID\[2\].FF_D A[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08666_ _08666_/A _08679_/Y vssd1 vssd1 vccd1 vccd1 _13706_/Z sky130_fd_sc_hd__ebufn_2
X_05878_ _13902_/X wr vssd1 vssd1 vccd1 vccd1 _05878_/X sky130_fd_sc_hd__and2_1
XPHY_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07617_ _07625_/CLK line[69] vssd1 vssd1 vccd1 vccd1 _07618_/A sky130_fd_sc_hd__dfxtp_1
X_08597_ _08605_/CLK line[5] vssd1 vssd1 vccd1 vccd1 _08598_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07548_ _07548_/A _07559_/Y vssd1 vssd1 vccd1 vccd1 _13708_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[18\].VALID\[6\].FF_D A[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07479_ _07485_/CLK line[6] vssd1 vssd1 vccd1 vccd1 _07480_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11033__D line[109] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09218_ _09218_/A _09239_/Y vssd1 vssd1 vccd1 vccd1 _13698_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_14_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06127__D line[42] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10490_ _10490_/A _10499_/Y vssd1 vssd1 vccd1 vccd1 _13850_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05031__D line[39] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[5\].VALID\[1\].FF OVHB\[5\].V/CLK A[8] vssd1 vssd1 vccd1 vccd1 OVHB\[5\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_09149_ _09165_/CLK line[1] vssd1 vssd1 vccd1 vccd1 _09150_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10872__D line[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05966__D line[82] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12160_ _12160_/A _12179_/Y vssd1 vssd1 vccd1 vccd1 _13840_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08342__D line[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11111_ _11125_/CLK line[2] vssd1 vssd1 vccd1 vccd1 _11112_/A sky130_fd_sc_hd__dfxtp_1
X_12091_ _12105_/CLK line[66] vssd1 vssd1 vccd1 vccd1 _12092_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_104_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11042_ _11042_/A _11059_/Y vssd1 vssd1 vccd1 vccd1 _13842_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12799__D line[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XOVHB\[13\].VALID\[4\].TOBUF OVHB\[13\].VALID\[4\].FF/Q OVHB\[13\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04925_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_76_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11058__A _13925_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11208__D line[61] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12993_ _13015_/CLK line[109] vssd1 vssd1 vccd1 vccd1 _12994_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_29_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11944_ _11944_/A _11969_/Y vssd1 vssd1 vccd1 vccd1 _13624_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_55_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05206__D line[119] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11875_ _11895_/CLK line[110] vssd1 vssd1 vccd1 vccd1 _11876_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_32_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13423__D line[35] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13614_ _13898_/Y vssd1 vssd1 vccd1 vccd1 _13614_/Y sky130_fd_sc_hd__inv_2
X_10826_ _10826_/A _10849_/Y vssd1 vssd1 vccd1 vccd1 _13626_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_60_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08517__D line[111] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10757_ _10775_/CLK line[111] vssd1 vssd1 vccd1 vccd1 _10758_/A sky130_fd_sc_hd__dfxtp_1
X_13545_ _13575_/CLK line[96] vssd1 vssd1 vccd1 vccd1 _13546_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_201_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13476_ _13476_/A _13509_/Y vssd1 vssd1 vccd1 vccd1 _13756_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_9_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10688_ _10688_/A _10709_/Y vssd1 vssd1 vccd1 vccd1 _13768_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10782__D line[122] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12427_ _12455_/CLK line[106] vssd1 vssd1 vccd1 vccd1 _12428_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[16\].CLKBUF\[1\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12358_ _12358_/A _12389_/Y vssd1 vssd1 vccd1 vccd1 _13758_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_126_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11309_ _11335_/CLK line[107] vssd1 vssd1 vccd1 vccd1 _11310_/A sky130_fd_sc_hd__dfxtp_1
X_12289_ _12315_/CLK line[43] vssd1 vssd1 vccd1 vccd1 _12290_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_113_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XOVHB\[3\].VALID\[3\].FF OVHB\[3\].V/CLK A[10] vssd1 vssd1 vccd1 vccd1 OVHB\[3\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_141_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06850_ _06850_/A _06859_/Y vssd1 vssd1 vccd1 vccd1 _13850_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09083__D line[99] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05801_ _05805_/CLK line[7] vssd1 vssd1 vccd1 vccd1 _05802_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_95_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06781_ _06785_/CLK line[71] vssd1 vssd1 vccd1 vccd1 _06782_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_209_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10022__D line[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08520_ _08520_/A _08539_/Y vssd1 vssd1 vccd1 vccd1 _13840_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[19\].VOBUF OVHB\[19\].V/Q OVHB\[19\].INV/Y vssd1 vssd1 vccd1 vccd1 _04912_/B1
+ sky130_fd_sc_hd__ebufn_2
X_05732_ _05732_/A _05739_/Y vssd1 vssd1 vccd1 vccd1 _13852_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_36_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05116__D line[92] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[9\].CLKBUF\[1\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08451_ _08465_/CLK line[66] vssd1 vssd1 vccd1 vccd1 _08452_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10957__D line[74] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05663_ _05665_/CLK line[72] vssd1 vssd1 vccd1 vccd1 _05664_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_35_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07402_ _07402_/A _07419_/Y vssd1 vssd1 vccd1 vccd1 _13842_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__04955__D line[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08382_ _08382_/A _08399_/Y vssd1 vssd1 vccd1 vccd1 _13702_/Z sky130_fd_sc_hd__ebufn_2
X_05594_ _05594_/A _05599_/Y vssd1 vssd1 vccd1 vccd1 _13714_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_50_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07331__D line[66] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07333_ _07345_/CLK line[67] vssd1 vssd1 vccd1 vccd1 _07334_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_109_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07264_ _07264_/A _07279_/Y vssd1 vssd1 vccd1 vccd1 _13704_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11788__D line[56] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09003_ _09025_/CLK line[77] vssd1 vssd1 vccd1 vccd1 _09004_/A sky130_fd_sc_hd__dfxtp_1
X_06215_ _06225_/CLK line[68] vssd1 vssd1 vccd1 vccd1 _06216_/A sky130_fd_sc_hd__dfxtp_1
X_07195_ _07205_/CLK line[4] vssd1 vssd1 vccd1 vccd1 _07196_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09258__D line[51] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06146_ _06146_/A _06159_/Y vssd1 vssd1 vccd1 vccd1 _13706_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_105_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06077_ _06085_/CLK line[5] vssd1 vssd1 vccd1 vccd1 _06078_/A sky130_fd_sc_hd__dfxtp_1
X_05028_ _05028_/A _05039_/Y vssd1 vssd1 vccd1 vccd1 _13708_/Z sky130_fd_sc_hd__ebufn_2
X_09905_ _09935_/CLK line[96] vssd1 vssd1 vccd1 vccd1 _09906_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12412__D line[85] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09836_ _09836_/A _09869_/Y vssd1 vssd1 vccd1 vccd1 _13756_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07506__D line[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06979_ _06995_/CLK line[33] vssd1 vssd1 vccd1 vccd1 _06980_/A sky130_fd_sc_hd__dfxtp_1
X_09767_ _09795_/CLK line[42] vssd1 vssd1 vccd1 vccd1 _09768_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07803__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08718_ _08718_/A _08749_/Y vssd1 vssd1 vccd1 vccd1 _13758_/Z sky130_fd_sc_hd__ebufn_2
X_09698_ _09698_/A _09729_/Y vssd1 vssd1 vccd1 vccd1 _13618_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09721__D line[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[1\].VALID\[5\].FF OVHB\[1\].V/CLK A[12] vssd1 vssd1 vccd1 vccd1 OVHB\[1\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08649_ _08675_/CLK line[43] vssd1 vssd1 vccd1 vccd1 _08650_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11660_ _11660_/A _11689_/Y vssd1 vssd1 vccd1 vccd1 _13620_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10611_ _10635_/CLK line[44] vssd1 vssd1 vccd1 vccd1 _10612_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11591_ _11615_/CLK line[108] vssd1 vssd1 vccd1 vccd1 _11592_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XOVHB\[11\].VALID\[9\].TOBUF OVHB\[11\].VALID\[9\].FF/Q OVHB\[11\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04914_/B2 sky130_fd_sc_hd__ebufn_2
XPHY_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13330_ _13330_/CLK line[121] vssd1 vssd1 vccd1 vccd1 _13331_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_183_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10542_ _10542_/A _10569_/Y vssd1 vssd1 vccd1 vccd1 _13622_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MUX.M\[3\].MUX\[6\]_A1 _13731_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11698__D line[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13261_ _13261_/A _13264_/Y vssd1 vssd1 vccd1 vccd1 _13821_/Z sky130_fd_sc_hd__ebufn_2
X_10473_ _10495_/CLK line[109] vssd1 vssd1 vccd1 vccd1 _10474_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_182_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05696__D line[87] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12212_ _12212_/CLK _12213_/X vssd1 vssd1 vccd1 vccd1 _12210_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__08072__D line[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13192_ _13192_/CLK _13193_/X vssd1 vssd1 vccd1 vccd1 _13190_/CLK sky130_fd_sc_hd__dlclkp_1
X_12143_ _13934_/X wr vssd1 vssd1 vccd1 vccd1 _12143_/X sky130_fd_sc_hd__and2_1
X_12074_ _13934_/X vssd1 vssd1 vccd1 vccd1 _12074_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12322__D line[58] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11025_ _11055_/CLK line[96] vssd1 vssd1 vccd1 vccd1 _11026_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06320__D line[116] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_MUX.M\[1\].MUX\[2\]_A2 _13758_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[20\].VOBUF OVHB\[20\].V/Q OVHB\[20\].INV/Y vssd1 vssd1 vccd1 vccd1 _04912_/B1
+ sky130_fd_sc_hd__ebufn_2
XFILLER_80_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12976_ _12980_/CLK line[87] vssd1 vssd1 vccd1 vccd1 _12977_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09631__D line[108] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11927_ _11927_/A _11934_/Y vssd1 vssd1 vccd1 vccd1 _13887_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_205_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13153__D line[40] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08247__D line[101] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11858_ _11860_/CLK line[88] vssd1 vssd1 vccd1 vccd1 _11859_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_82_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10809_ _10809_/A _10814_/Y vssd1 vssd1 vccd1 vccd1 _13889_/Z sky130_fd_sc_hd__ebufn_2
X_11789_ _11789_/A _11794_/Y vssd1 vssd1 vccd1 vccd1 _13749_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_9_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13528_ _13540_/CLK line[83] vssd1 vssd1 vccd1 vccd1 _13529_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_118_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13459_ _13459_/A _13474_/Y vssd1 vssd1 vccd1 vccd1 _13739_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11401__D line[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06000_ _06000_/A _06019_/Y vssd1 vssd1 vccd1 vccd1 _13840_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09055__TE_B _09064_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09806__D line[60] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08710__D line[57] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07951_ _07975_/CLK line[108] vssd1 vssd1 vccd1 vccd1 _07952_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_141_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13328__D line[120] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06902_ _06902_/A _06929_/Y vssd1 vssd1 vccd1 vccd1 _13622_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[14\].CLKBUF\[3\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13906__A A[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07882_ _07882_/A _07909_/Y vssd1 vssd1 vccd1 vccd1 _13762_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[21\].VALID\[5\].FF_D A[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09621_ _09621_/A _09624_/Y vssd1 vssd1 vccd1 vccd1 _13821_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[28\].VALID\[0\].FF OVHB\[28\].V/CLK A[7] vssd1 vssd1 vccd1 vccd1 OVHB\[28\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06230__D line[80] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06833_ _06855_/CLK line[109] vssd1 vssd1 vccd1 vccd1 _06834_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_28_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09552_ _09552_/CLK _09553_/X vssd1 vssd1 vccd1 vccd1 _09550_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_209_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06764_ _06764_/A _06789_/Y vssd1 vssd1 vccd1 vccd1 _13764_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_102_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08503_ _13913_/X wr vssd1 vssd1 vccd1 vccd1 _08503_/X sky130_fd_sc_hd__and2_1
XANTENNA__05424__A _13900_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10687__D line[79] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05715_ _05735_/CLK line[110] vssd1 vssd1 vccd1 vccd1 _05716_/A sky130_fd_sc_hd__dfxtp_1
X_09483_ _13920_/Y wr vssd1 vssd1 vccd1 vccd1 _09483_/X sky130_fd_sc_hd__and2_1
X_06695_ _06715_/CLK line[46] vssd1 vssd1 vccd1 vccd1 _06696_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13063__D line[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[14\].VALID\[9\].FF_D A[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05143__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08434_ _13913_/X vssd1 vssd1 vccd1 vccd1 _08434_/Y sky130_fd_sc_hd__inv_2
X_05646_ _05646_/A _05669_/Y vssd1 vssd1 vccd1 vccd1 _13766_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08157__D line[74] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07061__D line[71] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08365_ _08395_/CLK line[32] vssd1 vssd1 vccd1 vccd1 _08366_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05577_ _05595_/CLK line[47] vssd1 vssd1 vccd1 vccd1 _05578_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07996__D line[114] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07316_ _07316_/A _07349_/Y vssd1 vssd1 vccd1 vccd1 _13756_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[7\].CLKBUF\[3\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08296_ _08296_/A _08329_/Y vssd1 vssd1 vccd1 vccd1 _13616_/Z sky130_fd_sc_hd__ebufn_2
X_07247_ _07275_/CLK line[42] vssd1 vssd1 vccd1 vccd1 _07248_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11311__D line[108] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06405__D line[32] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07178_ _07178_/A _07209_/Y vssd1 vssd1 vccd1 vccd1 _13618_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_133_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13088__A _13938_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06129_ _06155_/CLK line[43] vssd1 vssd1 vccd1 vccd1 _06130_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_87_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08620__D line[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[11\].VALID\[13\].FF_D A[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13238__D line[93] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05318__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07236__D line[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[19\].CG_CLK clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09819_ _09819_/A _09834_/Y vssd1 vssd1 vccd1 vccd1 _13739_/Z sky130_fd_sc_hd__ebufn_2
X_12830_ _12840_/CLK line[20] vssd1 vssd1 vccd1 vccd1 _12831_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_36_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12761_ _12761_/A _12774_/Y vssd1 vssd1 vccd1 vccd1 _13881_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11712_ _11720_/CLK line[21] vssd1 vssd1 vccd1 vccd1 _11713_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_199_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12692_ _12700_/CLK line[85] vssd1 vssd1 vccd1 vccd1 _12693_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[26\].VALID\[2\].FF OVHB\[26\].V/CLK A[9] vssd1 vssd1 vccd1 vccd1 OVHB\[26\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[21\].VALID\[12\].FF_D A[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[1\].VALID\[0\].TOBUF OVHB\[1\].VALID\[0\].FF/Q OVHB\[1\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04924_/B2 sky130_fd_sc_hd__ebufn_2
XPHY_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11643_ _11643_/A _11654_/Y vssd1 vssd1 vccd1 vccd1 _13883_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[2\].VALID\[0\].FF_D A[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[26\].VALID\[3\].TOBUF OVHB\[26\].VALID\[3\].FF/Q OVHB\[26\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04919_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__13701__D line[34] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11574_ _11580_/CLK line[86] vssd1 vssd1 vccd1 vccd1 _11575_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10525_ _10525_/A _10534_/Y vssd1 vssd1 vccd1 vccd1 _13885_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_168_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13313_ _13313_/A _13334_/Y vssd1 vssd1 vccd1 vccd1 _13873_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_155_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13244_ _13260_/CLK line[81] vssd1 vssd1 vccd1 vccd1 _13245_/A sky130_fd_sc_hd__dfxtp_1
X_10456_ _10460_/CLK line[87] vssd1 vssd1 vccd1 vccd1 _10457_/A sky130_fd_sc_hd__dfxtp_1
X_13175_ _13175_/A _13194_/Y vssd1 vssd1 vccd1 vccd1 _13735_/Z sky130_fd_sc_hd__ebufn_2
X_10387_ _10387_/A _10394_/Y vssd1 vssd1 vccd1 vccd1 _13747_/Z sky130_fd_sc_hd__ebufn_2
X_12126_ _12140_/CLK line[82] vssd1 vssd1 vccd1 vccd1 _12127_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[31\].VALID\[11\].FF_D A[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12052__D line[63] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12057_ _12057_/A _12074_/Y vssd1 vssd1 vccd1 vccd1 _13737_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_111_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07146__D line[124] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[13\].V_D TIE/HI vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06050__D line[121] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11008_ _11020_/CLK line[83] vssd1 vssd1 vccd1 vccd1 _11009_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12987__D line[106] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11891__D line[103] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06985__D line[36] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[27\].CGAND _13923_/X wr vssd1 vssd1 vccd1 vccd1 OVHB\[27\].CGAND/X sky130_fd_sc_hd__and2_4
XANTENNA_OVHB\[27\].VALID\[9\].FF_D A[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09361__D line[98] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_OVHB\[28\].V_D TIE/HI vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12959_ _12959_/A _12984_/Y vssd1 vssd1 vccd1 vccd1 _13799_/Z sky130_fd_sc_hd__ebufn_2
X_05500_ _05500_/A _05529_/Y vssd1 vssd1 vccd1 vccd1 _13620_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.M\[0\].MUX\[3\]_A0 _13634_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10300__D line[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06480_ _06480_/A _06509_/Y vssd1 vssd1 vccd1 vccd1 _13760_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_178_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05431_ _05455_/CLK line[108] vssd1 vssd1 vccd1 vccd1 _05432_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_60_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08150_ _08150_/CLK line[57] vssd1 vssd1 vccd1 vccd1 _08151_/A sky130_fd_sc_hd__dfxtp_1
X_05362_ _05362_/A _05389_/Y vssd1 vssd1 vccd1 vccd1 _13762_/Z sky130_fd_sc_hd__ebufn_2
X_07101_ _07101_/A _07104_/Y vssd1 vssd1 vccd1 vccd1 _13821_/Z sky130_fd_sc_hd__ebufn_2
X_08081_ _08081_/A _08084_/Y vssd1 vssd1 vccd1 vccd1 _13681_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12227__D line[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05293_ _05315_/CLK line[45] vssd1 vssd1 vccd1 vccd1 _05294_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[18\].VALID\[9\].TOBUF OVHB\[18\].VALID\[9\].FF/Q OVHB\[18\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04914_/B2 sky130_fd_sc_hd__ebufn_2
XOVHB\[24\].VALID\[4\].FF OVHB\[24\].V/CLK A[11] vssd1 vssd1 vccd1 vccd1 OVHB\[24\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_07032_ _07032_/CLK _07033_/X vssd1 vssd1 vccd1 vccd1 _07030_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__06225__D line[73] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09536__D line[50] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08983_ _08983_/A _08994_/Y vssd1 vssd1 vccd1 vccd1 _13743_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_69_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09833__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07934_ _07940_/CLK line[86] vssd1 vssd1 vccd1 vccd1 _07935_/A sky130_fd_sc_hd__dfxtp_1
X_07865_ _07865_/A _07874_/Y vssd1 vssd1 vccd1 vccd1 _13745_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_95_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09604_ _09620_/CLK line[81] vssd1 vssd1 vccd1 vccd1 _09605_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06895__D line[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06816_ _06820_/CLK line[87] vssd1 vssd1 vccd1 vccd1 _06817_/A sky130_fd_sc_hd__dfxtp_1
X_07796_ _07800_/CLK line[23] vssd1 vssd1 vccd1 vccd1 _07797_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_113_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06747_ _06747_/A _06754_/Y vssd1 vssd1 vccd1 vccd1 _13747_/Z sky130_fd_sc_hd__ebufn_2
X_09535_ _09535_/A _09554_/Y vssd1 vssd1 vccd1 vccd1 _13735_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[12\].CLKBUF\[5\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09466_ _09480_/CLK line[18] vssd1 vssd1 vccd1 vccd1 _09467_/A sky130_fd_sc_hd__dfxtp_1
XPHY_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06678_ _06680_/CLK line[24] vssd1 vssd1 vccd1 vccd1 _06679_/A sky130_fd_sc_hd__dfxtp_1
XPHY_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08417_ _08417_/A _08434_/Y vssd1 vssd1 vccd1 vccd1 _13737_/Z sky130_fd_sc_hd__ebufn_2
X_05629_ _05629_/A _05634_/Y vssd1 vssd1 vccd1 vccd1 _13749_/Z sky130_fd_sc_hd__ebufn_2
X_09397_ _09397_/A _09414_/Y vssd1 vssd1 vccd1 vccd1 _13877_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08348_ _08360_/CLK line[19] vssd1 vssd1 vccd1 vccd1 _08349_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08279_ _08279_/A _08294_/Y vssd1 vssd1 vccd1 vccd1 _13879_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11041__D line[98] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[8\].VALID\[4\].FF_D A[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10310_ _10320_/CLK line[20] vssd1 vssd1 vccd1 vccd1 _10311_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_22_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06135__D line[46] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11290_ _11300_/CLK line[84] vssd1 vssd1 vccd1 vccd1 _11291_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11976__D line[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10241_ _10241_/A _10254_/Y vssd1 vssd1 vccd1 vccd1 _13881_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10880__D line[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_DATA\[5\].CLKBUF\[5\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05974__D line[86] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08350__D line[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10172_ _10180_/CLK line[85] vssd1 vssd1 vccd1 vccd1 _10173_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_120_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[22\].VALID\[6\].FF OVHB\[22\].V/CLK A[13] vssd1 vssd1 vccd1 vccd1 OVHB\[22\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XOVHB\[24\].VALID\[8\].TOBUF OVHB\[24\].VALID\[8\].FF/Q OVHB\[24\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04931_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[31\].CLKBUF\[7\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13931_ _13938_/A _13938_/B _13938_/C _13938_/D vssd1 vssd1 vccd1 vccd1 _13931_/Y
+ sky130_fd_sc_hd__nor4b_4
XFILLER_208_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XOVHB\[30\].VALID\[11\].FF OVHB\[30\].V/CLK A[18] vssd1 vssd1 vccd1 vccd1 OVHB\[30\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[28\].V_RESET_B rst_n vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12600__D line[48] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13862_ _13890_/CLK line[122] vssd1 vssd1 vccd1 vccd1 _13863_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12813_ _12813_/A _12844_/Y vssd1 vssd1 vccd1 vccd1 _13653_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_28_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13793_ _13793_/A _13824_/Y vssd1 vssd1 vccd1 vccd1 _13793_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11216__D line[50] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12744_ _12770_/CLK line[123] vssd1 vssd1 vccd1 vccd1 _12745_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_188_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11513__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12675_ _12675_/A _12704_/Y vssd1 vssd1 vccd1 vccd1 _13795_/Z sky130_fd_sc_hd__ebufn_2
XPHY_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13431__D line[39] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08525__D line[100] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11626_ _11650_/CLK line[124] vssd1 vssd1 vccd1 vccd1 _11627_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11557_ _11557_/A _11584_/Y vssd1 vssd1 vccd1 vccd1 _13797_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10508_ _10530_/CLK line[125] vssd1 vssd1 vccd1 vccd1 _10509_/A sky130_fd_sc_hd__dfxtp_1
X_11488_ _11510_/CLK line[61] vssd1 vssd1 vccd1 vccd1 _11489_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_155_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10790__D line[126] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13227_ _13227_/CLK _13228_/X vssd1 vssd1 vccd1 vccd1 _13225_/CLK sky130_fd_sc_hd__dlclkp_1
XOVHB\[20\].VALID\[13\].FF OVHB\[20\].V/CLK A[20] vssd1 vssd1 vccd1 vccd1 OVHB\[20\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_10439_ _10439_/A _10464_/Y vssd1 vssd1 vccd1 vccd1 _13799_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05884__D line[59] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08260__D line[112] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13158_ _13938_/X wr vssd1 vssd1 vccd1 vccd1 _13158_/X sky130_fd_sc_hd__and2_1
X_12109_ _13934_/X vssd1 vssd1 vccd1 vccd1 _12109_/Y sky130_fd_sc_hd__inv_2
X_13089_ _13938_/X vssd1 vssd1 vccd1 vccd1 _13089_/Y sky130_fd_sc_hd__inv_2
X_05980_ _05980_/CLK line[89] vssd1 vssd1 vccd1 vccd1 _05981_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07454__A _13910_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_04931_ A_h[13] _04931_/B2 A_h[13] _04931_/B2 vssd1 vssd1 vccd1 vccd1 _04933_/C sky130_fd_sc_hd__a2bb2oi_2
XANTENNA_OVHB\[18\].VALID\[13\].FF_D A[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13606__D line[119] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07173__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07650_ _07660_/CLK line[84] vssd1 vssd1 vccd1 vccd1 _07651_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_81_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09091__D line[103] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06601_ _06601_/A _06614_/Y vssd1 vssd1 vccd1 vccd1 _13881_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_80_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07581_ _07581_/A _07594_/Y vssd1 vssd1 vccd1 vccd1 _13741_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[3\].VALID\[11\].TOBUF OVHB\[3\].VALID\[11\].FF/Q OVHB\[3\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04915_/B2 sky130_fd_sc_hd__ebufn_2
X_09320_ _09340_/CLK line[94] vssd1 vssd1 vccd1 vccd1 _09321_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[20\].VALID\[8\].FF OVHB\[20\].V/CLK A[15] vssd1 vssd1 vccd1 vccd1 OVHB\[20\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10030__D line[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06532_ _06540_/CLK line[85] vssd1 vssd1 vccd1 vccd1 _06533_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05124__D line[81] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09251_ _09251_/A _09274_/Y vssd1 vssd1 vccd1 vccd1 _13731_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[30\].VALID\[7\].TOBUF OVHB\[30\].VALID\[7\].FF/Q OVHB\[30\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/A2 sky130_fd_sc_hd__ebufn_2
X_06463_ _06463_/A _06474_/Y vssd1 vssd1 vccd1 vccd1 _13743_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10965__D line[78] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13341__D line[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08202_ _08220_/CLK line[95] vssd1 vssd1 vccd1 vccd1 _08203_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__04963__D line[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05414_ _05420_/CLK line[86] vssd1 vssd1 vccd1 vccd1 _05415_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_166_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09182_ _09200_/CLK line[31] vssd1 vssd1 vccd1 vccd1 _09183_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08435__D line[64] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06394_ _06400_/CLK line[22] vssd1 vssd1 vccd1 vccd1 _06395_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[28\].VALID\[12\].FF_D A[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[8\].VALID\[0\].TOBUF OVHB\[8\].VALID\[0\].FF/Q OVHB\[8\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04924_/B2 sky130_fd_sc_hd__ebufn_2
X_08133_ _08133_/A _08154_/Y vssd1 vssd1 vccd1 vccd1 _13733_/Z sky130_fd_sc_hd__ebufn_2
X_05345_ _05345_/A _05354_/Y vssd1 vssd1 vccd1 vccd1 _13745_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_146_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08064_ _08080_/CLK line[17] vssd1 vssd1 vccd1 vccd1 _08065_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07629__A _13911_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05276_ _05280_/CLK line[23] vssd1 vssd1 vccd1 vccd1 _05277_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_162_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07015_ _07015_/A _07034_/Y vssd1 vssd1 vccd1 vccd1 _13735_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07348__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09266__D line[55] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10205__D line[100] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08966_ _08990_/CLK line[60] vssd1 vssd1 vccd1 vccd1 _08967_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[17\].INV _13954_/X vssd1 vssd1 vccd1 vccd1 OVHB\[17\].INV/Y sky130_fd_sc_hd__inv_2
XFILLER_130_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07917_ _07917_/A _07944_/Y vssd1 vssd1 vccd1 vccd1 _13797_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_187_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08897_ _08897_/A _08924_/Y vssd1 vssd1 vccd1 vccd1 _13657_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13516__D line[92] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12420__D line[89] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07848_ _07870_/CLK line[61] vssd1 vssd1 vccd1 vccd1 _07849_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07514__D line[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XOVHB\[19\].VALID\[9\].FF OVHB\[19\].V/CLK A[16] vssd1 vssd1 vccd1 vccd1 OVHB\[19\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_07779_ _07779_/A _07804_/Y vssd1 vssd1 vccd1 vccd1 _13659_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_140_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09518_ _13920_/Y wr vssd1 vssd1 vccd1 vccd1 _09518_/X sky130_fd_sc_hd__and2_1
X_10790_ _10810_/CLK line[126] vssd1 vssd1 vccd1 vccd1 _10791_/A sky130_fd_sc_hd__dfxtp_1
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09449_ _13920_/Y vssd1 vssd1 vccd1 vccd1 _09449_/Y sky130_fd_sc_hd__inv_2
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12460_ _12490_/CLK line[112] vssd1 vssd1 vccd1 vccd1 _12461_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_12_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08923__A _13915_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_DATA\[10\].CLKBUF\[7\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11411_ _11411_/A _11444_/Y vssd1 vssd1 vccd1 vccd1 _13651_/Z sky130_fd_sc_hd__ebufn_2
X_12391_ _12391_/A _12424_/Y vssd1 vssd1 vccd1 vccd1 _13791_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_165_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11342_ _11370_/CLK line[122] vssd1 vssd1 vccd1 vccd1 _11343_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_165_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[30\].VALID\[8\].FF_D A[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11273_ _11273_/A _11304_/Y vssd1 vssd1 vccd1 vccd1 _13793_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09176__D line[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10224_ _10250_/CLK line[123] vssd1 vssd1 vccd1 vccd1 _10225_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08080__D line[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MUX.M\[2\].MUX\[4\]_A2 _13811_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13012_ _13012_/A _13019_/Y vssd1 vssd1 vccd1 vccd1 _13852_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10115__D line[64] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10155_ _10155_/A _10184_/Y vssd1 vssd1 vccd1 vccd1 _13795_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_79_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10086_ _10110_/CLK line[60] vssd1 vssd1 vccd1 vccd1 _10087_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[3\].CLKBUF\[7\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12330__D line[62] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13914_ _13916_/B _13916_/A _13916_/C _13916_/D vssd1 vssd1 vccd1 vccd1 _13914_/X
+ sky130_fd_sc_hd__and4b_4
XANTENNA__07424__D line[123] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13845_ _13855_/CLK line[100] vssd1 vssd1 vccd1 vccd1 _13846_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_16_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XOVHB\[10\].CG clk OVHB\[10\].CGAND/X vssd1 vssd1 vccd1 vccd1 OVHB\[10\].V/CLK sky130_fd_sc_hd__dlclkp_1
X_13776_ _13776_/A _13789_/Y vssd1 vssd1 vccd1 vccd1 _13776_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_200_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10988_ _13925_/X wr vssd1 vssd1 vccd1 vccd1 _10988_/X sky130_fd_sc_hd__and2_1
XFILLER_203_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12727_ _12735_/CLK line[101] vssd1 vssd1 vccd1 vccd1 _12728_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_30_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_MUX.M\[0\].MUX\[0\]_A3 _13826_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[26\].VALID\[13\].TOBUF OVHB\[26\].VALID\[13\].FF/Q OVHB\[26\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04916_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_188_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08255__D line[105] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12658_ _12658_/A _12669_/Y vssd1 vssd1 vccd1 vccd1 _13778_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11609_ _11615_/CLK line[102] vssd1 vssd1 vccd1 vccd1 _11610_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12589_ _12595_/CLK line[38] vssd1 vssd1 vccd1 vccd1 _12590_/A sky130_fd_sc_hd__dfxtp_1
X_05130_ _05140_/CLK line[84] vssd1 vssd1 vccd1 vccd1 _05131_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[13\].VALID\[0\].FF_D A[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12505__D line[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05061_ _05061_/A _05074_/Y vssd1 vssd1 vccd1 vccd1 _13741_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06503__D line[72] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08820_ _08850_/CLK line[112] vssd1 vssd1 vccd1 vccd1 _08821_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10603__A _13924_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09814__D line[49] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08751_ _08751_/A _08784_/Y vssd1 vssd1 vccd1 vccd1 _13791_/Z sky130_fd_sc_hd__ebufn_2
X_05963_ _05963_/A _05984_/Y vssd1 vssd1 vccd1 vccd1 _13803_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_100_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XOVHB\[6\].VALID\[5\].TOBUF OVHB\[6\].VALID\[5\].FF/Q OVHB\[6\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04927_/B2 sky130_fd_sc_hd__ebufn_2
X_04914_ _04913_/Y _04922_/A2 _04911_/Y _04914_/B2 vssd1 vssd1 vccd1 vccd1 _04917_/B
+ sky130_fd_sc_hd__a22o_2
XFILLER_66_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07702_ _07730_/CLK line[122] vssd1 vssd1 vccd1 vccd1 _07703_/A sky130_fd_sc_hd__dfxtp_1
X_08682_ _08710_/CLK line[58] vssd1 vssd1 vccd1 vccd1 _08683_/A sky130_fd_sc_hd__dfxtp_1
X_05894_ _05910_/CLK line[49] vssd1 vssd1 vccd1 vccd1 _05895_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_54_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07633_ _07633_/A _07664_/Y vssd1 vssd1 vccd1 vccd1 _13793_/Z sky130_fd_sc_hd__ebufn_2
X_07564_ _07590_/CLK line[59] vssd1 vssd1 vccd1 vccd1 _07565_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_53_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09303_ _09305_/CLK line[72] vssd1 vssd1 vccd1 vccd1 _09304_/A sky130_fd_sc_hd__dfxtp_1
X_06515_ _06515_/A _06544_/Y vssd1 vssd1 vccd1 vccd1 _13795_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10695__D line[68] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07495_ _07495_/A _07524_/Y vssd1 vssd1 vccd1 vccd1 _13655_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13071__D line[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05789__D line[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06446_ _06470_/CLK line[60] vssd1 vssd1 vccd1 vccd1 _06447_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08165__D line[78] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09234_ _09234_/A _09239_/Y vssd1 vssd1 vccd1 vccd1 _13714_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[4\].VALID\[7\].FF_D A[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09165_ _09165_/CLK line[9] vssd1 vssd1 vccd1 vccd1 _09166_/A sky130_fd_sc_hd__dfxtp_1
X_06377_ _06377_/A _06404_/Y vssd1 vssd1 vccd1 vccd1 _13657_/Z sky130_fd_sc_hd__ebufn_2
X_08116_ _08116_/A _08119_/Y vssd1 vssd1 vccd1 vccd1 _13716_/Z sky130_fd_sc_hd__ebufn_2
X_05328_ _05350_/CLK line[61] vssd1 vssd1 vccd1 vccd1 _05329_/A sky130_fd_sc_hd__dfxtp_1
X_09096_ _09096_/A _09099_/Y vssd1 vssd1 vccd1 vccd1 _13856_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06263__A _13903_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08047_ _08047_/CLK _08048_/X vssd1 vssd1 vccd1 vccd1 _08045_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_79_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05259_ _05259_/A _05284_/Y vssd1 vssd1 vccd1 vccd1 _13659_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_135_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06413__D line[45] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09998_ _09998_/A _10009_/Y vssd1 vssd1 vccd1 vccd1 _13638_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05029__D line[38] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08949_ _08955_/CLK line[38] vssd1 vssd1 vccd1 vccd1 _08950_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_151_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13246__D line[82] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13824__A _13899_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11960_ _11960_/A _11969_/Y vssd1 vssd1 vccd1 vccd1 _13640_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_72_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10911_ _10915_/CLK line[39] vssd1 vssd1 vccd1 vccd1 _10912_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13543__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11891_ _11895_/CLK line[103] vssd1 vssd1 vccd1 vccd1 _11892_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_17_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13630_ _13630_/A _13649_/Y vssd1 vssd1 vccd1 vccd1 _13630_/Z sky130_fd_sc_hd__ebufn_2
X_10842_ _10842_/A _10849_/Y vssd1 vssd1 vccd1 vccd1 _13642_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_198_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06438__A _13904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13561_ _13575_/CLK line[98] vssd1 vssd1 vccd1 vccd1 _13562_/A sky130_fd_sc_hd__dfxtp_1
X_10773_ _10775_/CLK line[104] vssd1 vssd1 vccd1 vccd1 _10774_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[5\].CG clk OVHB\[5\].CGAND/X vssd1 vssd1 vccd1 vccd1 OVHB\[5\].V/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA_DATA\[24\].CLKBUF\[1\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[13\].VALID\[0\].TOBUF OVHB\[13\].VALID\[0\].FF/Q OVHB\[13\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04924_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_40_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12512_ _12512_/A _12529_/Y vssd1 vssd1 vccd1 vccd1 _13632_/Z sky130_fd_sc_hd__ebufn_2
X_13492_ _13492_/A _13509_/Y vssd1 vssd1 vccd1 vccd1 _13772_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_100_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_OVHB\[26\].VALID\[0\].FF_D A[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12443_ _12455_/CLK line[99] vssd1 vssd1 vccd1 vccd1 _12444_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_176_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_200_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08803__D line[99] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12374_ _12374_/A _12389_/Y vssd1 vssd1 vccd1 vccd1 _13774_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_138_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11325_ _11335_/CLK line[100] vssd1 vssd1 vccd1 vccd1 _11326_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_5_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09484__A _13920_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11256_ _11256_/A _11269_/Y vssd1 vssd1 vccd1 vccd1 _13776_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[19\].VALID\[4\].FF_D A[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13718__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10207_ _10215_/CLK line[101] vssd1 vssd1 vccd1 vccd1 _10208_/A sky130_fd_sc_hd__dfxtp_1
X_11187_ _11195_/CLK line[37] vssd1 vssd1 vccd1 vccd1 _11188_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10138_ _10138_/A _10149_/Y vssd1 vssd1 vccd1 vccd1 _13778_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.M\[1\].MUX\[5\]_A0 _13624_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12060__D line[52] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10069_ _10075_/CLK line[38] vssd1 vssd1 vccd1 vccd1 _10070_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_63_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07154__D line[113] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12995__D line[110] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06993__D line[40] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13828_ _13828_/A _13859_/Y vssd1 vssd1 vccd1 vccd1 _13828_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_189_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13759_ _13785_/CLK line[75] vssd1 vssd1 vccd1 vccd1 _13760_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06300_ _06330_/CLK line[112] vssd1 vssd1 vccd1 vccd1 _06301_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09659__A _13920_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07280_ _07310_/CLK line[48] vssd1 vssd1 vccd1 vccd1 _07281_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05402__D line[95] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06231_ _06231_/A _06264_/Y vssd1 vssd1 vccd1 vccd1 _13791_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09378__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06162_ _06190_/CLK line[58] vssd1 vssd1 vccd1 vccd1 _06163_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_163_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[15\].VOBUF OVHB\[15\].V/Q OVHB\[15\].INV/Y vssd1 vssd1 vccd1 vccd1 _04912_/B1
+ sky130_fd_sc_hd__ebufn_2
XFILLER_144_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_OVHB\[13\].CGAND_A _13903_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDATA\[19\].CLKBUF\[4\] clk vssd1 vssd1 vccd1 vccd1 _07907_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_117_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05113_ _05113_/A _05144_/Y vssd1 vssd1 vccd1 vccd1 _13793_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12235__D line[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06093_ _06093_/A _06124_/Y vssd1 vssd1 vccd1 vccd1 _13653_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_117_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07329__D line[65] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05044_ _05070_/CLK line[59] vssd1 vssd1 vccd1 vccd1 _05045_/A sky130_fd_sc_hd__dfxtp_1
X_09921_ _09935_/CLK line[98] vssd1 vssd1 vccd1 vccd1 _09922_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_98_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09852_ _09852_/A _09869_/Y vssd1 vssd1 vccd1 vccd1 _13772_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_86_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09544__D line[54] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08803_ _08815_/CLK line[99] vssd1 vssd1 vccd1 vccd1 _08804_/A sky130_fd_sc_hd__dfxtp_1
X_09783_ _09795_/CLK line[35] vssd1 vssd1 vccd1 vccd1 _09784_/A sky130_fd_sc_hd__dfxtp_1
X_06995_ _06995_/CLK line[41] vssd1 vssd1 vccd1 vccd1 _06996_/A sky130_fd_sc_hd__dfxtp_1
X_08734_ _08734_/A _08749_/Y vssd1 vssd1 vccd1 vccd1 _13774_/Z sky130_fd_sc_hd__ebufn_2
X_05946_ _05946_/A _05949_/Y vssd1 vssd1 vccd1 vccd1 _13786_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_66_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05877_ _05877_/CLK _05878_/X vssd1 vssd1 vccd1 vccd1 _05875_/CLK sky130_fd_sc_hd__dlclkp_1
X_08665_ _08675_/CLK line[36] vssd1 vssd1 vccd1 vccd1 _08666_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11164__A _13933_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07616_ _07616_/A _07629_/Y vssd1 vssd1 vccd1 vccd1 _13776_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_42_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08596_ _08596_/A _08609_/Y vssd1 vssd1 vccd1 vccd1 _13636_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_202_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07547_ _07555_/CLK line[37] vssd1 vssd1 vccd1 vccd1 _07548_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07478_ _07478_/A _07489_/Y vssd1 vssd1 vccd1 vccd1 _13638_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_10_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09217_ _09235_/CLK line[47] vssd1 vssd1 vccd1 vccd1 _09218_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_210_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06429_ _06435_/CLK line[38] vssd1 vssd1 vccd1 vccd1 _06430_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09719__D line[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09148_ _09148_/A _09169_/Y vssd1 vssd1 vccd1 vccd1 _13628_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_107_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12145__D line[96] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09079_ _09095_/CLK line[97] vssd1 vssd1 vccd1 vccd1 _09080_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_30_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11110_ _11110_/A _11129_/Y vssd1 vssd1 vccd1 vccd1 _13630_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_30_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06143__D line[35] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12090_ _12090_/A _12109_/Y vssd1 vssd1 vccd1 vccd1 _13770_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11984__D line[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11339__A _13933_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11041_ _11055_/CLK line[98] vssd1 vssd1 vccd1 vccd1 _11042_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[8\].VALID\[6\].FF OVHB\[8\].V/CLK A[13] vssd1 vssd1 vccd1 vccd1 OVHB\[8\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XDATA\[18\].CLKBUF\[1\] clk vssd1 vssd1 vccd1 vccd1 _07522_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_77_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09454__D line[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XOVHB\[11\].VALID\[5\].TOBUF OVHB\[11\].VALID\[5\].FF/Q OVHB\[11\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04927_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__11058__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12992_ _12992_/A _13019_/Y vssd1 vssd1 vccd1 vccd1 _13832_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_17_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11943_ _11965_/CLK line[13] vssd1 vssd1 vccd1 vccd1 _11944_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_84_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11874_ _11874_/A _11899_/Y vssd1 vssd1 vccd1 vccd1 _13834_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_32_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07702__D line[122] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13613_ _13898_/Y wr vssd1 vssd1 vccd1 vccd1 _13613_/X sky130_fd_sc_hd__and2_1
X_10825_ _10845_/CLK line[14] vssd1 vssd1 vccd1 vccd1 _10826_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11224__D line[54] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06318__D line[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13544_ _13898_/Y vssd1 vssd1 vccd1 vccd1 _13544_/Y sky130_fd_sc_hd__inv_2
X_10756_ _10756_/A _10779_/Y vssd1 vssd1 vccd1 vccd1 _13836_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[25\].VALID\[13\].FF OVHB\[25\].V/CLK A[20] vssd1 vssd1 vccd1 vccd1 OVHB\[25\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_185_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13475_ _13505_/CLK line[64] vssd1 vssd1 vccd1 vccd1 _13476_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_173_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10687_ _10705_/CLK line[79] vssd1 vssd1 vccd1 vccd1 _10688_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_145_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09629__D line[107] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08533__D line[104] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12426_ _12426_/A _12459_/Y vssd1 vssd1 vccd1 vccd1 _13826_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[22\].CLKBUF\[3\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12357_ _12385_/CLK line[74] vssd1 vssd1 vccd1 vccd1 _12358_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12633__A _13936_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11308_ _11308_/A _11339_/Y vssd1 vssd1 vccd1 vccd1 _13828_/Z sky130_fd_sc_hd__ebufn_2
X_12288_ _12288_/A _12319_/Y vssd1 vssd1 vccd1 vccd1 _13688_/Z sky130_fd_sc_hd__ebufn_2
X_11239_ _11265_/CLK line[75] vssd1 vssd1 vccd1 vccd1 _11240_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05892__D line[63] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05800_ _05800_/A _05809_/Y vssd1 vssd1 vccd1 vccd1 _13640_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_95_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06780_ _06780_/A _06789_/Y vssd1 vssd1 vccd1 vccd1 _13780_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_209_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05731_ _05735_/CLK line[103] vssd1 vssd1 vccd1 vccd1 _05732_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[6\].VALID\[8\].FF OVHB\[6\].V/CLK A[15] vssd1 vssd1 vccd1 vccd1 OVHB\[6\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_75_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08450_ _08450_/A _08469_/Y vssd1 vssd1 vccd1 vccd1 _13770_/Z sky130_fd_sc_hd__ebufn_2
X_05662_ _05662_/A _05669_/Y vssd1 vssd1 vccd1 vccd1 _13782_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_24_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08708__D line[56] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07401_ _07415_/CLK line[98] vssd1 vssd1 vccd1 vccd1 _07402_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_196_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08381_ _08395_/CLK line[34] vssd1 vssd1 vccd1 vccd1 _08382_/A sky130_fd_sc_hd__dfxtp_1
X_05593_ _05595_/CLK line[40] vssd1 vssd1 vccd1 vccd1 _05594_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[16\].VALID\[11\].TOBUF OVHB\[16\].VALID\[11\].FF/Q OVHB\[16\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04915_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__12808__A _13937_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11134__D line[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07332_ _07332_/A _07349_/Y vssd1 vssd1 vccd1 vccd1 _13772_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_176_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05132__D line[85] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08293__A _13932_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10973__D line[67] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07263_ _07275_/CLK line[35] vssd1 vssd1 vccd1 vccd1 _07264_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_176_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06214_ _06214_/A _06229_/Y vssd1 vssd1 vccd1 vccd1 _13774_/Z sky130_fd_sc_hd__ebufn_2
X_09002_ _09002_/A _09029_/Y vssd1 vssd1 vccd1 vccd1 _13762_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08443__D line[77] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07194_ _07194_/A _07209_/Y vssd1 vssd1 vccd1 vccd1 _13634_/Z sky130_fd_sc_hd__ebufn_2
X_06145_ _06155_/CLK line[36] vssd1 vssd1 vccd1 vccd1 _06146_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_145_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07059__D line[70] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06076_ _06076_/A _06089_/Y vssd1 vssd1 vccd1 vccd1 _13636_/Z sky130_fd_sc_hd__ebufn_2
X_09904_ _13921_/X vssd1 vssd1 vccd1 vccd1 _09904_/Y sky130_fd_sc_hd__inv_2
X_05027_ _05035_/CLK line[37] vssd1 vssd1 vccd1 vccd1 _05028_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_113_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09835_ _09865_/CLK line[64] vssd1 vssd1 vccd1 vccd1 _09836_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11309__D line[107] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10213__D line[104] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09766_ _09766_/A _09799_/Y vssd1 vssd1 vccd1 vccd1 _13686_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08468__A _13913_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06978_ _06978_/A _06999_/Y vssd1 vssd1 vccd1 vccd1 _13698_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05307__D line[37] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08717_ _08745_/CLK line[74] vssd1 vssd1 vccd1 vccd1 _08718_/A sky130_fd_sc_hd__dfxtp_1
X_05929_ _05945_/CLK line[65] vssd1 vssd1 vccd1 vccd1 _05930_/A sky130_fd_sc_hd__dfxtp_1
X_09697_ _09725_/CLK line[10] vssd1 vssd1 vccd1 vccd1 _09698_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_199_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13524__D line[81] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_199_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08618__D line[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08648_ _08648_/A _08679_/Y vssd1 vssd1 vccd1 vccd1 _13688_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08579_ _08605_/CLK line[11] vssd1 vssd1 vccd1 vccd1 _08580_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[22\].VALID\[3\].FF_D A[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10610_ _10610_/A _10639_/Y vssd1 vssd1 vccd1 vccd1 _13690_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05042__D line[58] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11590_ _11590_/A _11619_/Y vssd1 vssd1 vccd1 vccd1 _13830_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10541_ _10565_/CLK line[12] vssd1 vssd1 vccd1 vccd1 _10542_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MUX.M\[3\].MUX\[6\]_A2 _13801_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13260_ _13260_/CLK line[89] vssd1 vssd1 vccd1 vccd1 _13261_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_210_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10472_ _10472_/A _10499_/Y vssd1 vssd1 vccd1 vccd1 _13832_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_182_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12211_ _12211_/A _12214_/Y vssd1 vssd1 vccd1 vccd1 _13891_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[15\].VALID\[7\].FF_D A[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13191_ _13191_/A _13194_/Y vssd1 vssd1 vccd1 vccd1 _13751_/Z sky130_fd_sc_hd__ebufn_2
X_12142_ _12142_/CLK _12143_/X vssd1 vssd1 vccd1 vccd1 _12140_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_123_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12073_ _13934_/X wr vssd1 vssd1 vccd1 vccd1 _12073_/X sky130_fd_sc_hd__and2_1
XFILLER_151_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09184__D line[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11024_ _13925_/X vssd1 vssd1 vccd1 vccd1 _11024_/Y sky130_fd_sc_hd__inv_2
XANTENNA__10123__D line[77] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05217__D line[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_MUX.M\[1\].MUX\[2\]_A3 _13828_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12975_ _12975_/A _12984_/Y vssd1 vssd1 vccd1 vccd1 _13815_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_205_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11926_ _11930_/CLK line[119] vssd1 vssd1 vccd1 vccd1 _11927_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_206_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_OVHB\[8\].CG_CLK clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07432__D line[127] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[15\].VALID\[0\].FF OVHB\[15\].V/CLK A[7] vssd1 vssd1 vccd1 vccd1 OVHB\[15\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_11857_ _11857_/A _11864_/Y vssd1 vssd1 vccd1 vccd1 _13817_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_32_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10808_ _10810_/CLK line[120] vssd1 vssd1 vccd1 vccd1 _10809_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06048__D line[120] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11788_ _11790_/CLK line[56] vssd1 vssd1 vccd1 vccd1 _11789_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11889__D line[102] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13527_ _13527_/A _13544_/Y vssd1 vssd1 vccd1 vccd1 _13807_/Z sky130_fd_sc_hd__ebufn_2
X_10739_ _10739_/A _10744_/Y vssd1 vssd1 vccd1 vccd1 _13819_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10148__A _13922_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09359__D line[97] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13458_ _13470_/CLK line[51] vssd1 vssd1 vccd1 vccd1 _13459_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_146_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[23\].CGAND _13916_/X wr vssd1 vssd1 vccd1 vccd1 OVHB\[23\].CGAND/X sky130_fd_sc_hd__and2_4
X_12409_ _12409_/A _12424_/Y vssd1 vssd1 vccd1 vccd1 _13809_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[5\].VALID\[12\].FF_D A[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13389_ _13389_/A _13404_/Y vssd1 vssd1 vccd1 vccd1 _13669_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12513__D line[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07950_ _07950_/A _07979_/Y vssd1 vssd1 vccd1 vccd1 _13830_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07607__D line[79] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06901_ _06925_/CLK line[12] vssd1 vssd1 vccd1 vccd1 _06902_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[20\].CLKBUF\[5\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07881_ _07905_/CLK line[76] vssd1 vssd1 vccd1 vccd1 _07882_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_95_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09620_ _09620_/CLK line[89] vssd1 vssd1 vccd1 vccd1 _09621_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13194__A _13938_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06832_ _06832_/A _06859_/Y vssd1 vssd1 vccd1 vccd1 _13832_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09822__D line[53] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09551_ _09551_/A _09554_/Y vssd1 vssd1 vccd1 vccd1 _13751_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[18\].VALID\[5\].TOBUF OVHB\[18\].VALID\[5\].FF/Q OVHB\[18\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04927_/B2 sky130_fd_sc_hd__ebufn_2
X_06763_ _06785_/CLK line[77] vssd1 vssd1 vccd1 vccd1 _06764_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_48_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XOVHB\[21\].VALID\[11\].FF OVHB\[21\].V/CLK A[18] vssd1 vssd1 vccd1 vccd1 OVHB\[21\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_08502_ _08502_/CLK _08503_/X vssd1 vssd1 vccd1 vccd1 _08500_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05714_ _05714_/A _05739_/Y vssd1 vssd1 vccd1 vccd1 _13834_/Z sky130_fd_sc_hd__ebufn_2
X_09482_ _09482_/CLK _09483_/X vssd1 vssd1 vccd1 vccd1 _09480_/CLK sky130_fd_sc_hd__dlclkp_1
X_06694_ _06694_/A _06719_/Y vssd1 vssd1 vccd1 vccd1 _13694_/Z sky130_fd_sc_hd__ebufn_2
XPHY_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08433_ _13913_/X wr vssd1 vssd1 vccd1 vccd1 _08433_/X sky130_fd_sc_hd__and2_1
X_05645_ _05665_/CLK line[78] vssd1 vssd1 vccd1 vccd1 _05646_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08364_ _13913_/X vssd1 vssd1 vccd1 vccd1 _08364_/Y sky130_fd_sc_hd__inv_2
XPHY_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05576_ _05576_/A _05599_/Y vssd1 vssd1 vccd1 vccd1 _13696_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11799__D line[75] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07315_ _07345_/CLK line[64] vssd1 vssd1 vccd1 vccd1 _07316_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_149_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08295_ _08325_/CLK line[0] vssd1 vssd1 vccd1 vccd1 _08296_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05797__D line[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[28\].VALID\[7\].FF_D A[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08173__D line[67] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07246_ _07246_/A _07279_/Y vssd1 vssd1 vccd1 vccd1 _13686_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[13\].VALID\[2\].FF OVHB\[13\].V/CLK A[9] vssd1 vssd1 vccd1 vccd1 OVHB\[13\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13369__A _13898_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07177_ _07205_/CLK line[10] vssd1 vssd1 vccd1 vccd1 _07178_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_180_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XOVHB\[30\].VALID\[6\].FF OVHB\[30\].V/CLK A[13] vssd1 vssd1 vccd1 vccd1 OVHB\[30\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_06128_ _06128_/A _06159_/Y vssd1 vssd1 vccd1 vccd1 _13688_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13088__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06059_ _06085_/CLK line[11] vssd1 vssd1 vccd1 vccd1 _06060_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[11\].VALID\[13\].FF OVHB\[11\].V/CLK A[20] vssd1 vssd1 vccd1 vccd1 OVHB\[11\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_160_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06421__D line[34] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_OVHB\[27\].V_RESET_B rst_n vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11039__D line[97] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09818_ _09830_/CLK line[51] vssd1 vssd1 vccd1 vccd1 _09819_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09732__D line[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10878__D line[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09749_ _09749_/A _09764_/Y vssd1 vssd1 vccd1 vccd1 _13669_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13254__D line[86] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08348__D line[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12760_ _12770_/CLK line[116] vssd1 vssd1 vccd1 vccd1 _12761_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_160_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ _11711_/A _11724_/Y vssd1 vssd1 vccd1 vccd1 _13671_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12691_ _12691_/A _12704_/Y vssd1 vssd1 vccd1 vccd1 _13811_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_14_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11642_ _11650_/CLK line[117] vssd1 vssd1 vccd1 vccd1 _11643_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11573_ _11573_/A _11584_/Y vssd1 vssd1 vccd1 vccd1 _13813_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[24\].VALID\[4\].TOBUF OVHB\[24\].VALID\[4\].FF/Q OVHB\[24\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04925_/B2 sky130_fd_sc_hd__ebufn_2
XPHY_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11502__D line[53] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13312_ _13330_/CLK line[127] vssd1 vssd1 vccd1 vccd1 _13313_/A sky130_fd_sc_hd__dfxtp_1
X_10524_ _10530_/CLK line[118] vssd1 vssd1 vccd1 vccd1 _10525_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[29\].VALID\[7\].FF OVHB\[29\].V/CLK A[14] vssd1 vssd1 vccd1 vccd1 OVHB\[29\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_13243_ _13243_/A _13264_/Y vssd1 vssd1 vccd1 vccd1 _13803_/Z sky130_fd_sc_hd__ebufn_2
X_10455_ _10455_/A _10464_/Y vssd1 vssd1 vccd1 vccd1 _13815_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.M\[2\].MUX\[7\]_A0 _13677_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09907__D line[106] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08811__D line[103] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13174_ _13190_/CLK line[49] vssd1 vssd1 vccd1 vccd1 _13175_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[9\].CLKBUF\[5\] clk vssd1 vssd1 vccd1 vccd1 _13822_/CLK sky130_fd_sc_hd__clkbuf_4
X_10386_ _10390_/CLK line[55] vssd1 vssd1 vccd1 vccd1 _10387_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13429__D line[38] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12125_ _12125_/A _12144_/Y vssd1 vssd1 vccd1 vccd1 _13805_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[19\].CLKBUF\[6\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XOVHB\[11\].VALID\[4\].FF OVHB\[11\].V/CLK A[11] vssd1 vssd1 vccd1 vccd1 OVHB\[11\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_12056_ _12070_/CLK line[50] vssd1 vssd1 vccd1 vccd1 _12057_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[9\].VALID\[2\].FF_D A[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11007_ _11007_/A _11024_/Y vssd1 vssd1 vccd1 vccd1 _13807_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_65_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10788__D line[125] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13164__D line[59] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12958_ _12980_/CLK line[93] vssd1 vssd1 vccd1 vccd1 _12959_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07162__D line[117] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11909_ _11909_/A _11934_/Y vssd1 vssd1 vccd1 vccd1 _13869_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.M\[0\].MUX\[3\]_A1 _13704_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12889_ _12889_/A _12914_/Y vssd1 vssd1 vccd1 vccd1 _13729_/Z sky130_fd_sc_hd__ebufn_2
X_05430_ _05430_/A _05459_/Y vssd1 vssd1 vccd1 vccd1 _13830_/Z sky130_fd_sc_hd__ebufn_2
X_05361_ _05385_/CLK line[76] vssd1 vssd1 vccd1 vccd1 _05362_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_174_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11412__D line[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09089__D line[102] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07100_ _07100_/CLK line[89] vssd1 vssd1 vccd1 vccd1 _07101_/A sky130_fd_sc_hd__dfxtp_1
X_08080_ _08080_/CLK line[25] vssd1 vssd1 vccd1 vccd1 _08081_/A sky130_fd_sc_hd__dfxtp_1
X_05292_ _05292_/A _05319_/Y vssd1 vssd1 vccd1 vccd1 _13692_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05410__D line[84] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07031_ _07031_/A _07034_/Y vssd1 vssd1 vccd1 vccd1 _13751_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10028__D line[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08721__D line[76] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13339__D line[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12243__D line[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13917__A A[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08982_ _08990_/CLK line[53] vssd1 vssd1 vccd1 vccd1 _08983_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07337__D line[69] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[30\].VALID\[3\].TOBUF OVHB\[30\].VALID\[3\].FF/Q OVHB\[30\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04919_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_130_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XOVHB\[27\].VALID\[9\].FF OVHB\[27\].V/CLK A[16] vssd1 vssd1 vccd1 vccd1 OVHB\[27\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_87_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07933_ _07933_/A _07944_/Y vssd1 vssd1 vccd1 vccd1 _13813_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[8\].CLKBUF\[2\] clk vssd1 vssd1 vccd1 vccd1 _13437_/CLK sky130_fd_sc_hd__clkbuf_4
X_07864_ _07870_/CLK line[54] vssd1 vssd1 vccd1 vccd1 _07865_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_113_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09603_ _09603_/A _09624_/Y vssd1 vssd1 vccd1 vccd1 _13803_/Z sky130_fd_sc_hd__ebufn_2
X_06815_ _06815_/A _06824_/Y vssd1 vssd1 vccd1 vccd1 _13815_/Z sky130_fd_sc_hd__ebufn_2
X_07795_ _07795_/A _07804_/Y vssd1 vssd1 vccd1 vccd1 _13675_/Z sky130_fd_sc_hd__ebufn_2
X_09534_ _09550_/CLK line[49] vssd1 vssd1 vccd1 vccd1 _09535_/A sky130_fd_sc_hd__dfxtp_1
X_06746_ _06750_/CLK line[55] vssd1 vssd1 vccd1 vccd1 _06747_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07072__D line[90] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09465_ _09465_/A _09484_/Y vssd1 vssd1 vccd1 vccd1 _13665_/Z sky130_fd_sc_hd__ebufn_2
XPHY_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06677_ _06677_/A _06684_/Y vssd1 vssd1 vccd1 vccd1 _13677_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13802__D line[95] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08416_ _08430_/CLK line[50] vssd1 vssd1 vccd1 vccd1 _08417_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05628_ _05630_/CLK line[56] vssd1 vssd1 vccd1 vccd1 _05629_/A sky130_fd_sc_hd__dfxtp_1
X_09396_ _09410_/CLK line[114] vssd1 vssd1 vccd1 vccd1 _09397_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07800__D line[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08347_ _08347_/A _08364_/Y vssd1 vssd1 vccd1 vccd1 _13667_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12418__D line[88] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05559_ _05559_/A _05564_/Y vssd1 vssd1 vccd1 vccd1 _13679_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05320__D line[48] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08278_ _08290_/CLK line[115] vssd1 vssd1 vccd1 vccd1 _08279_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_22_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07229_ _07229_/A _07244_/Y vssd1 vssd1 vccd1 vccd1 _13669_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XDATA\[28\].CLKBUF\[6\] clk vssd1 vssd1 vccd1 vccd1 _10777_/CLK sky130_fd_sc_hd__clkbuf_4
X_10240_ _10250_/CLK line[116] vssd1 vssd1 vccd1 vccd1 _10241_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12153__D line[109] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10171_ _10171_/A _10184_/Y vssd1 vssd1 vccd1 vccd1 _13811_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07247__D line[42] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06151__D line[39] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11992__D line[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13930_ A[4] vssd1 vssd1 vccd1 vccd1 _13938_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_47_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09462__D line[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[22\].VALID\[9\].TOBUF OVHB\[22\].VALID\[9\].FF/Q OVHB\[22\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04914_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_207_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13861_ _13861_/A _13894_/Y vssd1 vssd1 vccd1 vccd1 _13861_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_207_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12812_ _12840_/CLK line[26] vssd1 vssd1 vccd1 vccd1 _12813_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10401__D line[76] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08078__D line[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13792_ _13820_/CLK line[90] vssd1 vssd1 vccd1 vccd1 _13793_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_55_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XOVHB\[6\].VALID\[13\].TOBUF OVHB\[6\].VALID\[13\].FF/Q OVHB\[6\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04916_/B2 sky130_fd_sc_hd__ebufn_2
X_12743_ _12743_/A _12774_/Y vssd1 vssd1 vccd1 vccd1 _13863_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12178__A _13934_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12674_ _12700_/CLK line[91] vssd1 vssd1 vccd1 vccd1 _12675_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_43_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07710__D line[126] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11625_ _11625_/A _11654_/Y vssd1 vssd1 vccd1 vccd1 _13865_/Z sky130_fd_sc_hd__ebufn_2
XPHY_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12328__D line[61] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06326__D line[119] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11556_ _11580_/CLK line[92] vssd1 vssd1 vccd1 vccd1 _11557_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_11_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10507_ _10507_/A _10534_/Y vssd1 vssd1 vccd1 vccd1 _13867_/Z sky130_fd_sc_hd__ebufn_2
X_11487_ _11487_/A _11514_/Y vssd1 vssd1 vccd1 vccd1 _13727_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_195_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09637__D line[111] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13226_ _13226_/A _13229_/Y vssd1 vssd1 vccd1 vccd1 _13786_/Z sky130_fd_sc_hd__ebufn_2
X_10438_ _10460_/CLK line[93] vssd1 vssd1 vccd1 vccd1 _10439_/A sky130_fd_sc_hd__dfxtp_1
X_13157_ _13157_/CLK _13158_/X vssd1 vssd1 vccd1 vccd1 _13155_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_112_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10369_ _10369_/A _10394_/Y vssd1 vssd1 vccd1 vccd1 _13729_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06061__D line[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12108_ _13934_/X wr vssd1 vssd1 vccd1 vccd1 _12108_/X sky130_fd_sc_hd__and2_1
X_13088_ _13938_/X wr vssd1 vssd1 vccd1 vccd1 _13088_/X sky130_fd_sc_hd__and2_1
XFILLER_85_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XDATA\[27\].CLKBUF\[3\] clk vssd1 vssd1 vccd1 vccd1 _10392_/CLK sky130_fd_sc_hd__clkbuf_4
XMUX.M\[3\].MUX\[4\] _13657_/Z _13727_/Z _13797_/Z _13867_/Z MUX.SEL0BUF\[3\]/X MUX.SEL1BUF\[3\]/X
+ vssd1 vssd1 vccd1 vccd1 Do[28] sky130_fd_sc_hd__mux4_1
X_04930_ A_h[7] _04930_/B2 A_h[7] _04930_/B2 vssd1 vssd1 vccd1 vccd1 _04933_/B sky130_fd_sc_hd__a2bb2oi_2
X_12039_ _13934_/X vssd1 vssd1 vccd1 vccd1 _12039_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[31\].VALID\[6\].FF_D A[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06600_ _06610_/CLK line[116] vssd1 vssd1 vccd1 vccd1 _06601_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_92_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07580_ _07590_/CLK line[52] vssd1 vssd1 vccd1 vccd1 _07581_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_179_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06531_ _06531_/A _06544_/Y vssd1 vssd1 vccd1 vccd1 _13811_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_179_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09250_ _09270_/CLK line[62] vssd1 vssd1 vccd1 vccd1 _09251_/A sky130_fd_sc_hd__dfxtp_1
X_06462_ _06470_/CLK line[53] vssd1 vssd1 vccd1 vccd1 _06463_/A sky130_fd_sc_hd__dfxtp_1
X_08201_ _08201_/A _08224_/Y vssd1 vssd1 vccd1 vccd1 _13801_/Z sky130_fd_sc_hd__ebufn_2
X_05413_ _05413_/A _05424_/Y vssd1 vssd1 vccd1 vccd1 _13813_/Z sky130_fd_sc_hd__ebufn_2
X_09181_ _09181_/A _09204_/Y vssd1 vssd1 vccd1 vccd1 _13661_/Z sky130_fd_sc_hd__ebufn_2
X_06393_ _06393_/A _06404_/Y vssd1 vssd1 vccd1 vccd1 _13673_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11142__D line[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05344_ _05350_/CLK line[54] vssd1 vssd1 vccd1 vccd1 _05345_/A sky130_fd_sc_hd__dfxtp_1
X_08132_ _08150_/CLK line[63] vssd1 vssd1 vccd1 vccd1 _08133_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06236__D line[92] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[6\].VALID\[1\].TOBUF OVHB\[6\].VALID\[1\].FF/Q OVHB\[6\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04926_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__05140__D line[89] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10981__D line[71] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08063_ _08063_/A _08084_/Y vssd1 vssd1 vccd1 vccd1 _13663_/Z sky130_fd_sc_hd__ebufn_2
X_05275_ _05275_/A _05284_/Y vssd1 vssd1 vccd1 vccd1 _13675_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_108_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07014_ _07030_/CLK line[49] vssd1 vssd1 vccd1 vccd1 _07015_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08451__D line[66] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13069__D line[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08965_ _08965_/A _08994_/Y vssd1 vssd1 vccd1 vccd1 _13725_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[12\].VALID\[14\].FF_D A[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07916_ _07940_/CLK line[92] vssd1 vssd1 vccd1 vccd1 _07917_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_57_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08896_ _08920_/CLK line[28] vssd1 vssd1 vccd1 vccd1 _08897_/A sky130_fd_sc_hd__dfxtp_1
X_07847_ _07847_/A _07874_/Y vssd1 vssd1 vccd1 vccd1 _13727_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_29_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11317__D line[111] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDATA\[26\].CLKBUF\[0\] clk vssd1 vssd1 vccd1 vccd1 _10007_/CLK sky130_fd_sc_hd__clkbuf_4
X_07778_ _07800_/CLK line[29] vssd1 vssd1 vccd1 vccd1 _07779_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05315__D line[41] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09517_ _09517_/CLK _09518_/X vssd1 vssd1 vccd1 vccd1 _09515_/CLK sky130_fd_sc_hd__dlclkp_1
X_06729_ _06729_/A _06754_/Y vssd1 vssd1 vccd1 vccd1 _13729_/Z sky130_fd_sc_hd__ebufn_2
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13532__D line[85] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDATA\[16\].CLKBUF\[6\] clk vssd1 vssd1 vccd1 vccd1 _07137_/CLK sky130_fd_sc_hd__clkbuf_4
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09448_ _13920_/Y wr vssd1 vssd1 vccd1 vccd1 _09448_/X sky130_fd_sc_hd__and2_1
XANTENNA__08626__D line[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMUX.M\[2\].MUX\[6\] _13675_/Z _13745_/Z _13815_/Z _13885_/Z MUX.SEL0BUF\[2\]/X MUX.SEL1BUF\[2\]/X
+ vssd1 vssd1 vccd1 vccd1 Do[22] sky130_fd_sc_hd__mux4_1
XFILLER_169_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09379_ _13916_/X vssd1 vssd1 vccd1 vccd1 _09379_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[22\].VALID\[13\].FF_D A[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08923__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11410_ _11440_/CLK line[16] vssd1 vssd1 vccd1 vccd1 _11411_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[12\].V_D TIE/HI vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05050__D line[62] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12390_ _12420_/CLK line[80] vssd1 vssd1 vccd1 vccd1 _12391_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_123_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10891__D line[44] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11341_ _11341_/A _11374_/Y vssd1 vssd1 vccd1 vccd1 _13861_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_125_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05985__D line[96] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[2\].VALID\[13\].FF OVHB\[2\].V/CLK A[20] vssd1 vssd1 vccd1 vccd1 OVHB\[2\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_11272_ _11300_/CLK line[90] vssd1 vssd1 vccd1 vccd1 _11273_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[27\].V_D TIE/HI vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13011_ _13015_/CLK line[103] vssd1 vssd1 vccd1 vccd1 _13012_/A sky130_fd_sc_hd__dfxtp_1
X_10223_ _10223_/A _10254_/Y vssd1 vssd1 vccd1 vccd1 _13863_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[5\].VALID\[5\].FF_D A[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MUX.M\[2\].MUX\[4\]_A3 _13881_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10154_ _10180_/CLK line[91] vssd1 vssd1 vccd1 vccd1 _10155_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13707__D line[37] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10085_ _10085_/A _10114_/Y vssd1 vssd1 vccd1 vccd1 _13725_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09192__D line[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13913_ _13916_/A _13916_/B _13916_/C _13916_/D vssd1 vssd1 vccd1 vccd1 _13913_/X
+ sky130_fd_sc_hd__and4bb_4
XOVHB\[22\].VALID\[14\].TOBUF OVHB\[22\].VALID\[14\].FF/Q OVHB\[22\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__10131__D line[66] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13844_ _13844_/A _13859_/Y vssd1 vssd1 vccd1 vccd1 _13844_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05225__D line[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13775_ _13785_/CLK line[68] vssd1 vssd1 vccd1 vccd1 _13776_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_16_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10987_ _10987_/CLK _10988_/X vssd1 vssd1 vccd1 vccd1 _10985_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__13442__D line[58] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12726_ _12726_/A _12739_/Y vssd1 vssd1 vccd1 vccd1 _13846_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_31_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07440__D line[116] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12058__D line[51] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12657_ _12665_/CLK line[69] vssd1 vssd1 vccd1 vccd1 _12658_/A sky130_fd_sc_hd__dfxtp_1
XPHY_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11608_ _11608_/A _11619_/Y vssd1 vssd1 vccd1 vccd1 _13848_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[15\].CLKBUF\[3\] clk vssd1 vssd1 vccd1 vccd1 _06752_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_129_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[0\].VALID\[1\].FF OVHB\[0\].V/CLK A[8] vssd1 vssd1 vccd1 vccd1 OVHB\[0\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_12588_ _12588_/A _12599_/Y vssd1 vssd1 vccd1 vccd1 _13708_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[14\].VALID\[10\].FF_D A[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11539_ _11545_/CLK line[70] vssd1 vssd1 vccd1 vccd1 _11540_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_209_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09367__D line[101] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05060_ _05070_/CLK line[52] vssd1 vssd1 vccd1 vccd1 _05061_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_143_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13209_ _13225_/CLK line[65] vssd1 vssd1 vccd1 vccd1 _13210_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10306__D line[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[26\].VALID\[11\].FF OVHB\[26\].V/CLK A[18] vssd1 vssd1 vccd1 vccd1 OVHB\[26\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13617__D line[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10603__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12521__D line[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08750_ _08780_/CLK line[80] vssd1 vssd1 vccd1 vccd1 _08751_/A sky130_fd_sc_hd__dfxtp_1
X_05962_ _05980_/CLK line[95] vssd1 vssd1 vccd1 vccd1 _05963_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_85_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07615__D line[68] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07701_ _07701_/A _07734_/Y vssd1 vssd1 vccd1 vccd1 _13861_/Z sky130_fd_sc_hd__ebufn_2
X_04913_ A_h[12] vssd1 vssd1 vccd1 vccd1 _04913_/Y sky130_fd_sc_hd__inv_2
X_08681_ _08681_/A _08714_/Y vssd1 vssd1 vccd1 vccd1 _13721_/Z sky130_fd_sc_hd__ebufn_2
X_05893_ _05893_/A _05914_/Y vssd1 vssd1 vccd1 vccd1 _13733_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[4\].VALID\[6\].TOBUF OVHB\[4\].VALID\[6\].FF/Q OVHB\[4\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04923_/A2 sky130_fd_sc_hd__ebufn_2
XFILLER_26_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XOVHB\[11\].VOBUF OVHB\[11\].V/Q OVHB\[11\].INV/Y vssd1 vssd1 vccd1 vccd1 _04912_/B1
+ sky130_fd_sc_hd__ebufn_2
X_07632_ _07660_/CLK line[90] vssd1 vssd1 vccd1 vccd1 _07633_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_19_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XOVHB\[29\].VALID\[9\].TOBUF OVHB\[29\].VALID\[9\].FF/Q OVHB\[29\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04914_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__09830__D line[57] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07563_ _07563_/A _07594_/Y vssd1 vssd1 vccd1 vccd1 _13723_/Z sky130_fd_sc_hd__ebufn_2
X_09302_ _09302_/A _09309_/Y vssd1 vssd1 vccd1 vccd1 _13782_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__04974__D line[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13930__A A[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06514_ _06540_/CLK line[91] vssd1 vssd1 vccd1 vccd1 _06515_/A sky130_fd_sc_hd__dfxtp_1
X_07494_ _07520_/CLK line[27] vssd1 vssd1 vccd1 vccd1 _07495_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_80_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07350__D line[80] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09233_ _09235_/CLK line[40] vssd1 vssd1 vccd1 vccd1 _09234_/A sky130_fd_sc_hd__dfxtp_1
X_06445_ _06445_/A _06474_/Y vssd1 vssd1 vccd1 vccd1 _13725_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_167_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09164_ _09164_/A _09169_/Y vssd1 vssd1 vccd1 vccd1 _13644_/Z sky130_fd_sc_hd__ebufn_2
X_06376_ _06400_/CLK line[28] vssd1 vssd1 vccd1 vccd1 _06377_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06544__A _13904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[11\].CLKBUF\[1\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08115_ _08115_/CLK line[41] vssd1 vssd1 vccd1 vccd1 _08116_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[16\].VALID\[13\].FF OVHB\[16\].V/CLK A[20] vssd1 vssd1 vccd1 vccd1 OVHB\[16\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_05327_ _05327_/A _05354_/Y vssd1 vssd1 vccd1 vccd1 _13727_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_135_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09095_ _09095_/CLK line[105] vssd1 vssd1 vccd1 vccd1 _09096_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_119_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06263__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09277__D line[74] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08181__D line[71] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08046_ _08046_/A _08049_/Y vssd1 vssd1 vccd1 vccd1 _13646_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_134_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05258_ _05280_/CLK line[29] vssd1 vssd1 vccd1 vccd1 _05259_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[14\].CLKBUF\[0\] clk vssd1 vssd1 vccd1 vccd1 _06367_/CLK sky130_fd_sc_hd__clkbuf_4
X_05189_ _05189_/A _05214_/Y vssd1 vssd1 vccd1 vccd1 _13869_/Z sky130_fd_sc_hd__ebufn_2
X_09997_ _10005_/CLK line[5] vssd1 vssd1 vccd1 vccd1 _09998_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_95_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12431__D line[108] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08948_ _08948_/A _08959_/Y vssd1 vssd1 vccd1 vccd1 _13708_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07525__D line[32] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08879_ _08885_/CLK line[6] vssd1 vssd1 vccd1 vccd1 _08880_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11047__D line[101] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10910_ _10910_/A _10919_/Y vssd1 vssd1 vccd1 vccd1 _13710_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_28_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11890_ _11890_/A _11899_/Y vssd1 vssd1 vccd1 vccd1 _13850_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[4\].CLKBUF\[1\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09740__D line[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06719__A _13905_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10841_ _10845_/CLK line[7] vssd1 vssd1 vccd1 vccd1 _10842_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06438__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13560_ _13560_/A _13579_/Y vssd1 vssd1 vccd1 vccd1 _13840_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08356__D line[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10772_ _10772_/A _10779_/Y vssd1 vssd1 vccd1 vccd1 _13852_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_44_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_DATA\[30\].CLKBUF\[3\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12511_ _12525_/CLK line[2] vssd1 vssd1 vccd1 vccd1 _12512_/A sky130_fd_sc_hd__dfxtp_1
X_13491_ _13505_/CLK line[66] vssd1 vssd1 vccd1 vccd1 _13492_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[11\].VALID\[1\].TOBUF OVHB\[11\].VALID\[1\].FF/Q OVHB\[11\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04926_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_157_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12442_ _12442_/A _12459_/Y vssd1 vssd1 vccd1 vccd1 _13842_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_60_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12373_ _12385_/CLK line[67] vssd1 vssd1 vccd1 vccd1 _12374_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12606__D line[60] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11510__D line[57] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08091__D line[44] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06604__D line[118] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11324_ _11324_/A _11339_/Y vssd1 vssd1 vccd1 vccd1 _13844_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_125_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11255_ _11265_/CLK line[68] vssd1 vssd1 vccd1 vccd1 _11256_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_69_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09915__D line[110] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10206_ _10206_/A _10219_/Y vssd1 vssd1 vccd1 vccd1 _13846_/Z sky130_fd_sc_hd__ebufn_2
X_11186_ _11186_/A _11199_/Y vssd1 vssd1 vccd1 vccd1 _13706_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_121_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10137_ _10145_/CLK line[69] vssd1 vssd1 vccd1 vccd1 _10138_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.M\[1\].MUX\[5\]_A1 _13694_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10068_ _10068_/A _10079_/Y vssd1 vssd1 vccd1 vccd1 _13708_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_48_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_OVHB\[19\].VALID\[14\].FF_D A[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10796__D line[114] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13827_ _13855_/CLK line[106] vssd1 vssd1 vccd1 vccd1 _13828_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_211_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13172__D line[63] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08266__D line[124] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13758_ _13758_/A _13789_/Y vssd1 vssd1 vccd1 vccd1 _13758_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07170__D line[121] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12709_ _12735_/CLK line[107] vssd1 vssd1 vccd1 vccd1 _12710_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_149_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13689_ _13715_/CLK line[43] vssd1 vssd1 vccd1 vccd1 _13690_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06230_ _06260_/CLK line[80] vssd1 vssd1 vccd1 vccd1 _06231_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[16\].INV _13953_/Y vssd1 vssd1 vccd1 vccd1 OVHB\[16\].INV/Y sky130_fd_sc_hd__inv_2
XANTENNA_OVHB\[29\].VALID\[13\].FF_D A[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06161_ _06161_/A _06194_/Y vssd1 vssd1 vccd1 vccd1 _13721_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_116_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11420__D line[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[13\].CGAND_B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05112_ _05140_/CLK line[90] vssd1 vssd1 vccd1 vccd1 _05113_/A sky130_fd_sc_hd__dfxtp_1
X_06092_ _06120_/CLK line[26] vssd1 vssd1 vccd1 vccd1 _06093_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06514__D line[91] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05043_ _05043_/A _05074_/Y vssd1 vssd1 vccd1 vccd1 _13723_/Z sky130_fd_sc_hd__ebufn_2
X_09920_ _09920_/A _09939_/Y vssd1 vssd1 vccd1 vccd1 _13840_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10036__D line[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_OVHB\[17\].CGAND_A _13910_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[10\].VALID\[1\].FF_D A[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09851_ _09865_/CLK line[66] vssd1 vssd1 vccd1 vccd1 _09852_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13347__D line[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08802_ _08802_/A _08819_/Y vssd1 vssd1 vccd1 vccd1 _13842_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_86_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09782_ _09782_/A _09799_/Y vssd1 vssd1 vccd1 vccd1 _13702_/Z sky130_fd_sc_hd__ebufn_2
X_06994_ _06994_/A _06999_/Y vssd1 vssd1 vccd1 vccd1 _13714_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07345__D line[73] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08733_ _08745_/CLK line[67] vssd1 vssd1 vccd1 vccd1 _08734_/A sky130_fd_sc_hd__dfxtp_1
X_05945_ _05945_/CLK line[73] vssd1 vssd1 vccd1 vccd1 _05946_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_73_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08664_ _08664_/A _08679_/Y vssd1 vssd1 vccd1 vccd1 _13704_/Z sky130_fd_sc_hd__ebufn_2
X_05876_ _05876_/A _05879_/Y vssd1 vssd1 vccd1 vccd1 _13716_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[18\].CGAND _13911_/X wr vssd1 vssd1 vccd1 vccd1 OVHB\[18\].CGAND/X sky130_fd_sc_hd__and2_4
XFILLER_54_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07615_ _07625_/CLK line[68] vssd1 vssd1 vccd1 vccd1 _07616_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08595_ _08605_/CLK line[4] vssd1 vssd1 vccd1 vccd1 _08596_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[29\].CLKBUF\[4\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07546_ _07546_/A _07559_/Y vssd1 vssd1 vccd1 vccd1 _13706_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07080__D line[94] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07477_ _07485_/CLK line[5] vssd1 vssd1 vccd1 vccd1 _07478_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_167_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13810__D line[84] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09216_ _09216_/A _09239_/Y vssd1 vssd1 vccd1 vccd1 _13696_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08904__D line[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06428_ _06428_/A _06439_/Y vssd1 vssd1 vccd1 vccd1 _13708_/Z sky130_fd_sc_hd__ebufn_2
X_09147_ _09165_/CLK line[15] vssd1 vssd1 vccd1 vccd1 _09148_/A sky130_fd_sc_hd__dfxtp_1
X_06359_ _06365_/CLK line[6] vssd1 vssd1 vccd1 vccd1 _06360_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_5_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[1\].VALID\[8\].FF_D A[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09078_ _09078_/A _09099_/Y vssd1 vssd1 vccd1 vccd1 _13838_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_190_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08029_ _08045_/CLK line[1] vssd1 vssd1 vccd1 vccd1 _08030_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_123_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11040_ _11040_/A _11059_/Y vssd1 vssd1 vccd1 vccd1 _13840_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_1_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12161__D line[98] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07255__D line[46] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[23\].VALID\[0\].FF OVHB\[23\].V/CLK A[7] vssd1 vssd1 vccd1 vccd1 OVHB\[23\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_12991_ _13015_/CLK line[108] vssd1 vssd1 vccd1 vccd1 _12992_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_29_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11942_ _11942_/A _11969_/Y vssd1 vssd1 vccd1 vccd1 _13622_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09470__D line[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05353__A _13900_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11873_ _11895_/CLK line[109] vssd1 vssd1 vccd1 vccd1 _11874_/A sky130_fd_sc_hd__dfxtp_1
X_13612_ _13612_/CLK _13613_/X vssd1 vssd1 vccd1 vccd1 _13610_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_72_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XOVHB\[12\].VALID\[11\].FF OVHB\[12\].V/CLK A[18] vssd1 vssd1 vccd1 vccd1 OVHB\[12\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_10824_ _10824_/A _10849_/Y vssd1 vssd1 vccd1 vccd1 _13624_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05503__D line[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[19\].VALID\[13\].TOBUF OVHB\[19\].VALID\[13\].FF/Q OVHB\[19\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04916_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_111_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13543_ _13898_/Y wr vssd1 vssd1 vccd1 vccd1 _13543_/X sky130_fd_sc_hd__and2_1
X_10755_ _10775_/CLK line[110] vssd1 vssd1 vccd1 vccd1 _10756_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[2\].CLKBUF\[3\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13720__D line[48] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13474_ _13898_/Y vssd1 vssd1 vccd1 vccd1 _13474_/Y sky130_fd_sc_hd__inv_2
X_10686_ _10686_/A _10709_/Y vssd1 vssd1 vccd1 vccd1 _13766_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_139_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12425_ _12455_/CLK line[96] vssd1 vssd1 vccd1 vccd1 _12426_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_173_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12336__D line[50] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12914__A _13937_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12356_ _12356_/A _12389_/Y vssd1 vssd1 vccd1 vccd1 _13756_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_154_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12633__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[23\].VALID\[1\].FF_D A[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11307_ _11335_/CLK line[106] vssd1 vssd1 vccd1 vccd1 _11308_/A sky130_fd_sc_hd__dfxtp_1
X_12287_ _12315_/CLK line[42] vssd1 vssd1 vccd1 vccd1 _12288_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_99_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09645__D line[100] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05528__A _13901_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11238_ _11238_/A _11269_/Y vssd1 vssd1 vccd1 vccd1 _13758_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_95_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11169_ _11195_/CLK line[43] vssd1 vssd1 vccd1 vccd1 _11170_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_OVHB\[16\].VALID\[5\].FF_D A[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[12\].VALID\[12\].TOBUF OVHB\[12\].VALID\[12\].FF/Q OVHB\[12\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04929_/B2 sky130_fd_sc_hd__ebufn_2
X_05730_ _05730_/A _05739_/Y vssd1 vssd1 vccd1 vccd1 _13850_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09380__D line[112] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05661_ _05665_/CLK line[71] vssd1 vssd1 vccd1 vccd1 _05662_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_35_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07400_ _07400_/A _07419_/Y vssd1 vssd1 vccd1 vccd1 _13840_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[21\].VALID\[2\].FF OVHB\[21\].V/CLK A[9] vssd1 vssd1 vccd1 vccd1 OVHB\[21\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_08380_ _08380_/A _08399_/Y vssd1 vssd1 vccd1 vccd1 _13700_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_211_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05592_ _05592_/A _05599_/Y vssd1 vssd1 vccd1 vccd1 _13712_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08574__A _13913_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12808__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07331_ _07345_/CLK line[66] vssd1 vssd1 vccd1 vccd1 _07332_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_189_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XDATA\[6\].CLKBUF\[7\] clk vssd1 vssd1 vccd1 vccd1 _13052_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__08293__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07262_ _07262_/A _07279_/Y vssd1 vssd1 vccd1 vccd1 _13702_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_149_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09001_ _09025_/CLK line[76] vssd1 vssd1 vccd1 vccd1 _09002_/A sky130_fd_sc_hd__dfxtp_1
X_06213_ _06225_/CLK line[67] vssd1 vssd1 vccd1 vccd1 _06214_/A sky130_fd_sc_hd__dfxtp_1
X_07193_ _07205_/CLK line[3] vssd1 vssd1 vccd1 vccd1 _07194_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_117_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11150__D line[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[18\].VALID\[1\].TOBUF OVHB\[18\].VALID\[1\].FF/Q OVHB\[18\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04926_/B2 sky130_fd_sc_hd__ebufn_2
XOVHB\[23\].CG clk OVHB\[23\].CGAND/X vssd1 vssd1 vccd1 vccd1 OVHB\[23\].V/CLK sky130_fd_sc_hd__dlclkp_1
X_06144_ _06144_/A _06159_/Y vssd1 vssd1 vccd1 vccd1 _13704_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06244__D line[81] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06075_ _06085_/CLK line[4] vssd1 vssd1 vccd1 vccd1 _06076_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09555__D line[64] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09903_ _13921_/X wr vssd1 vssd1 vccd1 vccd1 _09903_/X sky130_fd_sc_hd__and2_1
X_05026_ _05026_/A _05039_/Y vssd1 vssd1 vccd1 vccd1 _13706_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_160_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13077__D line[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[26\].V_RESET_B rst_n vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09834_ _13921_/X vssd1 vssd1 vccd1 vccd1 _09834_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08749__A _13914_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09765_ _09795_/CLK line[32] vssd1 vssd1 vccd1 vccd1 _09766_/A sky130_fd_sc_hd__dfxtp_1
X_06977_ _06995_/CLK line[47] vssd1 vssd1 vccd1 vccd1 _06978_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08468__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08716_ _08716_/A _08749_/Y vssd1 vssd1 vccd1 vccd1 _13756_/Z sky130_fd_sc_hd__ebufn_2
X_05928_ _05928_/A _05949_/Y vssd1 vssd1 vccd1 vccd1 _13768_/Z sky130_fd_sc_hd__ebufn_2
X_09696_ _09696_/A _09729_/Y vssd1 vssd1 vccd1 vccd1 _13616_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_26_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08647_ _08675_/CLK line[42] vssd1 vssd1 vccd1 vccd1 _08648_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05859_ _05875_/CLK line[33] vssd1 vssd1 vccd1 vccd1 _05860_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11325__D line[100] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06419__D line[33] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08578_ _08578_/A _08609_/Y vssd1 vssd1 vccd1 vccd1 _13618_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07529_ _07555_/CLK line[43] vssd1 vssd1 vccd1 vccd1 _07530_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13540__D line[89] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[7\].VALID\[13\].FF OVHB\[7\].V/CLK A[20] vssd1 vssd1 vccd1 vccd1 OVHB\[7\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_10540_ _10540_/A _10569_/Y vssd1 vssd1 vccd1 vccd1 _13620_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08634__D line[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_MUX.M\[3\].MUX\[6\]_A3 _13871_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10471_ _10495_/CLK line[108] vssd1 vssd1 vccd1 vccd1 _10472_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[27\].CLKBUF\[6\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11060__D line[112] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12210_ _12210_/CLK line[121] vssd1 vssd1 vccd1 vccd1 _12211_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[5\].CLKBUF\[4\] clk vssd1 vssd1 vccd1 vccd1 _12667_/CLK sky130_fd_sc_hd__clkbuf_4
X_13190_ _13190_/CLK line[57] vssd1 vssd1 vccd1 vccd1 _13191_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_203_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12141_ _12141_/A _12144_/Y vssd1 vssd1 vccd1 vccd1 _13821_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10254__A _13922_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05993__D line[109] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12072_ _12072_/CLK _12073_/X vssd1 vssd1 vccd1 vccd1 _12070_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA_OVHB\[29\].VALID\[5\].FF_D A[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11023_ _13925_/X wr vssd1 vssd1 vccd1 vccd1 _11023_/X sky130_fd_sc_hd__and2_1
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XOVHB\[24\].VALID\[0\].TOBUF OVHB\[24\].VALID\[0\].FF/Q OVHB\[24\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04924_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_66_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13715__D line[41] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08809__D line[102] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12974_ _12980_/CLK line[86] vssd1 vssd1 vccd1 vccd1 _12975_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_66_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11925_ _11925_/A _11934_/Y vssd1 vssd1 vccd1 vccd1 _13885_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11235__D line[64] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11856_ _11860_/CLK line[87] vssd1 vssd1 vccd1 vccd1 _11857_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_178_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05233__D line[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10807_ _10807_/A _10814_/Y vssd1 vssd1 vccd1 vccd1 _13887_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10429__A _13923_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11787_ _11787_/A _11794_/Y vssd1 vssd1 vccd1 vccd1 _13747_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13450__D line[62] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10738_ _10740_/CLK line[88] vssd1 vssd1 vccd1 vccd1 _10739_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08544__D line[123] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13526_ _13540_/CLK line[82] vssd1 vssd1 vccd1 vccd1 _13527_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_9_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10148__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[18\].VALID\[5\].FF OVHB\[18\].V/CLK A[12] vssd1 vssd1 vccd1 vccd1 OVHB\[18\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_174_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12066__D line[55] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13457_ _13457_/A _13474_/Y vssd1 vssd1 vccd1 vccd1 _13737_/Z sky130_fd_sc_hd__ebufn_2
X_10669_ _10669_/A _10674_/Y vssd1 vssd1 vccd1 vccd1 _13749_/Z sky130_fd_sc_hd__ebufn_2
X_12408_ _12420_/CLK line[83] vssd1 vssd1 vccd1 vccd1 _12409_/A sky130_fd_sc_hd__dfxtp_1
X_13388_ _13400_/CLK line[19] vssd1 vssd1 vccd1 vccd1 _13389_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_127_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_DATA\[0\].CLKBUF\[5\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12339_ _12339_/A _12354_/Y vssd1 vssd1 vccd1 vccd1 _13739_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[1\].V OVHB\[1\].V/CLK TIE/HI rst_n vssd1 vssd1 vccd1 vccd1 OVHB\[1\].V/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__09375__D line[105] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XDATA\[4\].CLKBUF\[1\] clk vssd1 vssd1 vccd1 vccd1 _12282_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_96_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06900_ _06900_/A _06929_/Y vssd1 vssd1 vccd1 vccd1 _13620_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10314__D line[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07880_ _07880_/A _07909_/Y vssd1 vssd1 vccd1 vccd1 _13760_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05408__D line[83] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06831_ _06855_/CLK line[108] vssd1 vssd1 vccd1 vccd1 _06832_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13625__D line[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09550_ _09550_/CLK line[57] vssd1 vssd1 vccd1 vccd1 _09551_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08719__D line[75] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06762_ _06762_/A _06789_/Y vssd1 vssd1 vccd1 vccd1 _13762_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06089__A _13903_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07623__D line[72] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08501_ _08501_/A _08504_/Y vssd1 vssd1 vccd1 vccd1 _13821_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[16\].VALID\[6\].TOBUF OVHB\[16\].VALID\[6\].FF/Q OVHB\[16\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04923_/A2 sky130_fd_sc_hd__ebufn_2
X_05713_ _05735_/CLK line[109] vssd1 vssd1 vccd1 vccd1 _05714_/A sky130_fd_sc_hd__dfxtp_1
X_09481_ _09481_/A _09484_/Y vssd1 vssd1 vccd1 vccd1 _13681_/Z sky130_fd_sc_hd__ebufn_2
X_06693_ _06715_/CLK line[45] vssd1 vssd1 vccd1 vccd1 _06694_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11723__A _13927_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08432_ _08432_/CLK _08433_/X vssd1 vssd1 vccd1 vccd1 _08430_/CLK sky130_fd_sc_hd__dlclkp_1
X_05644_ _05644_/A _05669_/Y vssd1 vssd1 vccd1 vccd1 _13764_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_211_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08363_ _13913_/X wr vssd1 vssd1 vccd1 vccd1 _08363_/X sky130_fd_sc_hd__and2_1
XFILLER_11_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05575_ _05595_/CLK line[46] vssd1 vssd1 vccd1 vccd1 _05576_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__04982__D line[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07314_ _13910_/X vssd1 vssd1 vccd1 vccd1 _07314_/Y sky130_fd_sc_hd__inv_2
X_08294_ _13932_/X vssd1 vssd1 vccd1 vccd1 _08294_/Y sky130_fd_sc_hd__inv_2
XFILLER_149_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07245_ _07275_/CLK line[32] vssd1 vssd1 vccd1 vccd1 _07246_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[24\].CLKBUF\[5\] clk vssd1 vssd1 vccd1 vccd1 _09622_/CLK sky130_fd_sc_hd__clkbuf_4
X_07176_ _07176_/A _07209_/Y vssd1 vssd1 vccd1 vccd1 _13616_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_117_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06127_ _06155_/CLK line[42] vssd1 vssd1 vccd1 vccd1 _06128_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_127_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09285__D line[78] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XOVHB\[16\].VALID\[7\].FF OVHB\[16\].V/CLK A[14] vssd1 vssd1 vccd1 vccd1 OVHB\[16\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_06058_ _06058_/A _06089_/Y vssd1 vssd1 vccd1 vccd1 _13618_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10224__D line[123] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05009_ _05035_/CLK line[43] vssd1 vssd1 vccd1 vccd1 _05010_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_160_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07383__A _13910_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09817_ _09817_/A _09834_/Y vssd1 vssd1 vccd1 vccd1 _13737_/Z sky130_fd_sc_hd__ebufn_2
X_09748_ _09760_/CLK line[19] vssd1 vssd1 vccd1 vccd1 _09749_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_39_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07533__D line[45] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09679_ _09679_/A _09694_/Y vssd1 vssd1 vccd1 vccd1 _13879_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_36_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11055__D line[105] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11710_ _11720_/CLK line[20] vssd1 vssd1 vccd1 vccd1 _11711_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_36_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06149__D line[38] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12690_ _12700_/CLK line[84] vssd1 vssd1 vccd1 vccd1 _12691_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11641_ _11641_/A _11654_/Y vssd1 vssd1 vccd1 vccd1 _13881_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11572_ _11580_/CLK line[85] vssd1 vssd1 vccd1 vccd1 _11573_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[28\].CG_CLK clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13311_ _13311_/A _13334_/Y vssd1 vssd1 vccd1 vccd1 _13871_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10523_ _10523_/A _10534_/Y vssd1 vssd1 vccd1 vccd1 _13883_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[22\].VALID\[5\].TOBUF OVHB\[22\].VALID\[5\].FF/Q OVHB\[22\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04927_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_6_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07558__A _13911_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13242_ _13260_/CLK line[95] vssd1 vssd1 vccd1 vccd1 _13243_/A sky130_fd_sc_hd__dfxtp_1
X_10454_ _10460_/CLK line[86] vssd1 vssd1 vccd1 vccd1 _10455_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_124_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MUX.M\[2\].MUX\[7\]_A1 _13747_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13173_ _13173_/A _13194_/Y vssd1 vssd1 vccd1 vccd1 _13733_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12614__D line[49] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10385_ _10385_/A _10394_/Y vssd1 vssd1 vccd1 vccd1 _13745_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_184_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07708__D line[125] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12124_ _12140_/CLK line[81] vssd1 vssd1 vccd1 vccd1 _12125_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[23\].CLKBUF\[2\] clk vssd1 vssd1 vccd1 vccd1 _09237_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_2_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[12\].VALID\[8\].FF_D A[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12055_ _12055_/A _12074_/Y vssd1 vssd1 vccd1 vccd1 _13735_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_77_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09923__D line[99] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11006_ _11020_/CLK line[82] vssd1 vssd1 vccd1 vccd1 _11007_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[14\].VALID\[9\].FF OVHB\[14\].V/CLK A[16] vssd1 vssd1 vccd1 vccd1 OVHB\[14\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XOVHB\[3\].VALID\[11\].FF OVHB\[3\].V/CLK A[18] vssd1 vssd1 vccd1 vccd1 OVHB\[3\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_12957_ _12957_/A _12984_/Y vssd1 vssd1 vccd1 vccd1 _13797_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_18_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06059__D line[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11908_ _11930_/CLK line[125] vssd1 vssd1 vccd1 vccd1 _11909_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.M\[0\].MUX\[3\]_A2 _13774_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12888_ _12910_/CLK line[61] vssd1 vssd1 vccd1 vccd1 _12889_/A sky130_fd_sc_hd__dfxtp_1
X_11839_ _11839_/A _11864_/Y vssd1 vssd1 vccd1 vccd1 _13799_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13180__D line[52] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05898__D line[51] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05360_ _05360_/A _05389_/Y vssd1 vssd1 vccd1 vccd1 _13760_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08274__D line[113] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13509_ _13898_/Y vssd1 vssd1 vccd1 vccd1 _13509_/Y sky130_fd_sc_hd__inv_2
X_05291_ _05315_/CLK line[44] vssd1 vssd1 vccd1 vccd1 _05292_/A sky130_fd_sc_hd__dfxtp_1
X_07030_ _07030_/CLK line[57] vssd1 vssd1 vccd1 vccd1 _07031_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_170_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06522__D line[95] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08981_ _08981_/A _08994_/Y vssd1 vssd1 vccd1 vccd1 _13741_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_114_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07932_ _07940_/CLK line[85] vssd1 vssd1 vccd1 vccd1 _07933_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05138__D line[88] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10979__D line[70] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07863_ _07863_/A _07874_/Y vssd1 vssd1 vccd1 vccd1 _13743_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13355__D line[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09602_ _09620_/CLK line[95] vssd1 vssd1 vccd1 vccd1 _09603_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_68_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06814_ _06820_/CLK line[86] vssd1 vssd1 vccd1 vccd1 _06815_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08449__D line[65] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07794_ _07800_/CLK line[22] vssd1 vssd1 vccd1 vccd1 _07795_/A sky130_fd_sc_hd__dfxtp_1
X_09533_ _09533_/A _09554_/Y vssd1 vssd1 vccd1 vccd1 _13733_/Z sky130_fd_sc_hd__ebufn_2
X_06745_ _06745_/A _06754_/Y vssd1 vssd1 vccd1 vccd1 _13745_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[12\].CLKBUF\[5\] clk vssd1 vssd1 vccd1 vccd1 _05982_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_24_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09464_ _09480_/CLK line[17] vssd1 vssd1 vccd1 vccd1 _09465_/A sky130_fd_sc_hd__dfxtp_1
X_06676_ _06680_/CLK line[23] vssd1 vssd1 vccd1 vccd1 _06677_/A sky130_fd_sc_hd__dfxtp_1
XPHY_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08415_ _08415_/A _08434_/Y vssd1 vssd1 vccd1 vccd1 _13735_/Z sky130_fd_sc_hd__ebufn_2
X_05627_ _05627_/A _05634_/Y vssd1 vssd1 vccd1 vccd1 _13747_/Z sky130_fd_sc_hd__ebufn_2
X_09395_ _09395_/A _09414_/Y vssd1 vssd1 vccd1 vccd1 _13875_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13090__D line[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11603__D line[99] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08346_ _08360_/CLK line[18] vssd1 vssd1 vccd1 vccd1 _08347_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05558_ _05560_/CLK line[24] vssd1 vssd1 vccd1 vccd1 _05559_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_11_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08277_ _08277_/A _08294_/Y vssd1 vssd1 vccd1 vccd1 _13877_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12284__A _13935_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05489_ _05489_/A _05494_/Y vssd1 vssd1 vccd1 vccd1 _13889_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_137_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07228_ _07240_/CLK line[19] vssd1 vssd1 vccd1 vccd1 _07229_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_138_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08912__D line[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07159_ _07159_/A _07174_/Y vssd1 vssd1 vccd1 vccd1 _13879_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[25\].VALID\[8\].FF_D A[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10170_ _10180_/CLK line[84] vssd1 vssd1 vccd1 vccd1 _10171_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_78_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[9\].VALID\[0\].FF OVHB\[9\].V/CLK A[7] vssd1 vssd1 vccd1 vccd1 OVHB\[9\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_120_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XOVHB\[29\].VALID\[11\].TOBUF OVHB\[29\].VALID\[11\].FF/Q OVHB\[29\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04915_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__05048__D line[61] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[2\].VALID\[14\].TOBUF OVHB\[2\].VALID\[14\].FF/Q OVHB\[2\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_75_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10889__D line[43] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[17\].VALID\[11\].FF OVHB\[17\].V/CLK A[18] vssd1 vssd1 vccd1 vccd1 OVHB\[17\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13265__D line[96] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13860_ _13890_/CLK line[112] vssd1 vssd1 vccd1 vccd1 _13861_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07263__D line[35] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12811_ _12811_/A _12844_/Y vssd1 vssd1 vccd1 vccd1 _13651_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_27_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12459__A _13935_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13791_ _13791_/A _13824_/Y vssd1 vssd1 vccd1 vccd1 _13791_/Z sky130_fd_sc_hd__ebufn_2
X_12742_ _12770_/CLK line[122] vssd1 vssd1 vccd1 vccd1 _12743_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12178__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12673_ _12673_/A _12704_/Y vssd1 vssd1 vccd1 vccd1 _13793_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XDATA\[11\].CLKBUF\[2\] clk vssd1 vssd1 vccd1 vccd1 _05597_/CLK sky130_fd_sc_hd__clkbuf_4
XPHY_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11624_ _11650_/CLK line[123] vssd1 vssd1 vccd1 vccd1 _11625_/A sky130_fd_sc_hd__dfxtp_1
XPHY_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05511__D line[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11555_ _11555_/A _11584_/Y vssd1 vssd1 vccd1 vccd1 _13795_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10129__D line[65] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10506_ _10530_/CLK line[124] vssd1 vssd1 vccd1 vccd1 _10507_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08822__D line[122] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11486_ _11510_/CLK line[60] vssd1 vssd1 vccd1 vccd1 _11487_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_109_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XOVHB\[22\].VALID\[10\].TOBUF OVHB\[22\].VALID\[10\].FF/Q OVHB\[22\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04932_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_6_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13225_ _13225_/CLK line[73] vssd1 vssd1 vccd1 vccd1 _13226_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_170_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12344__D line[54] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10437_ _10437_/A _10464_/Y vssd1 vssd1 vccd1 vccd1 _13797_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07438__D line[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[6\].VALID\[13\].FF_D A[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13156_ _13156_/A _13159_/Y vssd1 vssd1 vccd1 vccd1 _13716_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_112_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10368_ _10390_/CLK line[61] vssd1 vssd1 vccd1 vccd1 _10369_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_151_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12107_ _12107_/CLK _12108_/X vssd1 vssd1 vccd1 vccd1 _12105_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_97_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13087_ _13087_/CLK _13088_/X vssd1 vssd1 vccd1 vccd1 _13085_/CLK sky130_fd_sc_hd__dlclkp_1
X_10299_ _10299_/A _10324_/Y vssd1 vssd1 vccd1 vccd1 _13659_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09653__D line[104] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12038_ _13934_/X wr vssd1 vssd1 vccd1 vccd1 _12038_/X sky130_fd_sc_hd__and2_1
XFILLER_93_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13753__A _13899_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_OVHB\[6\].VALID\[3\].FF_D A[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XOVHB\[7\].VALID\[2\].FF OVHB\[7\].V/CLK A[9] vssd1 vssd1 vccd1 vccd1 OVHB\[7\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_06530_ _06540_/CLK line[84] vssd1 vssd1 vccd1 vccd1 _06531_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07901__D line[71] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12519__D line[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06461_ _06461_/A _06474_/Y vssd1 vssd1 vccd1 vccd1 _13741_/Z sky130_fd_sc_hd__ebufn_2
X_08200_ _08220_/CLK line[94] vssd1 vssd1 vccd1 vccd1 _08201_/A sky130_fd_sc_hd__dfxtp_1
X_05412_ _05420_/CLK line[85] vssd1 vssd1 vccd1 vccd1 _05413_/A sky130_fd_sc_hd__dfxtp_1
X_09180_ _09200_/CLK line[30] vssd1 vssd1 vccd1 vccd1 _09181_/A sky130_fd_sc_hd__dfxtp_1
X_06392_ _06400_/CLK line[21] vssd1 vssd1 vccd1 vccd1 _06393_/A sky130_fd_sc_hd__dfxtp_1
X_08131_ _08131_/A _08154_/Y vssd1 vssd1 vccd1 vccd1 _13731_/Z sky130_fd_sc_hd__ebufn_2
X_05343_ _05343_/A _05354_/Y vssd1 vssd1 vccd1 vccd1 _13743_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09828__D line[56] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[4\].VALID\[2\].TOBUF OVHB\[4\].VALID\[2\].FF/Q OVHB\[4\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04930_/B2 sky130_fd_sc_hd__ebufn_2
X_08062_ _08080_/CLK line[31] vssd1 vssd1 vccd1 vccd1 _08063_/A sky130_fd_sc_hd__dfxtp_1
X_05274_ _05280_/CLK line[22] vssd1 vssd1 vccd1 vccd1 _05275_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_134_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07013_ _07013_/A _07034_/Y vssd1 vssd1 vccd1 vccd1 _13733_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12254__D line[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13928__A A[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[29\].VALID\[5\].TOBUF OVHB\[29\].VALID\[5\].FF/Q OVHB\[29\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04927_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06252__D line[85] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08964_ _08990_/CLK line[59] vssd1 vssd1 vccd1 vccd1 _08965_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09563__D line[77] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07915_ _07915_/A _07944_/Y vssd1 vssd1 vccd1 vccd1 _13795_/Z sky130_fd_sc_hd__ebufn_2
X_08895_ _08895_/A _08924_/Y vssd1 vssd1 vccd1 vccd1 _13655_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13085__D line[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10502__D line[122] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07846_ _07870_/CLK line[60] vssd1 vssd1 vccd1 vccd1 _07847_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08179__D line[70] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07777_ _07777_/A _07804_/Y vssd1 vssd1 vccd1 vccd1 _13657_/Z sky130_fd_sc_hd__ebufn_2
X_04989_ _04989_/A _05004_/Y vssd1 vssd1 vccd1 vccd1 _13669_/Z sky130_fd_sc_hd__ebufn_2
X_09516_ _09516_/A _09519_/Y vssd1 vssd1 vccd1 vccd1 _13716_/Z sky130_fd_sc_hd__ebufn_2
X_06728_ _06750_/CLK line[61] vssd1 vssd1 vccd1 vccd1 _06729_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_197_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07811__D line[44] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09447_ _09447_/CLK _09448_/X vssd1 vssd1 vccd1 vccd1 _09445_/CLK sky130_fd_sc_hd__dlclkp_1
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06659_ _06659_/A _06684_/Y vssd1 vssd1 vccd1 vccd1 _13659_/Z sky130_fd_sc_hd__ebufn_2
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12429__D line[107] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11333__D line[104] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06427__D line[37] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09588__A _13920_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09378_ _13916_/X wr vssd1 vssd1 vccd1 vccd1 _09378_/X sky130_fd_sc_hd__and2_1
XFILLER_149_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XOVHB\[5\].VALID\[4\].FF OVHB\[5\].V/CLK A[11] vssd1 vssd1 vccd1 vccd1 OVHB\[5\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_08329_ _13913_/X vssd1 vssd1 vccd1 vccd1 _08329_/Y sky130_fd_sc_hd__inv_2
XANTENNA__09738__D line[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11340_ _11370_/CLK line[112] vssd1 vssd1 vccd1 vccd1 _11341_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_125_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11271_ _11271_/A _11304_/Y vssd1 vssd1 vccd1 vccd1 _13791_/Z sky130_fd_sc_hd__ebufn_2
X_13010_ _13010_/A _13019_/Y vssd1 vssd1 vccd1 vccd1 _13850_/Z sky130_fd_sc_hd__ebufn_2
X_10222_ _10250_/CLK line[122] vssd1 vssd1 vccd1 vccd1 _10223_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06162__D line[58] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10153_ _10153_/A _10184_/Y vssd1 vssd1 vccd1 vccd1 _13793_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_160_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10084_ _10110_/CLK line[59] vssd1 vssd1 vccd1 vccd1 _10085_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_47_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11508__D line[56] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08089__D line[43] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13912_ _13916_/C _13916_/B _13916_/A _13916_/D vssd1 vssd1 vccd1 vccd1 _13912_/X
+ sky130_fd_sc_hd__and4b_4
XFILLER_74_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13843_ _13855_/CLK line[99] vssd1 vssd1 vccd1 vccd1 _13844_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11093__A _13925_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[18\].CLKBUF\[2\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13774_ _13774_/A _13789_/Y vssd1 vssd1 vccd1 vccd1 _13774_/Z sky130_fd_sc_hd__ebufn_2
X_10986_ _10986_/A _10989_/Y vssd1 vssd1 vccd1 vccd1 _13786_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_15_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12725_ _12735_/CLK line[100] vssd1 vssd1 vccd1 vccd1 _12726_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11243__D line[77] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06337__D line[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05241__D line[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12656_ _12656_/A _12669_/Y vssd1 vssd1 vccd1 vccd1 _13776_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11607_ _11615_/CLK line[101] vssd1 vssd1 vccd1 vccd1 _11608_/A sky130_fd_sc_hd__dfxtp_1
X_12587_ _12595_/CLK line[37] vssd1 vssd1 vccd1 vccd1 _12588_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08552__D line[127] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11538_ _11538_/A _11549_/Y vssd1 vssd1 vccd1 vccd1 _13778_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_7_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11469_ _11475_/CLK line[38] vssd1 vssd1 vccd1 vccd1 _11470_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[28\].V OVHB\[28\].V/CLK TIE/HI rst_n vssd1 vssd1 vccd1 vccd1 OVHB\[28\].V/Q
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07168__D line[120] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13208_ _13208_/A _13229_/Y vssd1 vssd1 vccd1 vccd1 _13768_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[3\].VALID\[6\].FF OVHB\[3\].V/CLK A[13] vssd1 vssd1 vccd1 vccd1 OVHB\[3\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11268__A _13933_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13139_ _13155_/CLK line[33] vssd1 vssd1 vccd1 vccd1 _13140_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06800__D line[94] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05961_ _05961_/A _05984_/Y vssd1 vssd1 vccd1 vccd1 _13801_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11418__D line[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07700_ _07730_/CLK line[112] vssd1 vssd1 vccd1 vccd1 _07701_/A sky130_fd_sc_hd__dfxtp_1
X_04912_ _04911_/Y _04914_/B2 _04912_/B1 vssd1 vssd1 vccd1 vccd1 _04917_/A sky130_fd_sc_hd__o21ai_2
X_08680_ _08710_/CLK line[48] vssd1 vssd1 vccd1 vccd1 _08681_/A sky130_fd_sc_hd__dfxtp_1
X_05892_ _05910_/CLK line[63] vssd1 vssd1 vccd1 vccd1 _05893_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05416__D line[87] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07631_ _07631_/A _07664_/Y vssd1 vssd1 vccd1 vccd1 _13791_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[2\].VALID\[7\].TOBUF OVHB\[2\].VALID\[7\].FF/Q OVHB\[2\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/A2 sky130_fd_sc_hd__ebufn_2
XANTENNA__13633__D line[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08727__D line[79] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07562_ _07590_/CLK line[58] vssd1 vssd1 vccd1 vccd1 _07563_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_179_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09301_ _09305_/CLK line[71] vssd1 vssd1 vccd1 vccd1 _09302_/A sky130_fd_sc_hd__dfxtp_1
X_06513_ _06513_/A _06544_/Y vssd1 vssd1 vccd1 vccd1 _13793_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_179_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07493_ _07493_/A _07524_/Y vssd1 vssd1 vccd1 vccd1 _13653_/Z sky130_fd_sc_hd__ebufn_2
XMUX.SEL0BUF\[3\] A[0] vssd1 vssd1 vccd1 vccd1 MUX.SEL0BUF\[3\]/X sky130_fd_sc_hd__clkbuf_2
X_09232_ _09232_/A _09239_/Y vssd1 vssd1 vccd1 vccd1 _13712_/Z sky130_fd_sc_hd__ebufn_2
X_06444_ _06470_/CLK line[59] vssd1 vssd1 vccd1 vccd1 _06445_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_139_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05151__D line[108] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09163_ _09165_/CLK line[8] vssd1 vssd1 vccd1 vccd1 _09164_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10992__D line[90] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06375_ _06375_/A _06404_/Y vssd1 vssd1 vccd1 vccd1 _13655_/Z sky130_fd_sc_hd__ebufn_2
X_08114_ _08114_/A _08119_/Y vssd1 vssd1 vccd1 vccd1 _13714_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_108_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__04990__D line[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05326_ _05350_/CLK line[60] vssd1 vssd1 vccd1 vccd1 _05327_/A sky130_fd_sc_hd__dfxtp_1
X_09094_ _09094_/A _09099_/Y vssd1 vssd1 vccd1 vccd1 _13854_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_107_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[14\].CGAND _13904_/X wr vssd1 vssd1 vccd1 vccd1 OVHB\[14\].CGAND/X sky130_fd_sc_hd__and2_4
X_08045_ _08045_/CLK line[9] vssd1 vssd1 vccd1 vccd1 _08046_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_119_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05257_ _05257_/A _05284_/Y vssd1 vssd1 vccd1 vccd1 _13657_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07078__D line[93] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[19\].V OVHB\[19\].V/CLK TIE/HI rst_n vssd1 vssd1 vccd1 vccd1 OVHB\[19\].V/Q
+ sky130_fd_sc_hd__dfrtp_1
XOVHB\[31\].VALID\[0\].FF OVHB\[31\].V/CLK A[7] vssd1 vssd1 vccd1 vccd1 OVHB\[31\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__09053__TE_B _09064_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05188_ _05210_/CLK line[125] vssd1 vssd1 vccd1 vccd1 _05189_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_88_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13808__D line[83] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09996_ _09996_/A _10009_/Y vssd1 vssd1 vccd1 vccd1 _13636_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_88_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09293__D line[67] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08947_ _08955_/CLK line[37] vssd1 vssd1 vccd1 vccd1 _08948_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10232__D line[127] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08878_ _08878_/A _08889_/Y vssd1 vssd1 vccd1 vccd1 _13638_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05326__D line[60] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XOVHB\[1\].VALID\[8\].FF OVHB\[1\].V/CLK A[15] vssd1 vssd1 vccd1 vccd1 OVHB\[1\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_29_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07829_ _07835_/CLK line[38] vssd1 vssd1 vccd1 vccd1 _07830_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_205_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10840_ _10840_/A _10849_/Y vssd1 vssd1 vccd1 vccd1 _13640_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_72_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07541__D line[34] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10771_ _10775_/CLK line[103] vssd1 vssd1 vccd1 vccd1 _10772_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12159__D line[97] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12510_ _12510_/A _12529_/Y vssd1 vssd1 vccd1 vccd1 _13630_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_52_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13490_ _13490_/A _13509_/Y vssd1 vssd1 vccd1 vccd1 _13770_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_200_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11998__D line[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12441_ _12455_/CLK line[98] vssd1 vssd1 vccd1 vccd1 _12442_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09468__D line[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12372_ _12372_/A _12389_/Y vssd1 vssd1 vccd1 vccd1 _13772_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_60_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11323_ _11335_/CLK line[99] vssd1 vssd1 vccd1 vccd1 _11324_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10407__D line[79] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11254_ _11254_/A _11269_/Y vssd1 vssd1 vccd1 vccd1 _13774_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_122_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10205_ _10215_/CLK line[100] vssd1 vssd1 vccd1 vccd1 _10206_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12622__D line[53] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11185_ _11195_/CLK line[36] vssd1 vssd1 vccd1 vccd1 _11186_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[8\].VALID\[11\].FF OVHB\[8\].V/CLK A[18] vssd1 vssd1 vccd1 vccd1 OVHB\[8\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07716__D line[114] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10136_ _10136_/A _10149_/Y vssd1 vssd1 vccd1 vccd1 _13776_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.M\[1\].MUX\[5\]_A2 _13764_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10067_ _10075_/CLK line[37] vssd1 vssd1 vccd1 vccd1 _10068_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[2\].VALID\[6\].FF_D A[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09931__D line[103] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13826_ _13826_/A _13859_/Y vssd1 vssd1 vccd1 vccd1 _13826_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[2\].CLKBUF\[6\] clk vssd1 vssd1 vccd1 vccd1 _11337_/CLK sky130_fd_sc_hd__clkbuf_4
X_13757_ _13785_/CLK line[74] vssd1 vssd1 vccd1 vccd1 _13758_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_204_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10969_ _10985_/CLK line[65] vssd1 vssd1 vccd1 vccd1 _10970_/A sky130_fd_sc_hd__dfxtp_1
X_12708_ _12708_/A _12739_/Y vssd1 vssd1 vccd1 vccd1 _13828_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06067__D line[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13688_ _13688_/A _13719_/Y vssd1 vssd1 vccd1 vccd1 _13688_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_148_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12639_ _12665_/CLK line[75] vssd1 vssd1 vccd1 vccd1 _12640_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[16\].CLKBUF\[4\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06160_ _06190_/CLK line[48] vssd1 vssd1 vccd1 vccd1 _06161_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08282__D line[117] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05111_ _05111_/A _05144_/Y vssd1 vssd1 vccd1 vccd1 _13791_/Z sky130_fd_sc_hd__ebufn_2
X_06091_ _06091_/A _06124_/Y vssd1 vssd1 vccd1 vccd1 _13651_/Z sky130_fd_sc_hd__ebufn_2
X_05042_ _05070_/CLK line[58] vssd1 vssd1 vccd1 vccd1 _05043_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_131_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[17\].CGAND_B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12532__D line[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09850_ _09850_/A _09869_/Y vssd1 vssd1 vccd1 vccd1 _13770_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[25\].V_RESET_B rst_n vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08801_ _08815_/CLK line[98] vssd1 vssd1 vccd1 vccd1 _08802_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06530__D line[84] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[28\].VALID\[3\].FF OVHB\[28\].V/CLK A[10] vssd1 vssd1 vccd1 vccd1 OVHB\[28\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_06993_ _06995_/CLK line[40] vssd1 vssd1 vccd1 vccd1 _06994_/A sky130_fd_sc_hd__dfxtp_1
X_09781_ _09795_/CLK line[34] vssd1 vssd1 vccd1 vccd1 _09782_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11148__D line[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08732_ _08732_/A _08749_/Y vssd1 vssd1 vccd1 vccd1 _13772_/Z sky130_fd_sc_hd__ebufn_2
X_05944_ _05944_/A _05949_/Y vssd1 vssd1 vccd1 vccd1 _13784_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[11\].V_D TIE/HI vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[9\].CLKBUF\[4\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09841__D line[76] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08663_ _08675_/CLK line[35] vssd1 vssd1 vccd1 vccd1 _08664_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_26_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05875_ _05875_/CLK line[41] vssd1 vssd1 vccd1 vccd1 _05876_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13363__D line[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13941__A A_h[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08457__D line[69] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07614_ _07614_/A _07629_/Y vssd1 vssd1 vccd1 vccd1 _13774_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_121_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08594_ _08594_/A _08609_/Y vssd1 vssd1 vccd1 vccd1 _13634_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[10\].VALID\[0\].FF OVHB\[10\].V/CLK A[7] vssd1 vssd1 vccd1 vccd1 OVHB\[10\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07545_ _07555_/CLK line[36] vssd1 vssd1 vccd1 vccd1 _07546_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[26\].V_D TIE/HI vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07476_ _07476_/A _07489_/Y vssd1 vssd1 vccd1 vccd1 _13636_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[17\].VALID\[3\].FF_D A[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[8\].VOBUF OVHB\[8\].V/Q OVHB\[8\].INV/Y vssd1 vssd1 vccd1 vccd1 _04912_/B1
+ sky130_fd_sc_hd__ebufn_2
X_06427_ _06435_/CLK line[37] vssd1 vssd1 vccd1 vccd1 _06428_/A sky130_fd_sc_hd__dfxtp_1
X_09215_ _09235_/CLK line[46] vssd1 vssd1 vccd1 vccd1 _09216_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_210_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12707__D line[106] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDATA\[1\].CLKBUF\[3\] clk vssd1 vssd1 vccd1 vccd1 _08152_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_194_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11611__D line[103] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09146_ _09146_/A _09169_/Y vssd1 vssd1 vccd1 vccd1 _13626_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[23\].VALID\[14\].FF_D A[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08192__D line[90] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06358_ _06358_/A _06369_/Y vssd1 vssd1 vccd1 vccd1 _13638_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06705__D line[36] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05309_ _05315_/CLK line[38] vssd1 vssd1 vccd1 vccd1 _05310_/A sky130_fd_sc_hd__dfxtp_1
X_09077_ _09095_/CLK line[111] vssd1 vssd1 vccd1 vccd1 _09078_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_163_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06289_ _06295_/CLK line[102] vssd1 vssd1 vccd1 vccd1 _06290_/A sky130_fd_sc_hd__dfxtp_1
X_08028_ _08028_/A _08049_/Y vssd1 vssd1 vccd1 vccd1 _13628_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08920__D line[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13538__D line[88] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06440__D line[48] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09979_ _10005_/CLK line[11] vssd1 vssd1 vccd1 vccd1 _09980_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05056__D line[50] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[15\].VALID\[14\].TOBUF OVHB\[15\].VALID\[14\].FF/Q OVHB\[15\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/B2 sky130_fd_sc_hd__ebufn_2
X_12990_ _12990_/A _13019_/Y vssd1 vssd1 vccd1 vccd1 _13830_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_183_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05634__A _13901_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDATA\[31\].CLKBUF\[1\] clk vssd1 vssd1 vccd1 vccd1 _11722_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__10897__D line[47] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11941_ _11965_/CLK line[12] vssd1 vssd1 vccd1 vccd1 _11942_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_91_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13273__D line[109] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05353__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08367__D line[42] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11872_ _11872_/A _11899_/Y vssd1 vssd1 vccd1 vccd1 _13832_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07271__D line[39] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[26\].VALID\[5\].FF OVHB\[26\].V/CLK A[12] vssd1 vssd1 vccd1 vccd1 OVHB\[26\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_44_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XDATA\[21\].CLKBUF\[7\] clk vssd1 vssd1 vccd1 vccd1 _08852_/CLK sky130_fd_sc_hd__clkbuf_4
X_13611_ _13611_/A _13614_/Y vssd1 vssd1 vccd1 vccd1 _13891_/Z sky130_fd_sc_hd__ebufn_2
X_10823_ _10845_/CLK line[13] vssd1 vssd1 vccd1 vccd1 _10824_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[9\].VALID\[7\].TOBUF OVHB\[9\].VALID\[7\].FF/Q OVHB\[9\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/A2 sky130_fd_sc_hd__ebufn_2
XFILLER_60_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13542_ _13542_/CLK _13543_/X vssd1 vssd1 vccd1 vccd1 _13540_/CLK sky130_fd_sc_hd__dlclkp_1
X_10754_ _10754_/A _10779_/Y vssd1 vssd1 vccd1 vccd1 _13834_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_158_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10685_ _10705_/CLK line[78] vssd1 vssd1 vccd1 vccd1 _10686_/A sky130_fd_sc_hd__dfxtp_1
X_13473_ _13898_/Y wr vssd1 vssd1 vccd1 vccd1 _13473_/X sky130_fd_sc_hd__and2_1
XANTENNA__11521__D line[76] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09198__D line[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06615__D line[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12424_ _13935_/X vssd1 vssd1 vccd1 vccd1 _12424_/Y sky130_fd_sc_hd__inv_2
XFILLER_166_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10137__D line[69] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13298__A _13938_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12355_ _12385_/CLK line[64] vssd1 vssd1 vccd1 vccd1 _12356_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[15\].VALID\[11\].FF_D A[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XDATA\[0\].CLKBUF\[0\] clk vssd1 vssd1 vccd1 vccd1 _04967_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__05809__A _13902_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08830__D line[126] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11306_ _11306_/A _11339_/Y vssd1 vssd1 vccd1 vccd1 _13826_/Z sky130_fd_sc_hd__ebufn_2
X_12286_ _12286_/A _12319_/Y vssd1 vssd1 vccd1 vccd1 _13686_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_5_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13448__D line[61] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11237_ _11265_/CLK line[74] vssd1 vssd1 vccd1 vccd1 _11238_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05528__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07446__D line[119] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11168_ _11168_/A _11199_/Y vssd1 vssd1 vccd1 vccd1 _13688_/Z sky130_fd_sc_hd__ebufn_2
X_10119_ _10145_/CLK line[75] vssd1 vssd1 vccd1 vccd1 _10120_/A sky130_fd_sc_hd__dfxtp_1
X_11099_ _11125_/CLK line[11] vssd1 vssd1 vccd1 vccd1 _11100_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[25\].VALID\[10\].FF_D A[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10600__D line[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MUX.M\[0\].MUX\[6\]_A0 _13640_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05660_ _05660_/A _05669_/Y vssd1 vssd1 vccd1 vccd1 _13780_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07181__D line[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13809_ _13809_/A _13824_/Y vssd1 vssd1 vccd1 vccd1 _13809_/Z sky130_fd_sc_hd__ebufn_2
X_05591_ _05595_/CLK line[39] vssd1 vssd1 vccd1 vccd1 _05592_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_16_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07330_ _07330_/A _07349_/Y vssd1 vssd1 vccd1 vccd1 _13770_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[20\].CLKBUF\[4\] clk vssd1 vssd1 vccd1 vccd1 _08467_/CLK sky130_fd_sc_hd__clkbuf_4
X_07261_ _07275_/CLK line[34] vssd1 vssd1 vccd1 vccd1 _07262_/A sky130_fd_sc_hd__dfxtp_1
X_09000_ _09000_/A _09029_/Y vssd1 vssd1 vccd1 vccd1 _13760_/Z sky130_fd_sc_hd__ebufn_2
X_06212_ _06212_/A _06229_/Y vssd1 vssd1 vccd1 vccd1 _13772_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[24\].VALID\[7\].FF OVHB\[24\].V/CLK A[14] vssd1 vssd1 vccd1 vccd1 OVHB\[24\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_07192_ _07192_/A _07209_/Y vssd1 vssd1 vccd1 vccd1 _13632_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_176_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06143_ _06155_/CLK line[35] vssd1 vssd1 vccd1 vccd1 _06144_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10047__D line[42] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[16\].VALID\[2\].TOBUF OVHB\[16\].VALID\[2\].FF/Q OVHB\[16\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04930_/B2 sky130_fd_sc_hd__ebufn_2
X_06074_ _06074_/A _06089_/Y vssd1 vssd1 vccd1 vccd1 _13634_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[14\].CLKBUF\[6\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09902_ _09902_/CLK _09903_/X vssd1 vssd1 vccd1 vccd1 _09900_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__12262__D line[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05025_ _05035_/CLK line[36] vssd1 vssd1 vccd1 vccd1 _05026_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_116_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07356__D line[92] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06260__D line[89] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09833_ _13921_/X wr vssd1 vssd1 vccd1 vccd1 _09833_/X sky130_fd_sc_hd__and2_1
X_09764_ _13921_/X vssd1 vssd1 vccd1 vccd1 _09764_/Y sky130_fd_sc_hd__inv_2
X_06976_ _06976_/A _06999_/Y vssd1 vssd1 vccd1 vccd1 _13696_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09571__D line[66] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08715_ _08745_/CLK line[64] vssd1 vssd1 vccd1 vccd1 _08716_/A sky130_fd_sc_hd__dfxtp_1
X_05927_ _05945_/CLK line[79] vssd1 vssd1 vccd1 vccd1 _05928_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_73_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09695_ _09725_/CLK line[0] vssd1 vssd1 vccd1 vccd1 _09696_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_26_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10510__D line[126] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05858_ _05858_/A _05879_/Y vssd1 vssd1 vccd1 vccd1 _13698_/Z sky130_fd_sc_hd__ebufn_2
X_08646_ _08646_/A _08679_/Y vssd1 vssd1 vccd1 vccd1 _13686_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05604__D line[59] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_199_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08577_ _08605_/CLK line[10] vssd1 vssd1 vccd1 vccd1 _08578_/A sky130_fd_sc_hd__dfxtp_1
X_05789_ _05805_/CLK line[1] vssd1 vssd1 vccd1 vccd1 _05790_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07528_ _07528_/A _07559_/Y vssd1 vssd1 vccd1 vccd1 _13688_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_DATA\[7\].CLKBUF\[6\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07459_ _07485_/CLK line[11] vssd1 vssd1 vccd1 vccd1 _07460_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12437__D line[111] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10470_ _10470_/A _10499_/Y vssd1 vssd1 vccd1 vccd1 _13830_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06435__D line[41] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09129_ _09129_/A _09134_/Y vssd1 vssd1 vccd1 vccd1 _13889_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09746__D line[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12140_ _12140_/CLK line[89] vssd1 vssd1 vccd1 vccd1 _12141_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_190_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12071_ _12071_/A _12074_/Y vssd1 vssd1 vccd1 vccd1 _13751_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_151_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XOVHB\[22\].VALID\[9\].FF OVHB\[22\].V/CLK A[16] vssd1 vssd1 vccd1 vccd1 OVHB\[22\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06170__D line[62] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11022_ _11022_/CLK _11023_/X vssd1 vssd1 vccd1 vccd1 _11020_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_103_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XOVHB\[30\].VALID\[14\].FF OVHB\[30\].V/CLK A[21] vssd1 vssd1 vccd1 vccd1 OVHB\[30\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12900__D line[52] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[22\].VALID\[1\].TOBUF OVHB\[22\].VALID\[1\].FF/Q OVHB\[22\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04926_/B2 sky130_fd_sc_hd__ebufn_2
XOVHB\[15\].INV _13949_/X vssd1 vssd1 vccd1 vccd1 OVHB\[15\].INV/Y sky130_fd_sc_hd__inv_2
X_12973_ _12973_/A _12984_/Y vssd1 vssd1 vccd1 vccd1 _13813_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_206_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11924_ _11930_/CLK line[118] vssd1 vssd1 vccd1 vccd1 _11925_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08097__D line[47] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11855_ _11855_/A _11864_/Y vssd1 vssd1 vccd1 vccd1 _13815_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_72_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10806_ _10810_/CLK line[119] vssd1 vssd1 vccd1 vccd1 _10807_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_32_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11786_ _11790_/CLK line[55] vssd1 vssd1 vccd1 vccd1 _11787_/A sky130_fd_sc_hd__dfxtp_1
X_13525_ _13525_/A _13544_/Y vssd1 vssd1 vccd1 vccd1 _13805_/Z sky130_fd_sc_hd__ebufn_2
X_10737_ _10737_/A _10744_/Y vssd1 vssd1 vccd1 vccd1 _13817_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_186_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11251__D line[66] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06345__D line[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13456_ _13470_/CLK line[50] vssd1 vssd1 vccd1 vccd1 _13457_/A sky130_fd_sc_hd__dfxtp_1
X_10668_ _10670_/CLK line[56] vssd1 vssd1 vccd1 vccd1 _10669_/A sky130_fd_sc_hd__dfxtp_1
X_12407_ _12407_/A _12424_/Y vssd1 vssd1 vccd1 vccd1 _13807_/Z sky130_fd_sc_hd__ebufn_2
X_10599_ _10599_/A _10604_/Y vssd1 vssd1 vccd1 vccd1 _13679_/Z sky130_fd_sc_hd__ebufn_2
X_13387_ _13387_/A _13404_/Y vssd1 vssd1 vccd1 vccd1 _13667_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08560__D line[116] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12338_ _12350_/CLK line[51] vssd1 vssd1 vccd1 vccd1 _12339_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_99_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13178__D line[51] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12269_ _12269_/A _12284_/Y vssd1 vssd1 vccd1 vccd1 _13669_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[20\].VALID\[2\].FF_D A[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12810__D line[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06830_ _06830_/A _06859_/Y vssd1 vssd1 vccd1 vccd1 _13830_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_68_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06761_ _06785_/CLK line[76] vssd1 vssd1 vccd1 vccd1 _06762_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_55_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11426__D line[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08500_ _08500_/CLK line[89] vssd1 vssd1 vccd1 vccd1 _08501_/A sky130_fd_sc_hd__dfxtp_1
X_05712_ _05712_/A _05739_/Y vssd1 vssd1 vccd1 vccd1 _13832_/Z sky130_fd_sc_hd__ebufn_2
X_09480_ _09480_/CLK line[25] vssd1 vssd1 vccd1 vccd1 _09481_/A sky130_fd_sc_hd__dfxtp_1
X_06692_ _06692_/A _06719_/Y vssd1 vssd1 vccd1 vccd1 _13692_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[14\].VALID\[7\].TOBUF OVHB\[14\].VALID\[7\].FF/Q OVHB\[14\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/A2 sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[13\].VALID\[6\].FF_D A[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11723__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05643_ _05665_/CLK line[77] vssd1 vssd1 vccd1 vccd1 _05644_/A sky130_fd_sc_hd__dfxtp_1
X_08431_ _08431_/A _08434_/Y vssd1 vssd1 vccd1 vccd1 _13751_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_23_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13641__D line[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08362_ _08362_/CLK _08363_/X vssd1 vssd1 vccd1 vccd1 _08360_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__08735__D line[68] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05574_ _05574_/A _05599_/Y vssd1 vssd1 vccd1 vccd1 _13694_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_51_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07313_ _13910_/X wr vssd1 vssd1 vccd1 vccd1 _07313_/X sky130_fd_sc_hd__and2_1
X_08293_ _13932_/X wr vssd1 vssd1 vccd1 vccd1 _08293_/X sky130_fd_sc_hd__and2_1
XFILLER_165_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07244_ _13910_/X vssd1 vssd1 vccd1 vccd1 _07244_/Y sky130_fd_sc_hd__inv_2
XFILLER_177_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07175_ _07205_/CLK line[0] vssd1 vssd1 vccd1 vccd1 _07176_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[28\].CLKBUF\[0\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06126_ _06126_/A _06159_/Y vssd1 vssd1 vccd1 vccd1 _13686_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08470__D line[80] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[9\].VALID\[11\].TOBUF OVHB\[9\].VALID\[11\].FF/Q OVHB\[9\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04915_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_160_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06057_ _06085_/CLK line[10] vssd1 vssd1 vccd1 vccd1 _06058_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07086__D line[82] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05008_ _05008_/A _05039_/Y vssd1 vssd1 vccd1 vccd1 _13688_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_87_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07664__A _13911_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13816__D line[87] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09816_ _09830_/CLK line[50] vssd1 vssd1 vccd1 vccd1 _09817_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07383__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09747_ _09747_/A _09764_/Y vssd1 vssd1 vccd1 vccd1 _13667_/Z sky130_fd_sc_hd__ebufn_2
X_06959_ _06959_/A _06964_/Y vssd1 vssd1 vccd1 vccd1 _13679_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10240__D line[116] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09678_ _09690_/CLK line[115] vssd1 vssd1 vccd1 vccd1 _09679_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05334__D line[49] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08629_ _08629_/A _08644_/Y vssd1 vssd1 vccd1 vccd1 _13669_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_54_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13551__D line[108] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08645__D line[32] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11640_ _11650_/CLK line[116] vssd1 vssd1 vccd1 vccd1 _11641_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12167__D line[101] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11571_ _11571_/A _11584_/Y vssd1 vssd1 vccd1 vccd1 _13811_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[2\].VALID\[10\].TOBUF OVHB\[2\].VALID\[10\].FF/Q OVHB\[2\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04932_/B2 sky130_fd_sc_hd__ebufn_2
XPHY_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13310_ _13330_/CLK line[126] vssd1 vssd1 vccd1 vccd1 _13311_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07839__A _13912_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10522_ _10530_/CLK line[117] vssd1 vssd1 vccd1 vccd1 _10523_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[20\].VALID\[6\].TOBUF OVHB\[20\].VALID\[6\].FF/Q OVHB\[20\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04923_/A2 sky130_fd_sc_hd__ebufn_2
X_10453_ _10453_/A _10464_/Y vssd1 vssd1 vccd1 vccd1 _13813_/Z sky130_fd_sc_hd__ebufn_2
X_13241_ _13241_/A _13264_/Y vssd1 vssd1 vccd1 vccd1 _13801_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07558__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09476__D line[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MUX.M\[2\].MUX\[7\]_A2 _13817_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10384_ _10390_/CLK line[54] vssd1 vssd1 vccd1 vccd1 _10385_/A sky130_fd_sc_hd__dfxtp_1
X_13172_ _13190_/CLK line[63] vssd1 vssd1 vccd1 vccd1 _13173_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_123_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12123_ _12123_/A _12144_/Y vssd1 vssd1 vccd1 vccd1 _13803_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10415__D line[68] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05509__D line[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12054_ _12070_/CLK line[49] vssd1 vssd1 vccd1 vccd1 _12055_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13726__D line[60] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11005_ _11005_/A _11024_/Y vssd1 vssd1 vccd1 vccd1 _13805_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12630__D line[57] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07724__D line[118] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[26\].VALID\[6\].FF_D A[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10150__D line[80] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XOVHB\[13\].CG clk OVHB\[13\].CGAND/X vssd1 vssd1 vccd1 vccd1 OVHB\[13\].V/CLK sky130_fd_sc_hd__dlclkp_1
X_12956_ _12980_/CLK line[92] vssd1 vssd1 vccd1 vccd1 _12957_/A sky130_fd_sc_hd__dfxtp_1
X_11907_ _11907_/A _11934_/Y vssd1 vssd1 vccd1 vccd1 _13867_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_206_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12887_ _12887_/A _12914_/Y vssd1 vssd1 vccd1 vccd1 _13727_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.M\[0\].MUX\[3\]_A3 _13844_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11838_ _11860_/CLK line[93] vssd1 vssd1 vccd1 vccd1 _11839_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_61_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12077__D line[74] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11769_ _11769_/A _11794_/Y vssd1 vssd1 vccd1 vccd1 _13729_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06075__D line[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13508_ _13898_/Y wr vssd1 vssd1 vccd1 vccd1 _13508_/X sky130_fd_sc_hd__and2_1
X_05290_ _05290_/A _05319_/Y vssd1 vssd1 vccd1 vccd1 _13690_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_146_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12805__D line[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13439_ _13898_/Y vssd1 vssd1 vccd1 vccd1 _13439_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09386__D line[124] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08290__D line[121] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10325__D line[32] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08980_ _08990_/CLK line[52] vssd1 vssd1 vccd1 vccd1 _08981_/A sky130_fd_sc_hd__dfxtp_1
X_07931_ _07931_/A _07944_/Y vssd1 vssd1 vccd1 vccd1 _13811_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12540__D line[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07862_ _07870_/CLK line[53] vssd1 vssd1 vccd1 vccd1 _07863_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_3_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07634__D line[91] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09601_ _09601_/A _09624_/Y vssd1 vssd1 vccd1 vccd1 _13801_/Z sky130_fd_sc_hd__ebufn_2
X_06813_ _06813_/A _06824_/Y vssd1 vssd1 vccd1 vccd1 _13813_/Z sky130_fd_sc_hd__ebufn_2
X_07793_ _07793_/A _07804_/Y vssd1 vssd1 vccd1 vccd1 _13673_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11156__D line[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09532_ _09550_/CLK line[63] vssd1 vssd1 vccd1 vccd1 _09533_/A sky130_fd_sc_hd__dfxtp_1
X_06744_ _06750_/CLK line[54] vssd1 vssd1 vccd1 vccd1 _06745_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[29\].VALID\[1\].TOBUF OVHB\[29\].VALID\[1\].FF/Q OVHB\[29\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04926_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__09204__A _13916_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06675_ _06675_/A _06684_/Y vssd1 vssd1 vccd1 vccd1 _13675_/Z sky130_fd_sc_hd__ebufn_2
X_09463_ _09463_/A _09484_/Y vssd1 vssd1 vccd1 vccd1 _13663_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_64_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08414_ _08430_/CLK line[49] vssd1 vssd1 vccd1 vccd1 _08415_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08465__D line[73] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05626_ _05630_/CLK line[55] vssd1 vssd1 vccd1 vccd1 _05627_/A sky130_fd_sc_hd__dfxtp_1
X_09394_ _09410_/CLK line[113] vssd1 vssd1 vccd1 vccd1 _09395_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_24_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05557_ _05557_/A _05564_/Y vssd1 vssd1 vccd1 vccd1 _13677_/Z sky130_fd_sc_hd__ebufn_2
X_08345_ _08345_/A _08364_/Y vssd1 vssd1 vccd1 vccd1 _13665_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_177_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08276_ _08290_/CLK line[114] vssd1 vssd1 vccd1 vccd1 _08277_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_20_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05488_ _05490_/CLK line[120] vssd1 vssd1 vccd1 vccd1 _05489_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[7\].VALID\[1\].FF_D A[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12715__D line[110] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07227_ _07227_/A _07244_/Y vssd1 vssd1 vccd1 vccd1 _13667_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[25\].VALID\[12\].TOBUF OVHB\[25\].VALID\[12\].FF/Q OVHB\[25\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04929_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__07809__D line[43] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05179__A _13931_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07158_ _07170_/CLK line[115] vssd1 vssd1 vccd1 vccd1 _07159_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06713__D line[40] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06109_ _06109_/A _06124_/Y vssd1 vssd1 vccd1 vccd1 _13669_/Z sky130_fd_sc_hd__ebufn_2
X_07089_ _07089_/A _07104_/Y vssd1 vssd1 vccd1 vccd1 _13809_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10813__A _13924_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[26\].CLKBUF\[2\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11066__D line[124] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12810_ _12840_/CLK line[16] vssd1 vssd1 vccd1 vccd1 _12811_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_90_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13790_ _13820_/CLK line[80] vssd1 vssd1 vccd1 vccd1 _13791_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_43_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05064__D line[54] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12741_ _12741_/A _12774_/Y vssd1 vssd1 vccd1 vccd1 _13861_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[8\].CG clk OVHB\[8\].CGAND/X vssd1 vssd1 vccd1 vccd1 OVHB\[8\].V/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__13281__D line[98] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05999__D line[97] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08375__D line[46] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12672_ _12700_/CLK line[90] vssd1 vssd1 vccd1 vccd1 _12673_/A sky130_fd_sc_hd__dfxtp_1
XPHY_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11623_ _11623_/A _11654_/Y vssd1 vssd1 vccd1 vccd1 _13863_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11554_ _11580_/CLK line[91] vssd1 vssd1 vccd1 vccd1 _11555_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06473__A _13904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10505_ _10505_/A _10534_/Y vssd1 vssd1 vccd1 vccd1 _13865_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_195_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11485_ _11485_/A _11514_/Y vssd1 vssd1 vccd1 vccd1 _13725_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06623__D line[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13224_ _13224_/A _13229_/Y vssd1 vssd1 vccd1 vccd1 _13784_/Z sky130_fd_sc_hd__ebufn_2
X_10436_ _10460_/CLK line[92] vssd1 vssd1 vccd1 vccd1 _10437_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_136_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10145__D line[73] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13155_ _13155_/CLK line[41] vssd1 vssd1 vccd1 vccd1 _13156_/A sky130_fd_sc_hd__dfxtp_1
X_10367_ _10367_/A _10394_/Y vssd1 vssd1 vccd1 vccd1 _13727_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05239__D line[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12106_ _12106_/A _12109_/Y vssd1 vssd1 vccd1 vccd1 _13786_/Z sky130_fd_sc_hd__ebufn_2
X_13086_ _13086_/A _13089_/Y vssd1 vssd1 vccd1 vccd1 _13646_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_2_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10298_ _10320_/CLK line[29] vssd1 vssd1 vccd1 vccd1 _10299_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13456__D line[50] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12037_ _12037_/CLK _12038_/X vssd1 vssd1 vccd1 vccd1 _12035_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__13753__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06648__A _13905_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12939_ _12945_/CLK line[70] vssd1 vssd1 vccd1 vccd1 _12940_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_80_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11704__D line[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06460_ _06470_/CLK line[52] vssd1 vssd1 vccd1 vccd1 _06461_/A sky130_fd_sc_hd__dfxtp_1
X_05411_ _05411_/A _05424_/Y vssd1 vssd1 vccd1 vccd1 _13811_/Z sky130_fd_sc_hd__ebufn_2
X_06391_ _06391_/A _06404_/Y vssd1 vssd1 vccd1 vccd1 _13671_/Z sky130_fd_sc_hd__ebufn_2
X_08130_ _08150_/CLK line[62] vssd1 vssd1 vccd1 vccd1 _08131_/A sky130_fd_sc_hd__dfxtp_1
X_05342_ _05350_/CLK line[53] vssd1 vssd1 vccd1 vccd1 _05343_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_186_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08061_ _08061_/A _08084_/Y vssd1 vssd1 vccd1 vccd1 _13661_/Z sky130_fd_sc_hd__ebufn_2
X_05273_ _05273_/A _05284_/Y vssd1 vssd1 vccd1 vccd1 _13673_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[2\].VALID\[3\].TOBUF OVHB\[2\].VALID\[3\].FF/Q OVHB\[2\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04919_/B2 sky130_fd_sc_hd__ebufn_2
X_07012_ _07030_/CLK line[63] vssd1 vssd1 vccd1 vccd1 _07013_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09694__A _13920_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[0\].VALID\[14\].FF_D A[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[27\].VALID\[6\].TOBUF OVHB\[27\].VALID\[6\].FF/Q OVHB\[27\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04923_/A2 sky130_fd_sc_hd__ebufn_2
XANTENNA__10055__D line[46] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05149__D line[107] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08963_ _08963_/A _08994_/Y vssd1 vssd1 vccd1 vccd1 _13723_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12270__D line[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__04988__D line[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07914_ _07940_/CLK line[91] vssd1 vssd1 vccd1 vccd1 _07915_/A sky130_fd_sc_hd__dfxtp_1
X_08894_ _08920_/CLK line[27] vssd1 vssd1 vccd1 vccd1 _08895_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_84_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07364__D line[81] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07845_ _07845_/A _07874_/Y vssd1 vssd1 vccd1 vccd1 _13725_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_56_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[10\].CGAND _13900_/X wr vssd1 vssd1 vccd1 vccd1 OVHB\[10\].CGAND/X sky130_fd_sc_hd__and2_4
X_07776_ _07800_/CLK line[28] vssd1 vssd1 vccd1 vccd1 _07777_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_72_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_04988_ _05000_/CLK line[19] vssd1 vssd1 vccd1 vccd1 _04989_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_37_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09515_ _09515_/CLK line[41] vssd1 vssd1 vccd1 vccd1 _09516_/A sky130_fd_sc_hd__dfxtp_1
X_06727_ _06727_/A _06754_/Y vssd1 vssd1 vccd1 vccd1 _13727_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_25_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09446_ _09446_/A _09449_/Y vssd1 vssd1 vccd1 vccd1 _13646_/Z sky130_fd_sc_hd__ebufn_2
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09869__A _13921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06658_ _06680_/CLK line[29] vssd1 vssd1 vccd1 vccd1 _06659_/A sky130_fd_sc_hd__dfxtp_1
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05612__D line[63] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05609_ _05609_/A _05634_/Y vssd1 vssd1 vccd1 vccd1 _13729_/Z sky130_fd_sc_hd__ebufn_2
X_09377_ _09377_/CLK _09378_/X vssd1 vssd1 vccd1 vccd1 _09375_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_185_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09588__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06589_ _06589_/A _06614_/Y vssd1 vssd1 vccd1 vccd1 _13869_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_178_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08328_ _13913_/X wr vssd1 vssd1 vccd1 vccd1 _08328_/X sky130_fd_sc_hd__and2_1
XANTENNA__12445__D line[100] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08259_ _13932_/X vssd1 vssd1 vccd1 vccd1 _08259_/Y sky130_fd_sc_hd__inv_2
XANTENNA__07539__D line[33] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11270_ _11300_/CLK line[80] vssd1 vssd1 vccd1 vccd1 _11271_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_192_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10221_ _10221_/A _10254_/Y vssd1 vssd1 vccd1 vccd1 _13861_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_165_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[8\].VALID\[9\].FF OVHB\[8\].V/CLK A[16] vssd1 vssd1 vccd1 vccd1 OVHB\[8\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_133_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09754__D line[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10152_ _10180_/CLK line[90] vssd1 vssd1 vccd1 vccd1 _10153_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08013__A _13912_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12180__D line[112] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10083_ _10083_/A _10114_/Y vssd1 vssd1 vccd1 vccd1 _13723_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_94_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_OVHB\[22\].VALID\[9\].FF_D A[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13911_ _13916_/C _13916_/A _13916_/B _13916_/D vssd1 vssd1 vccd1 vccd1 _13911_/X
+ sky130_fd_sc_hd__and4bb_4
XFILLER_101_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11374__A _13933_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13842_ _13842_/A _13859_/Y vssd1 vssd1 vccd1 vccd1 _13842_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_16_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11093__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13773_ _13785_/CLK line[67] vssd1 vssd1 vccd1 vccd1 _13774_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[24\].CLKBUF\[4\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10985_ _10985_/CLK line[73] vssd1 vssd1 vccd1 vccd1 _10986_/A sky130_fd_sc_hd__dfxtp_1
X_12724_ _12724_/A _12739_/Y vssd1 vssd1 vccd1 vccd1 _13844_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[2\].VALID\[10\].FF_D A[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12655_ _12665_/CLK line[68] vssd1 vssd1 vccd1 vccd1 _12656_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09929__D line[102] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11606_ _11606_/A _11619_/Y vssd1 vssd1 vccd1 vccd1 _13846_/Z sky130_fd_sc_hd__ebufn_2
XPHY_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[12\].CG_CLK clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12586_ _12586_/A _12599_/Y vssd1 vssd1 vccd1 vccd1 _13706_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12355__D line[64] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11537_ _11545_/CLK line[69] vssd1 vssd1 vccd1 vccd1 _11538_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_7_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06353__D line[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11468_ _11468_/A _11479_/Y vssd1 vssd1 vccd1 vccd1 _13708_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_125_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11549__A _13926_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13207_ _13225_/CLK line[79] vssd1 vssd1 vccd1 vccd1 _13208_/A sky130_fd_sc_hd__dfxtp_1
X_10419_ _10425_/CLK line[70] vssd1 vssd1 vccd1 vccd1 _10420_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[24\].V_RESET_B rst_n vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11399_ _11405_/CLK line[6] vssd1 vssd1 vccd1 vccd1 _11400_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09664__D line[123] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11268__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13138_ _13138_/A _13159_/Y vssd1 vssd1 vccd1 vccd1 _13698_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13186__D line[55] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13069_ _13085_/CLK line[1] vssd1 vssd1 vccd1 vccd1 _13070_/A sky130_fd_sc_hd__dfxtp_1
X_05960_ _05980_/CLK line[94] vssd1 vssd1 vccd1 vccd1 _05961_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_04911_ A_h[14] vssd1 vssd1 vccd1 vccd1 _04911_/Y sky130_fd_sc_hd__inv_2
X_05891_ _05891_/A _05914_/Y vssd1 vssd1 vccd1 vccd1 _13731_/Z sky130_fd_sc_hd__ebufn_2
X_07630_ _07660_/CLK line[80] vssd1 vssd1 vccd1 vccd1 _07631_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_54_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07912__D line[90] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[0\].VALID\[8\].TOBUF OVHB\[0\].VALID\[8\].FF/Q OVHB\[0\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04931_/B2 sky130_fd_sc_hd__ebufn_2
X_07561_ _07561_/A _07594_/Y vssd1 vssd1 vccd1 vccd1 _13721_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_46_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11434__D line[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09300_ _09300_/A _09309_/Y vssd1 vssd1 vccd1 vccd1 _13780_/Z sky130_fd_sc_hd__ebufn_2
X_06512_ _06540_/CLK line[90] vssd1 vssd1 vccd1 vccd1 _06513_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_80_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06528__D line[83] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07492_ _07520_/CLK line[26] vssd1 vssd1 vccd1 vccd1 _07493_/A sky130_fd_sc_hd__dfxtp_1
X_09231_ _09235_/CLK line[39] vssd1 vssd1 vccd1 vccd1 _09232_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_167_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06443_ _06443_/A _06474_/Y vssd1 vssd1 vccd1 vccd1 _13723_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[3\].VALID\[4\].FF_D A[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09839__D line[75] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09162_ _09162_/A _09169_/Y vssd1 vssd1 vccd1 vccd1 _13642_/Z sky130_fd_sc_hd__ebufn_2
X_06374_ _06400_/CLK line[27] vssd1 vssd1 vccd1 vccd1 _06375_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_9_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08743__D line[72] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05325_ _05325_/A _05354_/Y vssd1 vssd1 vccd1 vccd1 _13725_/Z sky130_fd_sc_hd__ebufn_2
X_08113_ _08115_/CLK line[40] vssd1 vssd1 vccd1 vccd1 _08114_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_119_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13939__A A_h[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09093_ _09095_/CLK line[104] vssd1 vssd1 vccd1 vccd1 _09094_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12843__A _13937_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08044_ _08044_/A _08049_/Y vssd1 vssd1 vccd1 vccd1 _13644_/Z sky130_fd_sc_hd__ebufn_2
X_05256_ _05280_/CLK line[28] vssd1 vssd1 vccd1 vccd1 _05257_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_134_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05187_ _05187_/A _05214_/Y vssd1 vssd1 vccd1 vccd1 _13867_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_135_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XOVHB\[17\].VALID\[1\].FF OVHB\[17\].V/CLK A[8] vssd1 vssd1 vccd1 vccd1 OVHB\[17\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_09995_ _10005_/CLK line[4] vssd1 vssd1 vccd1 vccd1 _09996_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_142_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13096__D line[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11609__D line[102] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08946_ _08946_/A _08959_/Y vssd1 vssd1 vccd1 vccd1 _13706_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[4\].VOBUF OVHB\[4\].V/Q OVHB\[4\].INV/Y vssd1 vssd1 vccd1 vccd1 _04912_/B1
+ sky130_fd_sc_hd__ebufn_2
XFILLER_88_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07094__D line[86] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08877_ _08885_/CLK line[5] vssd1 vssd1 vccd1 vccd1 _08878_/A sky130_fd_sc_hd__dfxtp_1
X_07828_ _07828_/A _07839_/Y vssd1 vssd1 vccd1 vccd1 _13708_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08918__D line[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07759_ _07765_/CLK line[6] vssd1 vssd1 vccd1 vccd1 _07760_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11344__D line[123] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10770_ _10770_/A _10779_/Y vssd1 vssd1 vccd1 vccd1 _13850_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05342__D line[53] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09429_ _09445_/CLK line[1] vssd1 vssd1 vccd1 vccd1 _09430_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_201_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08653__D line[45] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12440_ _12440_/A _12459_/Y vssd1 vssd1 vccd1 vccd1 _13840_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_138_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XOVHB\[15\].VALID\[10\].TOBUF OVHB\[15\].VALID\[10\].FF/Q OVHB\[15\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04932_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__12175__D line[105] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12371_ _12385_/CLK line[66] vssd1 vssd1 vccd1 vccd1 _12372_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07269__D line[38] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11322_ _11322_/A _11339_/Y vssd1 vssd1 vccd1 vccd1 _13842_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_153_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11253_ _11265_/CLK line[67] vssd1 vssd1 vccd1 vccd1 _11254_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[18\].VALID\[1\].FF_D A[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[9\].VALID\[3\].TOBUF OVHB\[9\].VALID\[3\].FF/Q OVHB\[9\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04919_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_180_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10204_ _10204_/A _10219_/Y vssd1 vssd1 vccd1 vccd1 _13844_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06901__D line[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11184_ _11184_/A _11199_/Y vssd1 vssd1 vccd1 vccd1 _13704_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[7\].VALID\[14\].FF_D A[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11519__D line[75] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10423__D line[72] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10135_ _10145_/CLK line[68] vssd1 vssd1 vccd1 vccd1 _10136_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05517__D line[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08678__A _13914_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_MUX.M\[1\].MUX\[5\]_A3 _13834_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10066_ _10066_/A _10079_/Y vssd1 vssd1 vccd1 vccd1 _13706_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_208_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13734__D line[49] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08828__D line[125] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XOVHB\[15\].VALID\[3\].FF OVHB\[15\].V/CLK A[10] vssd1 vssd1 vccd1 vccd1 OVHB\[15\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_13825_ _13855_/CLK line[96] vssd1 vssd1 vccd1 vccd1 _13826_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_90_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13756_ _13756_/A _13789_/Y vssd1 vssd1 vccd1 vccd1 _13756_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05252__D line[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10968_ _10968_/A _10989_/Y vssd1 vssd1 vccd1 vccd1 _13768_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_203_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12707_ _12735_/CLK line[106] vssd1 vssd1 vccd1 vccd1 _12708_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_43_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XOVHB\[31\].VALID\[12\].FF OVHB\[31\].V/CLK A[19] vssd1 vssd1 vccd1 vccd1 OVHB\[31\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_13687_ _13715_/CLK line[42] vssd1 vssd1 vccd1 vccd1 _13688_/A sky130_fd_sc_hd__dfxtp_1
X_10899_ _10915_/CLK line[33] vssd1 vssd1 vccd1 vccd1 _10900_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_176_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12638_ _12638_/A _12669_/Y vssd1 vssd1 vccd1 vccd1 _13758_/Z sky130_fd_sc_hd__ebufn_2
XPHY_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_DATA\[22\].CLKBUF\[6\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12085__D line[78] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12569_ _12595_/CLK line[43] vssd1 vssd1 vccd1 vccd1 _12570_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[9\].VALID\[8\].FF_D A[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07179__D line[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05110_ _05140_/CLK line[80] vssd1 vssd1 vccd1 vccd1 _05111_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06083__D line[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06090_ _06120_/CLK line[16] vssd1 vssd1 vccd1 vccd1 _06091_/A sky130_fd_sc_hd__dfxtp_1
X_05041_ _05041_/A _05074_/Y vssd1 vssd1 vccd1 vccd1 _13721_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10183__A _13922_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09394__D line[113] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08800_ _08800_/A _08819_/Y vssd1 vssd1 vccd1 vccd1 _13840_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10333__D line[45] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09780_ _09780_/A _09799_/Y vssd1 vssd1 vccd1 vccd1 _13700_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_112_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06992_ _06992_/A _06999_/Y vssd1 vssd1 vccd1 vccd1 _13712_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05427__D line[106] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__04919__A1_N A_h[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08731_ _08745_/CLK line[66] vssd1 vssd1 vccd1 vccd1 _08732_/A sky130_fd_sc_hd__dfxtp_1
X_05943_ _05945_/CLK line[72] vssd1 vssd1 vccd1 vccd1 _05944_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[21\].VALID\[14\].FF OVHB\[21\].V/CLK A[21] vssd1 vssd1 vccd1 vccd1 OVHB\[21\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_08662_ _08662_/A _08679_/Y vssd1 vssd1 vccd1 vccd1 _13702_/Z sky130_fd_sc_hd__ebufn_2
X_05874_ _05874_/A _05879_/Y vssd1 vssd1 vccd1 vccd1 _13714_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07642__D line[95] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07613_ _07625_/CLK line[67] vssd1 vssd1 vccd1 vccd1 _07614_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08593_ _08605_/CLK line[3] vssd1 vssd1 vccd1 vccd1 _08594_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_121_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07544_ _07544_/A _07559_/Y vssd1 vssd1 vccd1 vccd1 _13704_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06258__D line[88] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07475_ _07485_/CLK line[4] vssd1 vssd1 vccd1 vccd1 _07476_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10358__A _13923_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09569__D line[65] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09214_ _09214_/A _09239_/Y vssd1 vssd1 vccd1 vccd1 _13694_/Z sky130_fd_sc_hd__ebufn_2
X_06426_ _06426_/A _06439_/Y vssd1 vssd1 vccd1 vccd1 _13706_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[9\].VALID\[10\].FF_D A[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[13\].VALID\[5\].FF OVHB\[13\].V/CLK A[12] vssd1 vssd1 vccd1 vccd1 OVHB\[13\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_09145_ _09165_/CLK line[14] vssd1 vssd1 vccd1 vccd1 _09146_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10508__D line[125] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[30\].VALID\[9\].FF OVHB\[30\].V/CLK A[16] vssd1 vssd1 vccd1 vccd1 OVHB\[30\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_06357_ _06365_/CLK line[5] vssd1 vssd1 vccd1 vccd1 _06358_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_175_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05308_ _05308_/A _05319_/Y vssd1 vssd1 vccd1 vccd1 _13708_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_107_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09076_ _09076_/A _09099_/Y vssd1 vssd1 vccd1 vccd1 _13836_/Z sky130_fd_sc_hd__ebufn_2
X_06288_ _06288_/A _06299_/Y vssd1 vssd1 vccd1 vccd1 _13848_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_190_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12723__D line[99] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08027_ _08045_/CLK line[15] vssd1 vssd1 vccd1 vccd1 _08028_/A sky130_fd_sc_hd__dfxtp_1
X_05239_ _05245_/CLK line[6] vssd1 vssd1 vccd1 vccd1 _05240_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07817__D line[47] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09978_ _09978_/A _10009_/Y vssd1 vssd1 vccd1 vccd1 _13618_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_131_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08929_ _08955_/CLK line[43] vssd1 vssd1 vccd1 vccd1 _08930_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_69_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11940_ _11940_/A _11969_/Y vssd1 vssd1 vccd1 vccd1 _13620_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_18_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11871_ _11895_/CLK line[108] vssd1 vssd1 vccd1 vccd1 _11872_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_44_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11074__D line[113] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13610_ _13610_/CLK line[121] vssd1 vssd1 vccd1 vccd1 _13611_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_55_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10822_ _10822_/A _10849_/Y vssd1 vssd1 vccd1 vccd1 _13622_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06168__D line[61] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[7\].VALID\[8\].TOBUF OVHB\[7\].VALID\[8\].FF/Q OVHB\[7\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04931_/B2 sky130_fd_sc_hd__ebufn_2
X_13541_ _13541_/A _13544_/Y vssd1 vssd1 vccd1 vccd1 _13821_/Z sky130_fd_sc_hd__ebufn_2
X_10753_ _10775_/CLK line[109] vssd1 vssd1 vccd1 vccd1 _10754_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DECH.DEC0.AND2_B A_h[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08383__D line[35] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13472_ _13472_/CLK _13473_/X vssd1 vssd1 vccd1 vccd1 _13470_/CLK sky130_fd_sc_hd__dlclkp_1
X_10684_ _10684_/A _10709_/Y vssd1 vssd1 vccd1 vccd1 _13764_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_187_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13579__A _13898_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12423_ _13935_/X wr vssd1 vssd1 vccd1 vccd1 _12423_/X sky130_fd_sc_hd__and2_1
XFILLER_138_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12354_ _13935_/X vssd1 vssd1 vccd1 vccd1 _12354_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13298__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11305_ _11335_/CLK line[96] vssd1 vssd1 vccd1 vccd1 _11306_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12285_ _12315_/CLK line[32] vssd1 vssd1 vccd1 vccd1 _12286_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[11\].VALID\[7\].FF OVHB\[11\].V/CLK A[14] vssd1 vssd1 vccd1 vccd1 OVHB\[11\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06631__D line[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11236_ _11236_/A _11269_/Y vssd1 vssd1 vccd1 vccd1 _13756_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11249__D line[65] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11167_ _11195_/CLK line[42] vssd1 vssd1 vccd1 vccd1 _11168_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09942__D line[122] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10118_ _10118_/A _10149_/Y vssd1 vssd1 vccd1 vccd1 _13758_/Z sky130_fd_sc_hd__ebufn_2
X_11098_ _11098_/A _11129_/Y vssd1 vssd1 vccd1 vccd1 _13618_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_95_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13464__D line[54] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10049_ _10075_/CLK line[43] vssd1 vssd1 vccd1 vccd1 _10050_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08558__D line[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MUX.M\[0\].MUX\[6\]_A1 _13710_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05590_ _05590_/A _05599_/Y vssd1 vssd1 vccd1 vccd1 _13710_/Z sky130_fd_sc_hd__ebufn_2
X_13808_ _13820_/CLK line[83] vssd1 vssd1 vccd1 vccd1 _13809_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_204_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13739_ _13739_/A _13754_/Y vssd1 vssd1 vccd1 vccd1 _13739_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11712__D line[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07260_ _07260_/A _07279_/Y vssd1 vssd1 vccd1 vccd1 _13700_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06806__D line[82] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06211_ _06225_/CLK line[66] vssd1 vssd1 vccd1 vccd1 _06212_/A sky130_fd_sc_hd__dfxtp_1
X_07191_ _07205_/CLK line[2] vssd1 vssd1 vccd1 vccd1 _07192_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_157_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06142_ _06142_/A _06159_/Y vssd1 vssd1 vccd1 vccd1 _13702_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_129_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13639__D line[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDATA\[19\].CLKBUF\[2\] clk vssd1 vssd1 vccd1 vccd1 _07837_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_105_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06073_ _06085_/CLK line[3] vssd1 vssd1 vccd1 vccd1 _06074_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[14\].VALID\[3\].TOBUF OVHB\[14\].VALID\[3\].FF/Q OVHB\[14\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04919_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_144_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09901_ _09901_/A _09904_/Y vssd1 vssd1 vccd1 vccd1 _13821_/Z sky130_fd_sc_hd__ebufn_2
X_05024_ _05024_/A _05039_/Y vssd1 vssd1 vccd1 vccd1 _13704_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_132_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XDEC.DEC0.AND0 A[5] A[6] vssd1 vssd1 vccd1 vccd1 _13938_/D sky130_fd_sc_hd__nor2_2
XANTENNA__10063__D line[35] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09832_ _09832_/CLK _09833_/X vssd1 vssd1 vccd1 vccd1 _09830_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_101_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05157__D line[111] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09763_ _13921_/X wr vssd1 vssd1 vccd1 vccd1 _09763_/X sky130_fd_sc_hd__and2_1
XANTENNA__10998__D line[93] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06975_ _06995_/CLK line[46] vssd1 vssd1 vccd1 vccd1 _06976_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13374__D line[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__04996__D line[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08714_ _13914_/X vssd1 vssd1 vccd1 vccd1 _08714_/Y sky130_fd_sc_hd__inv_2
XFILLER_132_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13952__A A_h[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05926_ _05926_/A _05949_/Y vssd1 vssd1 vccd1 vccd1 _13766_/Z sky130_fd_sc_hd__ebufn_2
X_09694_ _13920_/Y vssd1 vssd1 vccd1 vccd1 _09694_/Y sky130_fd_sc_hd__inv_2
XANTENNA__07372__D line[85] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08645_ _08675_/CLK line[32] vssd1 vssd1 vccd1 vccd1 _08646_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_26_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05857_ _05875_/CLK line[47] vssd1 vssd1 vccd1 vccd1 _05858_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08576_ _08576_/A _08609_/Y vssd1 vssd1 vccd1 vccd1 _13616_/Z sky130_fd_sc_hd__ebufn_2
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05788_ _05788_/A _05809_/Y vssd1 vssd1 vccd1 vccd1 _13628_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[21\].VALID\[0\].FF_D A[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07527_ _07555_/CLK line[42] vssd1 vssd1 vccd1 vccd1 _07528_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11622__D line[122] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09299__D line[70] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07458_ _07458_/A _07489_/Y vssd1 vssd1 vccd1 vccd1 _13618_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05620__D line[52] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10238__D line[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06409_ _06435_/CLK line[43] vssd1 vssd1 vccd1 vccd1 _06410_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_210_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07389_ _07415_/CLK line[107] vssd1 vssd1 vccd1 vccd1 _07390_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[14\].VALID\[4\].FF_D A[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09128_ _09130_/CLK line[120] vssd1 vssd1 vccd1 vccd1 _09129_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08931__D line[44] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13549__D line[107] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12453__D line[104] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09059_ _09059_/A _09064_/Y vssd1 vssd1 vccd1 vccd1 _13819_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_2_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07547__D line[37] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12070_ _12070_/CLK line[57] vssd1 vssd1 vccd1 vccd1 _12071_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_173_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11021_ _11021_/A _11024_/Y vssd1 vssd1 vccd1 vccd1 _13821_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_89_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10701__D line[71] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[20\].VALID\[2\].TOBUF OVHB\[20\].VALID\[2\].FF/Q OVHB\[20\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04930_/B2 sky130_fd_sc_hd__ebufn_2
X_12972_ _12980_/CLK line[85] vssd1 vssd1 vccd1 vccd1 _12973_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07282__D line[58] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11923_ _11923_/A _11934_/Y vssd1 vssd1 vccd1 vccd1 _13883_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_122_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11854_ _11860_/CLK line[86] vssd1 vssd1 vccd1 vccd1 _11855_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_82_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10805_ _10805_/A _10814_/Y vssd1 vssd1 vccd1 vccd1 _13885_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12628__D line[56] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11785_ _11785_/A _11794_/Y vssd1 vssd1 vccd1 vccd1 _13745_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_13_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13524_ _13540_/CLK line[81] vssd1 vssd1 vccd1 vccd1 _13525_/A sky130_fd_sc_hd__dfxtp_1
X_10736_ _10740_/CLK line[87] vssd1 vssd1 vccd1 vccd1 _10737_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_41_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05530__D line[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13455_ _13455_/A _13474_/Y vssd1 vssd1 vccd1 vccd1 _13735_/Z sky130_fd_sc_hd__ebufn_2
X_10667_ _10667_/A _10674_/Y vssd1 vssd1 vccd1 vccd1 _13747_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[10\].V_D TIE/HI vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12406_ _12420_/CLK line[82] vssd1 vssd1 vccd1 vccd1 _12407_/A sky130_fd_sc_hd__dfxtp_1
X_13386_ _13400_/CLK line[18] vssd1 vssd1 vccd1 vccd1 _13387_/A sky130_fd_sc_hd__dfxtp_1
X_10598_ _10600_/CLK line[24] vssd1 vssd1 vccd1 vccd1 _10599_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_154_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12363__D line[77] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12337_ _12337_/A _12354_/Y vssd1 vssd1 vccd1 vccd1 _13737_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07457__D line[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06361__D line[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12268_ _12280_/CLK line[19] vssd1 vssd1 vccd1 vccd1 _12269_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[25\].V_D TIE/HI vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[4\].VALID\[0\].FF OVHB\[4\].V/CLK A[7] vssd1 vssd1 vccd1 vccd1 OVHB\[4\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[15\].CLKBUF\[0\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11219_ _11219_/A _11234_/Y vssd1 vssd1 vccd1 vccd1 _13739_/Z sky130_fd_sc_hd__ebufn_2
X_12199_ _12199_/A _12214_/Y vssd1 vssd1 vccd1 vccd1 _13879_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_150_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09672__D line[127] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10611__D line[44] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06760_ _06760_/A _06789_/Y vssd1 vssd1 vccd1 vccd1 _13760_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08288__D line[120] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05705__D line[96] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05711_ _05735_/CLK line[108] vssd1 vssd1 vccd1 vccd1 _05712_/A sky130_fd_sc_hd__dfxtp_1
X_06691_ _06715_/CLK line[44] vssd1 vssd1 vccd1 vccd1 _06692_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12388__A _13935_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08430_ _08430_/CLK line[57] vssd1 vssd1 vccd1 vccd1 _08431_/A sky130_fd_sc_hd__dfxtp_1
X_05642_ _05642_/A _05669_/Y vssd1 vssd1 vccd1 vccd1 _13762_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[12\].VALID\[8\].TOBUF OVHB\[12\].VALID\[8\].FF/Q OVHB\[12\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04931_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__07920__D line[94] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12538__D line[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08361_ _08361_/A _08364_/Y vssd1 vssd1 vccd1 vccd1 _13681_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_16_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05573_ _05595_/CLK line[45] vssd1 vssd1 vccd1 vccd1 _05574_/A sky130_fd_sc_hd__dfxtp_1
X_07312_ _07312_/CLK _07313_/X vssd1 vssd1 vccd1 vccd1 _07310_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__06536__D line[87] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08292_ _08292_/CLK _08293_/X vssd1 vssd1 vccd1 vccd1 _08290_/CLK sky130_fd_sc_hd__dlclkp_1
XOVHB\[5\].VALID\[12\].TOBUF OVHB\[5\].VALID\[12\].FF/Q OVHB\[5\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04929_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[8\].CLKBUF\[0\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[27\].VALID\[4\].FF_D A[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07243_ _13910_/X wr vssd1 vssd1 vccd1 vccd1 _07243_/X sky130_fd_sc_hd__and2_1
XANTENNA__09847__D line[79] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07174_ _13909_/Y vssd1 vssd1 vccd1 vccd1 _07174_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06125_ _06155_/CLK line[32] vssd1 vssd1 vccd1 vccd1 _06126_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_127_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06271__D line[108] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06056_ _06056_/A _06089_/Y vssd1 vssd1 vccd1 vccd1 _13616_/Z sky130_fd_sc_hd__ebufn_2
X_05007_ _05035_/CLK line[42] vssd1 vssd1 vccd1 vccd1 _05008_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_143_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09815_ _09815_/A _09834_/Y vssd1 vssd1 vccd1 vccd1 _13735_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_101_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09746_ _09760_/CLK line[18] vssd1 vssd1 vccd1 vccd1 _09747_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08198__D line[93] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06958_ _06960_/CLK line[24] vssd1 vssd1 vccd1 vccd1 _06959_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_67_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05909_ _05909_/A _05914_/Y vssd1 vssd1 vccd1 vccd1 _13749_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[2\].VALID\[2\].FF OVHB\[2\].V/CLK A[9] vssd1 vssd1 vccd1 vccd1 OVHB\[2\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_09677_ _09677_/A _09694_/Y vssd1 vssd1 vccd1 vccd1 _13877_/Z sky130_fd_sc_hd__ebufn_2
X_06889_ _06889_/A _06894_/Y vssd1 vssd1 vccd1 vccd1 _13889_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_199_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08628_ _08640_/CLK line[19] vssd1 vssd1 vccd1 vccd1 _08629_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_15_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08559_ _08559_/A _08574_/Y vssd1 vssd1 vccd1 vccd1 _13879_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11352__D line[127] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06446__D line[60] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11570_ _11580_/CLK line[84] vssd1 vssd1 vccd1 vccd1 _11571_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05350__D line[57] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10521_ _10521_/A _10534_/Y vssd1 vssd1 vccd1 vccd1 _13881_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_7_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08661__D line[34] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13240_ _13260_/CLK line[94] vssd1 vssd1 vccd1 vccd1 _13241_/A sky130_fd_sc_hd__dfxtp_1
X_10452_ _10460_/CLK line[85] vssd1 vssd1 vccd1 vccd1 _10453_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13279__D line[97] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13171_ _13171_/A _13194_/Y vssd1 vssd1 vccd1 vccd1 _13731_/Z sky130_fd_sc_hd__ebufn_2
X_10383_ _10383_/A _10394_/Y vssd1 vssd1 vccd1 vccd1 _13743_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.M\[2\].MUX\[7\]_A3 _13887_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12122_ _12140_/CLK line[95] vssd1 vssd1 vccd1 vccd1 _12123_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[16\].VALID\[12\].FF_D A[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12053_ _12053_/A _12074_/Y vssd1 vssd1 vccd1 vccd1 _13733_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_2_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11004_ _11020_/CLK line[81] vssd1 vssd1 vccd1 vccd1 _11005_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11527__D line[79] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05525__D line[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12955_ _12955_/A _12984_/Y vssd1 vssd1 vccd1 vccd1 _13795_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13742__D line[53] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11906_ _11930_/CLK line[124] vssd1 vssd1 vccd1 vccd1 _11907_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[26\].VALID\[11\].FF_D A[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08836__D line[114] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12886_ _12910_/CLK line[60] vssd1 vssd1 vccd1 vccd1 _12887_/A sky130_fd_sc_hd__dfxtp_1
X_11837_ _11837_/A _11864_/Y vssd1 vssd1 vccd1 vccd1 _13797_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_14_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05260__D line[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11768_ _11790_/CLK line[61] vssd1 vssd1 vccd1 vccd1 _11769_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_202_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XOVHB\[0\].VALID\[4\].FF OVHB\[0\].V/CLK A[11] vssd1 vssd1 vccd1 vccd1 OVHB\[0\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_186_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10719_ _10719_/A _10744_/Y vssd1 vssd1 vccd1 vccd1 _13799_/Z sky130_fd_sc_hd__ebufn_2
X_13507_ _13507_/CLK _13508_/X vssd1 vssd1 vccd1 vccd1 _13505_/CLK sky130_fd_sc_hd__dlclkp_1
XPHY_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11699_ _11699_/A _11724_/Y vssd1 vssd1 vccd1 vccd1 _13659_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_173_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13438_ _13898_/Y wr vssd1 vssd1 vccd1 vccd1 _13438_/X sky130_fd_sc_hd__and2_1
XOVHB\[28\].VALID\[14\].TOBUF OVHB\[28\].VALID\[14\].FF/Q OVHB\[28\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__12093__D line[67] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13369_ _13898_/Y vssd1 vssd1 vccd1 vccd1 _13369_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07187__D line[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[26\].VALID\[14\].FF OVHB\[26\].V/CLK A[21] vssd1 vssd1 vccd1 vccd1 OVHB\[26\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_07930_ _07940_/CLK line[84] vssd1 vssd1 vccd1 vccd1 _07931_/A sky130_fd_sc_hd__dfxtp_1
X_07861_ _07861_/A _07874_/Y vssd1 vssd1 vccd1 vccd1 _13741_/Z sky130_fd_sc_hd__ebufn_2
X_09600_ _09620_/CLK line[94] vssd1 vssd1 vccd1 vccd1 _09601_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_3_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10341__D line[34] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06812_ _06820_/CLK line[85] vssd1 vssd1 vccd1 vccd1 _06813_/A sky130_fd_sc_hd__dfxtp_1
X_07792_ _07800_/CLK line[21] vssd1 vssd1 vccd1 vccd1 _07793_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_37_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05435__D line[110] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09531_ _09531_/A _09554_/Y vssd1 vssd1 vccd1 vccd1 _13731_/Z sky130_fd_sc_hd__ebufn_2
X_06743_ _06743_/A _06754_/Y vssd1 vssd1 vccd1 vccd1 _13743_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_37_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13652__D line[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[13\].CLKBUF\[2\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09462_ _09480_/CLK line[31] vssd1 vssd1 vccd1 vccd1 _09463_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[27\].VALID\[2\].TOBUF OVHB\[27\].VALID\[2\].FF/Q OVHB\[27\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04930_/B2 sky130_fd_sc_hd__ebufn_2
X_06674_ _06680_/CLK line[22] vssd1 vssd1 vccd1 vccd1 _06675_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07650__D line[84] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08413_ _08413_/A _08434_/Y vssd1 vssd1 vccd1 vccd1 _13733_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12268__D line[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05625_ _05625_/A _05634_/Y vssd1 vssd1 vccd1 vccd1 _13745_/Z sky130_fd_sc_hd__ebufn_2
X_09393_ _09393_/A _09414_/Y vssd1 vssd1 vccd1 vccd1 _13873_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[21\].VALID\[13\].TOBUF OVHB\[21\].VALID\[13\].FF/Q OVHB\[21\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04916_/B2 sky130_fd_sc_hd__ebufn_2
XPHY_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08344_ _08360_/CLK line[17] vssd1 vssd1 vccd1 vccd1 _08345_/A sky130_fd_sc_hd__dfxtp_1
X_05556_ _05560_/CLK line[23] vssd1 vssd1 vccd1 vccd1 _05557_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_32_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[10\].VALID\[7\].FF_D A[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08275_ _08275_/A _08294_/Y vssd1 vssd1 vccd1 vccd1 _13875_/Z sky130_fd_sc_hd__ebufn_2
X_05487_ _05487_/A _05494_/Y vssd1 vssd1 vccd1 vccd1 _13887_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11900__D line[112] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09577__D line[69] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07226_ _07240_/CLK line[18] vssd1 vssd1 vccd1 vccd1 _07227_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[14\].INV _13948_/X vssd1 vssd1 vccd1 vccd1 OVHB\[14\].INV/Y sky130_fd_sc_hd__inv_2
XFILLER_180_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10516__D line[114] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07157_ _07157_/A _07174_/Y vssd1 vssd1 vccd1 vccd1 _13877_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_106_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06108_ _06120_/CLK line[19] vssd1 vssd1 vccd1 vccd1 _06109_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[6\].CLKBUF\[2\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07088_ _07100_/CLK line[83] vssd1 vssd1 vccd1 vccd1 _07089_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_106_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10813__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13827__D line[106] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[29\].INV _13969_/X vssd1 vssd1 vccd1 vccd1 OVHB\[29\].INV/Y sky130_fd_sc_hd__inv_2
XANTENNA__12731__D line[103] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06039_ _06039_/A _06054_/Y vssd1 vssd1 vccd1 vccd1 _13879_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07825__D line[36] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09729_ _13921_/X vssd1 vssd1 vccd1 vccd1 _09729_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12740_ _12770_/CLK line[112] vssd1 vssd1 vccd1 vccd1 _12741_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_28_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07560__D line[48] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12671_ _12671_/A _12704_/Y vssd1 vssd1 vccd1 vccd1 _13791_/Z sky130_fd_sc_hd__ebufn_2
XPHY_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11082__D line[117] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11622_ _11650_/CLK line[122] vssd1 vssd1 vccd1 vccd1 _11623_/A sky130_fd_sc_hd__dfxtp_1
XPHY_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06176__D line[50] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06754__A _13905_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[19\].VALID\[8\].TOBUF OVHB\[19\].VALID\[8\].FF/Q OVHB\[19\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04931_/B2 sky130_fd_sc_hd__ebufn_2
XPHY_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11553_ _11553_/A _11584_/Y vssd1 vssd1 vccd1 vccd1 _13793_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_183_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12906__D line[55] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06473__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09487__D line[42] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08391__D line[39] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10504_ _10530_/CLK line[123] vssd1 vssd1 vccd1 vccd1 _10505_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11484_ _11510_/CLK line[59] vssd1 vssd1 vccd1 vccd1 _11485_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_183_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13223_ _13225_/CLK line[72] vssd1 vssd1 vccd1 vccd1 _13224_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_155_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10435_ _10435_/A _10464_/Y vssd1 vssd1 vccd1 vccd1 _13795_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[23\].V_RESET_B rst_n vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13154_ _13154_/A _13159_/Y vssd1 vssd1 vccd1 vccd1 _13714_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[9\].CLKBUF\[3\] clk vssd1 vssd1 vccd1 vccd1 _13752_/CLK sky130_fd_sc_hd__clkbuf_4
X_10366_ _10390_/CLK line[60] vssd1 vssd1 vccd1 vccd1 _10367_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_151_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12105_ _12105_/CLK line[73] vssd1 vssd1 vccd1 vccd1 _12106_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12641__D line[76] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13085_ _13085_/CLK line[9] vssd1 vssd1 vccd1 vccd1 _13086_/A sky130_fd_sc_hd__dfxtp_1
X_10297_ _10297_/A _10324_/Y vssd1 vssd1 vccd1 vccd1 _13657_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07735__D line[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12036_ _12036_/A _12039_/Y vssd1 vssd1 vccd1 vccd1 _13716_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11257__D line[69] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[30\].VALID\[3\].FF_D A[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09950__D line[126] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06929__A _13909_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06648__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08566__D line[119] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12938_ _12938_/A _12949_/Y vssd1 vssd1 vccd1 vccd1 _13778_/Z sky130_fd_sc_hd__ebufn_2
X_12869_ _12875_/CLK line[38] vssd1 vssd1 vccd1 vccd1 _12870_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_21_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_OVHB\[23\].VALID\[7\].FF_D A[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05410_ _05420_/CLK line[84] vssd1 vssd1 vccd1 vccd1 _05411_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_178_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06390_ _06400_/CLK line[20] vssd1 vssd1 vccd1 vccd1 _06391_/A sky130_fd_sc_hd__dfxtp_1
X_05341_ _05341_/A _05354_/Y vssd1 vssd1 vccd1 vccd1 _13741_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_186_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12816__D line[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11720__D line[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDATA\[29\].CLKBUF\[7\] clk vssd1 vssd1 vccd1 vccd1 _11092_/CLK sky130_fd_sc_hd__clkbuf_4
X_08060_ _08080_/CLK line[30] vssd1 vssd1 vccd1 vccd1 _08061_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06814__D line[86] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[25\].VALID\[1\].FF OVHB\[25\].V/CLK A[8] vssd1 vssd1 vccd1 vccd1 OVHB\[25\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_05272_ _05280_/CLK line[21] vssd1 vssd1 vccd1 vccd1 _05273_/A sky130_fd_sc_hd__dfxtp_1
X_07011_ _07011_/A _07034_/Y vssd1 vssd1 vccd1 vccd1 _13731_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[0\].VALID\[4\].TOBUF OVHB\[0\].VALID\[4\].FF/Q OVHB\[0\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04925_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[1\].CG_CLK clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[25\].VALID\[7\].TOBUF OVHB\[25\].VALID\[7\].FF/Q OVHB\[25\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/A2 sky130_fd_sc_hd__ebufn_2
X_08962_ _08990_/CLK line[58] vssd1 vssd1 vccd1 vccd1 _08963_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_142_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07913_ _07913_/A _07944_/Y vssd1 vssd1 vccd1 vccd1 _13793_/Z sky130_fd_sc_hd__ebufn_2
X_08893_ _08893_/A _08924_/Y vssd1 vssd1 vccd1 vccd1 _13653_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11167__D line[42] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDATA\[8\].CLKBUF\[0\] clk vssd1 vssd1 vccd1 vccd1 _13367_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__10071__D line[39] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07844_ _07870_/CLK line[59] vssd1 vssd1 vccd1 vccd1 _07845_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_68_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05165__D line[100] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07775_ _07775_/A _07804_/Y vssd1 vssd1 vccd1 vccd1 _13655_/Z sky130_fd_sc_hd__ebufn_2
X_04987_ _04987_/A _05004_/Y vssd1 vssd1 vccd1 vccd1 _13667_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13382__D line[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09514_ _09514_/A _09519_/Y vssd1 vssd1 vccd1 vccd1 _13714_/Z sky130_fd_sc_hd__ebufn_2
X_06726_ _06750_/CLK line[60] vssd1 vssd1 vccd1 vccd1 _06727_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08476__D line[92] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07380__D line[89] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09445_ _09445_/CLK line[9] vssd1 vssd1 vccd1 vccd1 _09446_/A sky130_fd_sc_hd__dfxtp_1
X_06657_ _06657_/A _06684_/Y vssd1 vssd1 vccd1 vccd1 _13657_/Z sky130_fd_sc_hd__ebufn_2
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05608_ _05630_/CLK line[61] vssd1 vssd1 vccd1 vccd1 _05609_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_169_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09376_ _09376_/A _09379_/Y vssd1 vssd1 vccd1 vccd1 _13856_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_52_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06588_ _06610_/CLK line[125] vssd1 vssd1 vccd1 vccd1 _06589_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[0\].VOBUF OVHB\[0\].V/Q OVHB\[0\].INV/Y vssd1 vssd1 vccd1 vccd1 _04912_/B1
+ sky130_fd_sc_hd__ebufn_2
XFILLER_33_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_DATA\[11\].CLKBUF\[4\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08327_ _08327_/CLK _08328_/X vssd1 vssd1 vccd1 vccd1 _08325_/CLK sky130_fd_sc_hd__dlclkp_1
X_05539_ _05539_/A _05564_/Y vssd1 vssd1 vccd1 vccd1 _13659_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[22\].VALID\[12\].FF OVHB\[22\].V/CLK A[19] vssd1 vssd1 vccd1 vccd1 OVHB\[22\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_137_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11630__D line[126] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06724__D line[59] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08258_ _13932_/X wr vssd1 vssd1 vccd1 vccd1 _08258_/X sky130_fd_sc_hd__and2_1
XANTENNA__09100__D line[112] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07209_ _13910_/X vssd1 vssd1 vccd1 vccd1 _07209_/Y sky130_fd_sc_hd__inv_2
XANTENNA__10246__D line[119] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08189_ _13932_/X vssd1 vssd1 vccd1 vccd1 _08189_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10220_ _10250_/CLK line[112] vssd1 vssd1 vccd1 vccd1 _10221_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[28\].CLKBUF\[4\] clk vssd1 vssd1 vccd1 vccd1 _10707_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA_OVHB\[4\].VALID\[2\].FF_D A[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13557__D line[111] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10151_ _10151_/A _10184_/Y vssd1 vssd1 vccd1 vccd1 _13791_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07555__D line[41] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08013__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[23\].VALID\[3\].FF OVHB\[23\].V/CLK A[10] vssd1 vssd1 vccd1 vccd1 OVHB\[23\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_10082_ _10110_/CLK line[58] vssd1 vssd1 vccd1 vccd1 _10083_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_121_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13910_ _13916_/C _13916_/B _13916_/A _13916_/D vssd1 vssd1 vccd1 vccd1 _13910_/X
+ sky130_fd_sc_hd__and4bb_4
XANTENNA_DATA\[4\].CLKBUF\[4\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05075__D line[64] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13841_ _13855_/CLK line[98] vssd1 vssd1 vccd1 vccd1 _13842_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11805__D line[78] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XOVHB\[12\].VALID\[14\].FF OVHB\[12\].V/CLK A[21] vssd1 vssd1 vccd1 vccd1 OVHB\[12\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_16_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XOVHB\[31\].VALID\[6\].TOBUF OVHB\[31\].VALID\[6\].FF/Q OVHB\[31\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04923_/A2 sky130_fd_sc_hd__ebufn_2
X_13772_ _13772_/A _13789_/Y vssd1 vssd1 vccd1 vccd1 _13772_/Z sky130_fd_sc_hd__ebufn_2
X_10984_ _10984_/A _10989_/Y vssd1 vssd1 vccd1 vccd1 _13784_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07290__D line[62] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05803__D line[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_DATA\[30\].CLKBUF\[6\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12723_ _12735_/CLK line[99] vssd1 vssd1 vccd1 vccd1 _12724_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_200_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12654_ _12654_/A _12669_/Y vssd1 vssd1 vccd1 vccd1 _13774_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_90_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11605_ _11615_/CLK line[100] vssd1 vssd1 vccd1 vccd1 _11606_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_30_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12585_ _12595_/CLK line[36] vssd1 vssd1 vccd1 vccd1 _12586_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_169_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11536_ _11536_/A _11549_/Y vssd1 vssd1 vccd1 vccd1 _13776_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10156__D line[92] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11467_ _11475_/CLK line[37] vssd1 vssd1 vccd1 vccd1 _11468_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_99_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13206_ _13206_/A _13229_/Y vssd1 vssd1 vccd1 vccd1 _13766_/Z sky130_fd_sc_hd__ebufn_2
X_10418_ _10418_/A _10429_/Y vssd1 vssd1 vccd1 vccd1 _13778_/Z sky130_fd_sc_hd__ebufn_2
X_11398_ _11398_/A _11409_/Y vssd1 vssd1 vccd1 vccd1 _13638_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12371__D line[66] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13137_ _13155_/CLK line[47] vssd1 vssd1 vccd1 vccd1 _13138_/A sky130_fd_sc_hd__dfxtp_1
X_10349_ _10355_/CLK line[38] vssd1 vssd1 vccd1 vccd1 _10350_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07465__D line[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13068_ _13068_/A _13089_/Y vssd1 vssd1 vccd1 vccd1 _13628_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_85_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XDATA\[27\].CLKBUF\[1\] clk vssd1 vssd1 vccd1 vccd1 _10322_/CLK sky130_fd_sc_hd__clkbuf_4
XMUX.M\[3\].MUX\[2\] _13653_/Z _13723_/Z _13793_/Z _13863_/Z MUX.SEL0BUF\[3\]/X MUX.SEL1BUF\[3\]/X
+ vssd1 vssd1 vccd1 vccd1 Do[26] sky130_fd_sc_hd__mux4_1
XFILLER_78_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12019_ _12035_/CLK line[33] vssd1 vssd1 vccd1 vccd1 _12020_/A sky130_fd_sc_hd__dfxtp_1
X_05890_ _05910_/CLK line[62] vssd1 vssd1 vccd1 vccd1 _05891_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09680__D line[116] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05563__A _13901_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDATA\[17\].CLKBUF\[7\] clk vssd1 vssd1 vccd1 vccd1 _07452_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_81_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07560_ _07590_/CLK line[48] vssd1 vssd1 vccd1 vccd1 _07561_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[21\].VALID\[5\].FF OVHB\[21\].V/CLK A[12] vssd1 vssd1 vccd1 vccd1 OVHB\[21\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_207_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05713__D line[109] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06511_ _06511_/A _06544_/Y vssd1 vssd1 vccd1 vccd1 _13791_/Z sky130_fd_sc_hd__ebufn_2
X_07491_ _07491_/A _07524_/Y vssd1 vssd1 vccd1 vccd1 _13651_/Z sky130_fd_sc_hd__ebufn_2
X_09230_ _09230_/A _09239_/Y vssd1 vssd1 vccd1 vccd1 _13710_/Z sky130_fd_sc_hd__ebufn_2
X_06442_ _06470_/CLK line[58] vssd1 vssd1 vccd1 vccd1 _06443_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09161_ _09165_/CLK line[7] vssd1 vssd1 vccd1 vccd1 _09162_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12546__D line[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06373_ _06373_/A _06404_/Y vssd1 vssd1 vccd1 vccd1 _13653_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_147_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[26\].CG clk OVHB\[26\].CGAND/X vssd1 vssd1 vccd1 vccd1 OVHB\[26\].V/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_9_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08112_ _08112_/A _08119_/Y vssd1 vssd1 vccd1 vccd1 _13712_/Z sky130_fd_sc_hd__ebufn_2
X_05324_ _05350_/CLK line[59] vssd1 vssd1 vccd1 vccd1 _05325_/A sky130_fd_sc_hd__dfxtp_1
X_09092_ _09092_/A _09099_/Y vssd1 vssd1 vccd1 vccd1 _13852_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[18\].VALID\[12\].TOBUF OVHB\[18\].VALID\[12\].FF/Q OVHB\[18\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04929_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_119_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12843__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08043_ _08045_/CLK line[8] vssd1 vssd1 vccd1 vccd1 _08044_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_135_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05255_ _05255_/A _05284_/Y vssd1 vssd1 vccd1 vccd1 _13655_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09855__D line[68] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05738__A _13901_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05186_ _05210_/CLK line[124] vssd1 vssd1 vccd1 vccd1 _05187_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_115_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09994_ _09994_/A _10009_/Y vssd1 vssd1 vccd1 vccd1 _13634_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_143_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08945_ _08955_/CLK line[36] vssd1 vssd1 vccd1 vccd1 _08946_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_103_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08876_ _08876_/A _08889_/Y vssd1 vssd1 vccd1 vccd1 _13636_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09590__D line[80] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07827_ _07835_/CLK line[37] vssd1 vssd1 vccd1 vccd1 _07828_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_45_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_DATA\[29\].CLKBUF\[7\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07758_ _07758_/A _07769_/Y vssd1 vssd1 vccd1 vccd1 _13638_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08784__A _13914_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XOVHB\[11\].VALID\[11\].TOBUF OVHB\[11\].VALID\[11\].FF/Q OVHB\[11\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04915_/B2 sky130_fd_sc_hd__ebufn_2
X_06709_ _06715_/CLK line[38] vssd1 vssd1 vccd1 vccd1 _06710_/A sky130_fd_sc_hd__dfxtp_1
X_07689_ _07695_/CLK line[102] vssd1 vssd1 vccd1 vccd1 _07690_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_52_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XDATA\[16\].CLKBUF\[4\] clk vssd1 vssd1 vccd1 vccd1 _07067_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_12_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09428_ _09428_/A _09449_/Y vssd1 vssd1 vccd1 vccd1 _13628_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_197_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09359_ _09375_/CLK line[97] vssd1 vssd1 vccd1 vccd1 _09360_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_12_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XMUX.M\[2\].MUX\[4\] _13671_/Z _13741_/Z _13811_/Z _13881_/Z MUX.SEL0BUF\[2\]/X MUX.SEL1BUF\[2\]/X
+ vssd1 vssd1 vccd1 vccd1 Do[20] sky130_fd_sc_hd__mux4_1
XOVHB\[7\].CGAND _13938_/X wr vssd1 vssd1 vccd1 vccd1 OVHB\[7\].CGAND/X sky130_fd_sc_hd__and2_4
XANTENNA__11360__D line[116] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12370_ _12370_/A _12389_/Y vssd1 vssd1 vccd1 vccd1 _13770_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06454__D line[49] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11321_ _11335_/CLK line[98] vssd1 vssd1 vccd1 vccd1 _11322_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_176_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09765__D line[32] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11252_ _11252_/A _11269_/Y vssd1 vssd1 vccd1 vccd1 _13772_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_125_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13287__D line[101] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10203_ _10215_/CLK line[99] vssd1 vssd1 vccd1 vccd1 _10204_/A sky130_fd_sc_hd__dfxtp_1
X_11183_ _11195_/CLK line[35] vssd1 vssd1 vccd1 vccd1 _11184_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[7\].VALID\[4\].TOBUF OVHB\[7\].VALID\[4\].FF/Q OVHB\[7\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04925_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__08959__A _13915_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10134_ _10134_/A _10149_/Y vssd1 vssd1 vccd1 vccd1 _13774_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_67_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08678__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10065_ _10075_/CLK line[36] vssd1 vssd1 vccd1 vccd1 _10066_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_125_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11535__D line[68] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06629__D line[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13824_ _13899_/X vssd1 vssd1 vccd1 vccd1 _13824_/Y sky130_fd_sc_hd__inv_2
XANTENNA__09005__D line[78] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13755_ _13785_/CLK line[64] vssd1 vssd1 vccd1 vccd1 _13756_/A sky130_fd_sc_hd__dfxtp_1
X_10967_ _10985_/CLK line[79] vssd1 vssd1 vccd1 vccd1 _10968_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_16_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13750__D line[57] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_DATA\[2\].CLKBUF\[6\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12706_ _12706_/A _12739_/Y vssd1 vssd1 vccd1 vccd1 _13826_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08844__D line[118] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13686_ _13686_/A _13719_/Y vssd1 vssd1 vccd1 vccd1 _13686_/Z sky130_fd_sc_hd__ebufn_2
X_10898_ _10898_/A _10919_/Y vssd1 vssd1 vccd1 vccd1 _13698_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[18\].VALID\[8\].FF OVHB\[18\].V/CLK A[15] vssd1 vssd1 vccd1 vccd1 OVHB\[18\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07103__A _13909_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12637_ _12665_/CLK line[74] vssd1 vssd1 vccd1 vccd1 _12638_/A sky130_fd_sc_hd__dfxtp_1
XPHY_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11270__D line[80] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XDATA\[15\].CLKBUF\[1\] clk vssd1 vssd1 vccd1 vccd1 _06682_/CLK sky130_fd_sc_hd__clkbuf_4
X_12568_ _12568_/A _12599_/Y vssd1 vssd1 vccd1 vccd1 _13688_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11519_ _11545_/CLK line[75] vssd1 vssd1 vccd1 vccd1 _11520_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_157_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12499_ _12525_/CLK line[11] vssd1 vssd1 vccd1 vccd1 _12500_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10464__A _13923_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05040_ _05070_/CLK line[48] vssd1 vssd1 vccd1 vccd1 _05041_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_172_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13197__D line[74] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10183__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07195__D line[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06991_ _06995_/CLK line[39] vssd1 vssd1 vccd1 vccd1 _06992_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_86_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMUX.M\[1\].MUX\[6\] _13626_/Z _13696_/Z _13766_/Z _13836_/Z MUX.SEL0BUF\[1\]/X MUX.SEL1BUF\[1\]/X
+ vssd1 vssd1 vccd1 vccd1 Do[14] sky130_fd_sc_hd__mux4_1
XOVHB\[31\].VALID\[11\].TOBUF OVHB\[31\].VALID\[11\].FF/Q OVHB\[31\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04915_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_39_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08730_ _08730_/A _08749_/Y vssd1 vssd1 vccd1 vccd1 _13770_/Z sky130_fd_sc_hd__ebufn_2
X_05942_ _05942_/A _05949_/Y vssd1 vssd1 vccd1 vccd1 _13782_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_38_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08661_ _08675_/CLK line[34] vssd1 vssd1 vccd1 vccd1 _08662_/A sky130_fd_sc_hd__dfxtp_1
X_05873_ _05875_/CLK line[40] vssd1 vssd1 vccd1 vccd1 _05874_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11445__D line[32] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07612_ _07612_/A _07629_/Y vssd1 vssd1 vccd1 vccd1 _13772_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_38_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08592_ _08592_/A _08609_/Y vssd1 vssd1 vccd1 vccd1 _13632_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05443__D line[99] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07543_ _07555_/CLK line[35] vssd1 vssd1 vccd1 vccd1 _07544_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13660__D line[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10639__A _13924_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07474_ _07474_/A _07489_/Y vssd1 vssd1 vccd1 vccd1 _13634_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08754__D line[91] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10358__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09213_ _09235_/CLK line[45] vssd1 vssd1 vccd1 vccd1 _09214_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12276__D line[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06425_ _06435_/CLK line[36] vssd1 vssd1 vccd1 vccd1 _06426_/A sky130_fd_sc_hd__dfxtp_1
X_09144_ _09144_/A _09169_/Y vssd1 vssd1 vccd1 vccd1 _13624_/Z sky130_fd_sc_hd__ebufn_2
X_06356_ _06356_/A _06369_/Y vssd1 vssd1 vccd1 vccd1 _13636_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_30_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05307_ _05315_/CLK line[37] vssd1 vssd1 vccd1 vccd1 _05308_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[0\].VALID\[5\].FF_D A[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09075_ _09095_/CLK line[110] vssd1 vssd1 vccd1 vccd1 _09076_/A sky130_fd_sc_hd__dfxtp_1
X_06287_ _06295_/CLK line[101] vssd1 vssd1 vccd1 vccd1 _06288_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09585__D line[73] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08026_ _08026_/A _08049_/Y vssd1 vssd1 vccd1 vccd1 _13626_/Z sky130_fd_sc_hd__ebufn_2
X_05238_ _05238_/A _05249_/Y vssd1 vssd1 vccd1 vccd1 _13638_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_163_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10524__D line[118] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05169_ _05175_/CLK line[102] vssd1 vssd1 vccd1 vccd1 _05170_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05618__D line[51] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09977_ _10005_/CLK line[10] vssd1 vssd1 vccd1 vccd1 _09978_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_89_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13835__D line[110] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08928_ _08928_/A _08959_/Y vssd1 vssd1 vccd1 vccd1 _13688_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08929__D line[43] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06299__A _13903_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07833__D line[40] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08859_ _08885_/CLK line[11] vssd1 vssd1 vccd1 vccd1 _08860_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_57_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11933__A _13927_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11870_ _11870_/A _11899_/Y vssd1 vssd1 vccd1 vccd1 _13830_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_169_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10821_ _10845_/CLK line[12] vssd1 vssd1 vccd1 vccd1 _10822_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_60_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10752_ _10752_/A _10779_/Y vssd1 vssd1 vccd1 vccd1 _13832_/Z sky130_fd_sc_hd__ebufn_2
X_13540_ _13540_/CLK line[89] vssd1 vssd1 vccd1 vccd1 _13541_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_198_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[5\].VALID\[9\].TOBUF OVHB\[5\].VALID\[9\].FF/Q OVHB\[5\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04914_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[3\].VALID\[11\].FF_D A[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12186__D line[124] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13471_ _13471_/A _13474_/Y vssd1 vssd1 vccd1 vccd1 _13751_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11090__D line[121] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10683_ _10705_/CLK line[77] vssd1 vssd1 vccd1 vccd1 _10684_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06184__D line[54] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12422_ _12422_/CLK _12423_/X vssd1 vssd1 vccd1 vccd1 _12420_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_166_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_DATA\[23\].CLKBUF\[0\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12353_ _13935_/X wr vssd1 vssd1 vccd1 vccd1 _12353_/X sky130_fd_sc_hd__and2_1
XFILLER_138_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09495__D line[46] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11304_ _13933_/X vssd1 vssd1 vccd1 vccd1 _11304_/Y sky130_fd_sc_hd__inv_2
X_12284_ _13935_/X vssd1 vssd1 vccd1 vccd1 _12284_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11235_ _11265_/CLK line[64] vssd1 vssd1 vccd1 vccd1 _11236_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_107_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10434__D line[91] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07593__A _13911_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11166_ _11166_/A _11199_/Y vssd1 vssd1 vccd1 vccd1 _13686_/Z sky130_fd_sc_hd__ebufn_2
X_10117_ _10145_/CLK line[74] vssd1 vssd1 vccd1 vccd1 _10118_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[15\].VALID\[2\].FF_D A[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12004__A _13934_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11097_ _11125_/CLK line[10] vssd1 vssd1 vccd1 vccd1 _11098_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07743__D line[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[3\].VALID\[14\].FF OVHB\[3\].V/CLK A[21] vssd1 vssd1 vccd1 vccd1 OVHB\[3\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_10048_ _10048_/A _10079_/Y vssd1 vssd1 vccd1 vccd1 _13688_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11265__D line[73] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06359__D line[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MUX.M\[0\].MUX\[6\]_A2 _13780_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13807_ _13807_/A _13824_/Y vssd1 vssd1 vccd1 vccd1 _13807_/Z sky130_fd_sc_hd__ebufn_2
X_11999_ _11999_/A _12004_/Y vssd1 vssd1 vccd1 vccd1 _13679_/Z sky130_fd_sc_hd__ebufn_2
X_13738_ _13750_/CLK line[51] vssd1 vssd1 vccd1 vccd1 _13739_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_204_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10609__D line[43] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13669_ _13669_/A _13684_/Y vssd1 vssd1 vccd1 vccd1 _13669_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06210_ _06210_/A _06229_/Y vssd1 vssd1 vccd1 vccd1 _13770_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06094__D line[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07768__A _13912_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07190_ _07190_/A _07209_/Y vssd1 vssd1 vccd1 vccd1 _13630_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_157_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06141_ _06155_/CLK line[34] vssd1 vssd1 vccd1 vccd1 _06142_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[4\].V OVHB\[4\].V/CLK TIE/HI rst_n vssd1 vssd1 vccd1 vccd1 OVHB\[4\].V/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12824__D line[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07918__D line[93] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06072_ _06072_/A _06089_/Y vssd1 vssd1 vccd1 vccd1 _13632_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[12\].VALID\[4\].TOBUF OVHB\[12\].VALID\[4\].FF/Q OVHB\[12\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04925_/B2 sky130_fd_sc_hd__ebufn_2
X_09900_ _09900_/CLK line[89] vssd1 vssd1 vccd1 vccd1 _09901_/A sky130_fd_sc_hd__dfxtp_1
X_05023_ _05035_/CLK line[35] vssd1 vssd1 vccd1 vccd1 _05024_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[6\].VALID\[9\].FF_D A[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDEC.DEC0.AND1 A[6] A[5] vssd1 vssd1 vccd1 vccd1 _13905_/D sky130_fd_sc_hd__and2b_2
X_09831_ _09831_/A _09834_/Y vssd1 vssd1 vccd1 vccd1 _13751_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__04920__A A_h[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09762_ _09762_/CLK _09763_/X vssd1 vssd1 vccd1 vccd1 _09760_/CLK sky130_fd_sc_hd__dlclkp_1
X_06974_ _06974_/A _06999_/Y vssd1 vssd1 vccd1 vccd1 _13694_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_39_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08713_ _13914_/X wr vssd1 vssd1 vccd1 vccd1 _08713_/X sky130_fd_sc_hd__and2_1
X_05925_ _05945_/CLK line[78] vssd1 vssd1 vccd1 vccd1 _05926_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_100_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09693_ _13920_/Y wr vssd1 vssd1 vccd1 vccd1 _09693_/X sky130_fd_sc_hd__and2_1
XANTENNA__11175__D line[46] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08644_ _13914_/X vssd1 vssd1 vccd1 vccd1 _08644_/Y sky130_fd_sc_hd__inv_2
XANTENNA__06269__D line[107] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05856_ _05856_/A _05879_/Y vssd1 vssd1 vccd1 vccd1 _13696_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05173__D line[104] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XOVHB\[27\].VALID\[12\].FF OVHB\[27\].V/CLK A[19] vssd1 vssd1 vccd1 vccd1 OVHB\[27\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08575_ _08605_/CLK line[0] vssd1 vssd1 vccd1 vccd1 _08576_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05787_ _05805_/CLK line[15] vssd1 vssd1 vccd1 vccd1 _05788_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13390__D line[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07526_ _07526_/A _07559_/Y vssd1 vssd1 vccd1 vccd1 _13686_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08484__D line[81] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07457_ _07485_/CLK line[10] vssd1 vssd1 vccd1 vccd1 _07458_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06408_ _06408_/A _06439_/Y vssd1 vssd1 vccd1 vccd1 _13688_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_155_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07388_ _07388_/A _07419_/Y vssd1 vssd1 vccd1 vccd1 _13828_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_210_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09127_ _09127_/A _09134_/Y vssd1 vssd1 vccd1 vccd1 _13887_/Z sky130_fd_sc_hd__ebufn_2
X_06339_ _06365_/CLK line[11] vssd1 vssd1 vccd1 vccd1 _06340_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06732__D line[63] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09058_ _09060_/CLK line[88] vssd1 vssd1 vccd1 vccd1 _09059_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_2_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08009_ _08009_/A _08014_/Y vssd1 vssd1 vccd1 vccd1 _13889_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[9\].VALID\[3\].FF OVHB\[9\].V/CLK A[10] vssd1 vssd1 vccd1 vccd1 OVHB\[9\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__05348__D line[56] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11020_ _11020_/CLK line[89] vssd1 vssd1 vccd1 vccd1 _11021_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_150_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[28\].VALID\[2\].FF_D A[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[17\].VALID\[14\].FF OVHB\[17\].V/CLK A[21] vssd1 vssd1 vccd1 vccd1 OVHB\[17\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13565__D line[100] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08659__D line[33] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12971_ _12971_/A _12984_/Y vssd1 vssd1 vccd1 vccd1 _13811_/Z sky130_fd_sc_hd__ebufn_2
X_11922_ _11930_/CLK line[117] vssd1 vssd1 vccd1 vccd1 _11923_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05083__D line[77] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09133__A _13915_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11853_ _11853_/A _11864_/Y vssd1 vssd1 vccd1 vccd1 _13813_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_73_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11813__D line[67] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10804_ _10810_/CLK line[118] vssd1 vssd1 vccd1 vccd1 _10805_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06907__D line[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11784_ _11790_/CLK line[54] vssd1 vssd1 vccd1 vccd1 _11785_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_82_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13523_ _13523_/A _13544_/Y vssd1 vssd1 vccd1 vccd1 _13803_/Z sky130_fd_sc_hd__ebufn_2
X_10735_ _10735_/A _10744_/Y vssd1 vssd1 vccd1 vccd1 _13815_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12494__A _13935_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[8\].VALID\[14\].TOBUF OVHB\[8\].VALID\[14\].FF/Q OVHB\[8\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/B2 sky130_fd_sc_hd__ebufn_2
X_13454_ _13470_/CLK line[49] vssd1 vssd1 vccd1 vccd1 _13455_/A sky130_fd_sc_hd__dfxtp_1
X_10666_ _10670_/CLK line[55] vssd1 vssd1 vccd1 vccd1 _10667_/A sky130_fd_sc_hd__dfxtp_1
X_12405_ _12405_/A _12424_/Y vssd1 vssd1 vccd1 vccd1 _13805_/Z sky130_fd_sc_hd__ebufn_2
X_13385_ _13385_/A _13404_/Y vssd1 vssd1 vccd1 vccd1 _13665_/Z sky130_fd_sc_hd__ebufn_2
X_10597_ _10597_/A _10604_/Y vssd1 vssd1 vccd1 vccd1 _13677_/Z sky130_fd_sc_hd__ebufn_2
X_12336_ _12350_/CLK line[50] vssd1 vssd1 vccd1 vccd1 _12337_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10164__D line[81] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12267_ _12267_/A _12284_/Y vssd1 vssd1 vccd1 vccd1 _13667_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05258__D line[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11218_ _11230_/CLK line[51] vssd1 vssd1 vccd1 vccd1 _11219_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09308__A _13916_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12198_ _12210_/CLK line[115] vssd1 vssd1 vccd1 vccd1 _12199_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[21\].CLKBUF\[2\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13475__D line[64] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11149_ _11149_/A _11164_/Y vssd1 vssd1 vccd1 vccd1 _13669_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07473__D line[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12669__A _13936_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[7\].VALID\[5\].FF OVHB\[7\].V/CLK A[12] vssd1 vssd1 vccd1 vccd1 OVHB\[7\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_05710_ _05710_/A _05739_/Y vssd1 vssd1 vccd1 vccd1 _13830_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[28\].VALID\[10\].TOBUF OVHB\[28\].VALID\[10\].FF/Q OVHB\[28\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04932_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_36_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06690_ _06690_/A _06719_/Y vssd1 vssd1 vccd1 vccd1 _13690_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[1\].VALID\[13\].TOBUF OVHB\[1\].VALID\[13\].FF/Q OVHB\[1\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04916_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__12388__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05641_ _05665_/CLK line[76] vssd1 vssd1 vccd1 vccd1 _05642_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_23_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08360_ _08360_/CLK line[25] vssd1 vssd1 vccd1 vccd1 _08361_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[10\].VALID\[9\].TOBUF OVHB\[10\].VALID\[9\].FF/Q OVHB\[10\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04914_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_23_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05572_ _05572_/A _05599_/Y vssd1 vssd1 vccd1 vccd1 _13692_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05721__D line[98] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07311_ _07311_/A _07314_/Y vssd1 vssd1 vccd1 vccd1 _13751_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_20_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10339__D line[33] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08291_ _08291_/A _08294_/Y vssd1 vssd1 vccd1 vccd1 _13891_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[6\].CLKBUF\[5\] clk vssd1 vssd1 vccd1 vccd1 _12982_/CLK sky130_fd_sc_hd__clkbuf_4
X_07242_ _07242_/CLK _07243_/X vssd1 vssd1 vccd1 vccd1 _07240_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_177_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07173_ _13909_/Y wr vssd1 vssd1 vccd1 vccd1 _07173_/X sky130_fd_sc_hd__and2_1
XANTENNA__12554__D line[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07648__D line[83] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06124_ _13903_/X vssd1 vssd1 vccd1 vccd1 _06124_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06055_ _06085_/CLK line[0] vssd1 vssd1 vccd1 vccd1 _06056_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_105_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09863__D line[72] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05006_ _05006_/A _05039_/Y vssd1 vssd1 vccd1 vccd1 _13686_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13963__A A_h[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10802__D line[117] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09814_ _09830_/CLK line[49] vssd1 vssd1 vccd1 vccd1 _09815_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_98_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09745_ _09745_/A _09764_/Y vssd1 vssd1 vccd1 vccd1 _13665_/Z sky130_fd_sc_hd__ebufn_2
X_06957_ _06957_/A _06964_/Y vssd1 vssd1 vccd1 vccd1 _13677_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_39_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05908_ _05910_/CLK line[56] vssd1 vssd1 vccd1 vccd1 _05909_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_100_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06888_ _06890_/CLK line[120] vssd1 vssd1 vccd1 vccd1 _06889_/A sky130_fd_sc_hd__dfxtp_1
X_09676_ _09690_/CLK line[114] vssd1 vssd1 vccd1 vccd1 _09677_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_55_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12729__D line[102] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08627_ _08627_/A _08644_/Y vssd1 vssd1 vccd1 vccd1 _13667_/Z sky130_fd_sc_hd__ebufn_2
X_05839_ _05839_/A _05844_/Y vssd1 vssd1 vccd1 vccd1 _13679_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_55_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08558_ _08570_/CLK line[115] vssd1 vssd1 vccd1 vccd1 _08559_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[5\].VALID\[7\].FF OVHB\[5\].V/CLK A[14] vssd1 vssd1 vccd1 vccd1 OVHB\[5\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_07509_ _07509_/A _07524_/Y vssd1 vssd1 vccd1 vccd1 _13669_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08489_ _08489_/A _08504_/Y vssd1 vssd1 vccd1 vccd1 _13809_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10520_ _10530_/CLK line[116] vssd1 vssd1 vccd1 vccd1 _10521_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12464__D line[123] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10451_ _10451_/A _10464_/Y vssd1 vssd1 vccd1 vccd1 _13811_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_164_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XDATA\[5\].CLKBUF\[2\] clk vssd1 vssd1 vccd1 vccd1 _12597_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__06462__D line[53] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13170_ _13190_/CLK line[62] vssd1 vssd1 vccd1 vccd1 _13171_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_201_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10382_ _10390_/CLK line[53] vssd1 vssd1 vccd1 vccd1 _10383_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[22\].V_RESET_B rst_n vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12121_ _12121_/A _12144_/Y vssd1 vssd1 vccd1 vccd1 _13801_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_151_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09773__D line[45] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12052_ _12070_/CLK line[63] vssd1 vssd1 vccd1 vccd1 _12053_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_111_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_OVHB\[11\].VALID\[5\].FF_D A[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09051__TE_B _09064_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13295__D line[105] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11003_ _11003_/A _11024_/Y vssd1 vssd1 vccd1 vccd1 _13803_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[19\].VALID\[4\].TOBUF OVHB\[19\].VALID\[4\].FF/Q OVHB\[19\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04925_/B2 sky130_fd_sc_hd__ebufn_2
XOVHB\[23\].VALID\[10\].FF OVHB\[23\].V/CLK A[17] vssd1 vssd1 vccd1 vccd1 OVHB\[23\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10712__D line[90] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08389__D line[38] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12954_ _12980_/CLK line[91] vssd1 vssd1 vccd1 vccd1 _12955_/A sky130_fd_sc_hd__dfxtp_1
X_11905_ _11905_/A _11934_/Y vssd1 vssd1 vccd1 vccd1 _13865_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12639__D line[75] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11543__D line[72] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12885_ _12885_/A _12914_/Y vssd1 vssd1 vccd1 vccd1 _13725_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_45_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06637__D line[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09798__A _13921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11836_ _11860_/CLK line[92] vssd1 vssd1 vccd1 vccd1 _11837_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09013__D line[67] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[3\].CGAND_A _13934_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XDATA\[25\].CLKBUF\[6\] clk vssd1 vssd1 vccd1 vccd1 _09937_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_159_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11767_ _11767_/A _11794_/Y vssd1 vssd1 vccd1 vccd1 _13727_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09948__D line[125] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13506_ _13506_/A _13509_/Y vssd1 vssd1 vccd1 vccd1 _13786_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10718_ _10740_/CLK line[93] vssd1 vssd1 vccd1 vccd1 _10719_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11698_ _11720_/CLK line[29] vssd1 vssd1 vccd1 vccd1 _11699_/A sky130_fd_sc_hd__dfxtp_1
X_13437_ _13437_/CLK _13438_/X vssd1 vssd1 vccd1 vccd1 _13435_/CLK sky130_fd_sc_hd__dlclkp_1
X_10649_ _10649_/A _10674_/Y vssd1 vssd1 vccd1 vccd1 _13729_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[13\].VALID\[12\].FF OVHB\[13\].V/CLK A[19] vssd1 vssd1 vccd1 vccd1 OVHB\[13\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06372__D line[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13368_ _13898_/Y wr vssd1 vssd1 vccd1 vccd1 _13368_/X sky130_fd_sc_hd__and2_1
XOVHB\[3\].VALID\[9\].FF OVHB\[3\].V/CLK A[16] vssd1 vssd1 vccd1 vccd1 OVHB\[3\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[10\].VALID\[13\].FF_D A[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12319_ _13935_/X vssd1 vssd1 vccd1 vccd1 _12319_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13299_ _13938_/X vssd1 vssd1 vccd1 vccd1 _13299_/Y sky130_fd_sc_hd__inv_2
XFILLER_114_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11718__D line[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08299__D line[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07860_ _07870_/CLK line[52] vssd1 vssd1 vccd1 vccd1 _07861_/A sky130_fd_sc_hd__dfxtp_1
X_06811_ _06811_/A _06824_/Y vssd1 vssd1 vccd1 vccd1 _13811_/Z sky130_fd_sc_hd__ebufn_2
X_07791_ _07791_/A _07804_/Y vssd1 vssd1 vccd1 vccd1 _13671_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_68_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09530_ _09550_/CLK line[62] vssd1 vssd1 vccd1 vccd1 _09531_/A sky130_fd_sc_hd__dfxtp_1
X_06742_ _06750_/CLK line[53] vssd1 vssd1 vccd1 vccd1 _06743_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[0\].VALID\[0\].TOBUF OVHB\[0\].VALID\[0\].FF/Q OVHB\[0\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04924_/B2 sky130_fd_sc_hd__ebufn_2
X_09461_ _09461_/A _09484_/Y vssd1 vssd1 vccd1 vccd1 _13661_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[20\].VALID\[12\].FF_D A[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06673_ _06673_/A _06684_/Y vssd1 vssd1 vccd1 vccd1 _13673_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11453__D line[45] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08412_ _08430_/CLK line[63] vssd1 vssd1 vccd1 vccd1 _08413_/A sky130_fd_sc_hd__dfxtp_1
X_05624_ _05630_/CLK line[54] vssd1 vssd1 vccd1 vccd1 _05625_/A sky130_fd_sc_hd__dfxtp_1
X_09392_ _09410_/CLK line[127] vssd1 vssd1 vccd1 vccd1 _09393_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[25\].VALID\[3\].TOBUF OVHB\[25\].VALID\[3\].FF/Q OVHB\[25\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04919_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__06547__D line[106] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05451__D line[103] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08343_ _08343_/A _08364_/Y vssd1 vssd1 vccd1 vccd1 _13663_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10069__D line[38] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05555_ _05555_/A _05564_/Y vssd1 vssd1 vccd1 vccd1 _13675_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[31\].VALID\[1\].FF_D A[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08762__D line[95] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08274_ _08290_/CLK line[113] vssd1 vssd1 vccd1 vccd1 _08275_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_165_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05486_ _05490_/CLK line[119] vssd1 vssd1 vccd1 vccd1 _05487_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_192_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07225_ _07225_/A _07244_/Y vssd1 vssd1 vccd1 vccd1 _13665_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XDATA\[24\].CLKBUF\[3\] clk vssd1 vssd1 vccd1 vccd1 _09552_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_146_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XOVHB\[31\].VALID\[3\].FF OVHB\[31\].V/CLK A[10] vssd1 vssd1 vccd1 vccd1 OVHB\[31\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_192_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07378__D line[88] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07156_ _07170_/CLK line[114] vssd1 vssd1 vccd1 vccd1 _07157_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[30\].VALID\[11\].FF_D A[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[24\].VALID\[5\].FF_D A[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06107_ _06107_/A _06124_/Y vssd1 vssd1 vccd1 vccd1 _13667_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11478__A _13926_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07087_ _07087_/A _07104_/Y vssd1 vssd1 vccd1 vccd1 _13807_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_105_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06038_ _06050_/CLK line[115] vssd1 vssd1 vccd1 vccd1 _06039_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11628__D line[125] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05626__D line[55] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[17\].VALID\[9\].FF_D A[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08002__D line[117] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13843__D line[99] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07989_ _07989_/A _08014_/Y vssd1 vssd1 vccd1 vccd1 _13869_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09728_ _13921_/X wr vssd1 vssd1 vccd1 vccd1 _09728_/X sky130_fd_sc_hd__and2_1
XANTENNA__08937__D line[47] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09659_ _13920_/Y vssd1 vssd1 vccd1 vccd1 _09659_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12670_ _12700_/CLK line[80] vssd1 vssd1 vccd1 vccd1 _12671_/A sky130_fd_sc_hd__dfxtp_1
XPHY_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05361__D line[76] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11621_ _11621_/A _11654_/Y vssd1 vssd1 vccd1 vccd1 _13861_/Z sky130_fd_sc_hd__ebufn_2
XPHY_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[24\].V_D TIE/HI vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[17\].VALID\[9\].TOBUF OVHB\[17\].VALID\[9\].FF/Q OVHB\[17\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04914_/B2 sky130_fd_sc_hd__ebufn_2
X_11552_ _11580_/CLK line[90] vssd1 vssd1 vccd1 vccd1 _11553_/A sky130_fd_sc_hd__dfxtp_1
XPHY_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12194__D line[113] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10503_ _10503_/A _10534_/Y vssd1 vssd1 vccd1 vccd1 _13863_/Z sky130_fd_sc_hd__ebufn_2
X_11483_ _11483_/A _11514_/Y vssd1 vssd1 vccd1 vccd1 _13723_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07288__D line[61] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13222_ _13222_/A _13229_/Y vssd1 vssd1 vccd1 vccd1 _13782_/Z sky130_fd_sc_hd__ebufn_2
X_10434_ _10460_/CLK line[91] vssd1 vssd1 vccd1 vccd1 _10435_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[31\].VALID\[2\].TOBUF OVHB\[31\].VALID\[2\].FF/Q OVHB\[31\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04930_/B2 sky130_fd_sc_hd__ebufn_2
X_10365_ _10365_/A _10394_/Y vssd1 vssd1 vccd1 vccd1 _13725_/Z sky130_fd_sc_hd__ebufn_2
X_13153_ _13155_/CLK line[40] vssd1 vssd1 vccd1 vccd1 _13154_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_128_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XOVHB\[8\].VALID\[14\].FF OVHB\[8\].V/CLK A[21] vssd1 vssd1 vccd1 vccd1 OVHB\[8\].VALID\[14\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_88_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XOVHB\[12\].VALID\[1\].FF OVHB\[12\].V/CLK A[8] vssd1 vssd1 vccd1 vccd1 OVHB\[12\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XDATA\[23\].CLKBUF\[0\] clk vssd1 vssd1 vccd1 vccd1 _09167_/CLK sky130_fd_sc_hd__clkbuf_4
X_12104_ _12104_/A _12109_/Y vssd1 vssd1 vccd1 vccd1 _13784_/Z sky130_fd_sc_hd__ebufn_2
X_13084_ _13084_/A _13089_/Y vssd1 vssd1 vccd1 vccd1 _13644_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_97_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10296_ _10320_/CLK line[28] vssd1 vssd1 vccd1 vccd1 _10297_/A sky130_fd_sc_hd__dfxtp_1
X_12035_ _12035_/CLK line[41] vssd1 vssd1 vccd1 vccd1 _12036_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10442__D line[95] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05536__D line[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDATA\[13\].CLKBUF\[6\] clk vssd1 vssd1 vccd1 vccd1 _06297_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_92_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_DATA\[18\].CLKBUF\[5\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[5\].VALID\[0\].FF_D A[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07751__D line[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12369__D line[65] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12937_ _12945_/CLK line[69] vssd1 vssd1 vccd1 vccd1 _12938_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_73_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12868_ _12868_/A _12879_/Y vssd1 vssd1 vccd1 vccd1 _13708_/Z sky130_fd_sc_hd__ebufn_2
X_11819_ _11825_/CLK line[70] vssd1 vssd1 vccd1 vccd1 _11820_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12799_ _12805_/CLK line[6] vssd1 vssd1 vccd1 vccd1 _12800_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09678__D line[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05340_ _05350_/CLK line[52] vssd1 vssd1 vccd1 vccd1 _05341_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_119_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05271_ _05271_/A _05284_/Y vssd1 vssd1 vccd1 vccd1 _13671_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10617__D line[47] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07010_ _07030_/CLK line[62] vssd1 vssd1 vccd1 vccd1 _07011_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_155_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12832__D line[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07926__D line[82] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[28\].VALID\[6\].FF OVHB\[28\].V/CLK A[13] vssd1 vssd1 vccd1 vccd1 OVHB\[28\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_08961_ _08961_/A _08994_/Y vssd1 vssd1 vccd1 vccd1 _13721_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_88_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XOVHB\[23\].VALID\[8\].TOBUF OVHB\[23\].VALID\[8\].FF/Q OVHB\[23\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04931_/B2 sky130_fd_sc_hd__ebufn_2
X_07912_ _07940_/CLK line[90] vssd1 vssd1 vccd1 vccd1 _07913_/A sky130_fd_sc_hd__dfxtp_1
X_08892_ _08920_/CLK line[26] vssd1 vssd1 vccd1 vccd1 _08893_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_111_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07843_ _07843_/A _07874_/Y vssd1 vssd1 vccd1 vccd1 _13723_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_96_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13018__A _13937_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XOVHB\[10\].VALID\[3\].FF OVHB\[10\].V/CLK A[10] vssd1 vssd1 vccd1 vccd1 OVHB\[10\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_04986_ _05000_/CLK line[18] vssd1 vssd1 vccd1 vccd1 _04987_/A sky130_fd_sc_hd__dfxtp_1
X_07774_ _07800_/CLK line[27] vssd1 vssd1 vccd1 vccd1 _07775_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_209_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XDATA\[12\].CLKBUF\[3\] clk vssd1 vssd1 vccd1 vccd1 _05912_/CLK sky130_fd_sc_hd__clkbuf_4
X_09513_ _09515_/CLK line[40] vssd1 vssd1 vccd1 vccd1 _09514_/A sky130_fd_sc_hd__dfxtp_1
X_06725_ _06725_/A _06754_/Y vssd1 vssd1 vccd1 vccd1 _13725_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_24_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11183__D line[35] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09444_ _09444_/A _09449_/Y vssd1 vssd1 vccd1 vccd1 _13644_/Z sky130_fd_sc_hd__ebufn_2
X_06656_ _06680_/CLK line[28] vssd1 vssd1 vccd1 vccd1 _06657_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06277__D line[111] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05607_ _05607_/A _05634_/Y vssd1 vssd1 vccd1 vccd1 _13727_/Z sky130_fd_sc_hd__ebufn_2
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09375_ _09375_/CLK line[105] vssd1 vssd1 vccd1 vccd1 _09376_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_12_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06587_ _06587_/A _06614_/Y vssd1 vssd1 vccd1 vccd1 _13867_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_149_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05538_ _05560_/CLK line[29] vssd1 vssd1 vccd1 vccd1 _05539_/A sky130_fd_sc_hd__dfxtp_1
X_08326_ _08326_/A _08329_/Y vssd1 vssd1 vccd1 vccd1 _13646_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08492__D line[85] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08257_ _08257_/CLK _08258_/X vssd1 vssd1 vccd1 vccd1 _08255_/CLK sky130_fd_sc_hd__dlclkp_1
X_05469_ _05469_/A _05494_/Y vssd1 vssd1 vccd1 vccd1 _13869_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_137_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07208_ _13910_/X wr vssd1 vssd1 vccd1 vccd1 _07208_/X sky130_fd_sc_hd__and2_1
X_08188_ _13932_/X wr vssd1 vssd1 vccd1 vccd1 _08188_/X sky130_fd_sc_hd__and2_1
XFILLER_118_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07139_ _13909_/Y vssd1 vssd1 vccd1 vccd1 _07139_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12742__D line[122] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06740__D line[52] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10150_ _10180_/CLK line[80] vssd1 vssd1 vccd1 vccd1 _10151_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_79_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_OVHB\[17\].VALID\[13\].FF_D A[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11358__D line[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10081_ _10081_/A _10114_/Y vssd1 vssd1 vccd1 vccd1 _13721_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[3\].CGAND _13934_/X wr vssd1 vssd1 vccd1 vccd1 OVHB\[3\].CGAND/X sky130_fd_sc_hd__and2_4
XANTENNA_OVHB\[9\].V_D TIE/HI vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_199_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13573__D line[104] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08667__D line[37] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13840_ _13840_/A _13859_/Y vssd1 vssd1 vccd1 vccd1 _13840_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[26\].VALID\[8\].FF OVHB\[26\].V/CLK A[15] vssd1 vssd1 vccd1 vccd1 OVHB\[26\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_13771_ _13785_/CLK line[66] vssd1 vssd1 vccd1 vccd1 _13772_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_204_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10983_ _10985_/CLK line[72] vssd1 vssd1 vccd1 vccd1 _10984_/A sky130_fd_sc_hd__dfxtp_1
X_12722_ _12722_/A _12739_/Y vssd1 vssd1 vccd1 vccd1 _13842_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_43_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05091__D line[66] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[7\].VALID\[0\].TOBUF OVHB\[7\].VALID\[0\].FF/Q OVHB\[7\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04924_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[27\].VALID\[12\].FF_D A[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12653_ _12665_/CLK line[67] vssd1 vssd1 vccd1 vccd1 _12654_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12917__D line[74] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XDATA\[11\].CLKBUF\[0\] clk vssd1 vssd1 vccd1 vccd1 _05527_/CLK sky130_fd_sc_hd__clkbuf_4
XPHY_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11821__D line[71] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11604_ _11604_/A _11619_/Y vssd1 vssd1 vccd1 vccd1 _13844_/Z sky130_fd_sc_hd__ebufn_2
XPHY_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06915__D line[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12584_ _12584_/A _12599_/Y vssd1 vssd1 vccd1 vccd1 _13704_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_196_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11535_ _11545_/CLK line[68] vssd1 vssd1 vccd1 vccd1 _11536_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11466_ _11466_/A _11479_/Y vssd1 vssd1 vccd1 vccd1 _13706_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13748__D line[56] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13205_ _13225_/CLK line[78] vssd1 vssd1 vccd1 vccd1 _13206_/A sky130_fd_sc_hd__dfxtp_1
X_10417_ _10425_/CLK line[69] vssd1 vssd1 vccd1 vccd1 _10418_/A sky130_fd_sc_hd__dfxtp_1
X_11397_ _11405_/CLK line[5] vssd1 vssd1 vccd1 vccd1 _11398_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06650__D line[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13136_ _13136_/A _13159_/Y vssd1 vssd1 vccd1 vccd1 _13696_/Z sky130_fd_sc_hd__ebufn_2
X_10348_ _10348_/A _10359_/Y vssd1 vssd1 vccd1 vccd1 _13708_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_151_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10172__D line[85] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10279_ _10285_/CLK line[6] vssd1 vssd1 vccd1 vccd1 _10280_/A sky130_fd_sc_hd__dfxtp_1
X_13067_ _13085_/CLK line[15] vssd1 vssd1 vccd1 vccd1 _13068_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05266__D line[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[21\].CG_CLK clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05844__A _13902_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12018_ _12018_/A _12039_/Y vssd1 vssd1 vccd1 vccd1 _13698_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_38_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13483__D line[77] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05563__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08577__D line[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07481__D line[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XOVHB\[13\].INV _13947_/X vssd1 vssd1 vccd1 vccd1 OVHB\[13\].INV/Y sky130_fd_sc_hd__inv_2
XANTENNA__12099__D line[70] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13969_ _13971_/B _13971_/A _13971_/C _13971_/D vssd1 vssd1 vccd1 vccd1 _13969_/X
+ sky130_fd_sc_hd__and4b_4
XFILLER_53_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06510_ _06540_/CLK line[80] vssd1 vssd1 vccd1 vccd1 _06511_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_207_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07490_ _07520_/CLK line[16] vssd1 vssd1 vccd1 vccd1 _07491_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[14\].VALID\[13\].TOBUF OVHB\[14\].VALID\[13\].FF/Q OVHB\[14\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04916_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_206_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06441_ _06441_/A _06474_/Y vssd1 vssd1 vccd1 vccd1 _13721_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_21_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_DATA\[16\].CLKBUF\[7\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XOVHB\[28\].INV _13968_/X vssd1 vssd1 vccd1 vccd1 OVHB\[28\].INV/Y sky130_fd_sc_hd__inv_2
XANTENNA__11731__D line[44] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09160_ _09160_/A _09169_/Y vssd1 vssd1 vccd1 vccd1 _13640_/Z sky130_fd_sc_hd__ebufn_2
X_06372_ _06400_/CLK line[26] vssd1 vssd1 vccd1 vccd1 _06373_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[4\].VALID\[12\].FF OVHB\[4\].V/CLK A[19] vssd1 vssd1 vccd1 vccd1 OVHB\[4\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__06825__D line[96] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08111_ _08115_/CLK line[39] vssd1 vssd1 vccd1 vccd1 _08112_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_30_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05323_ _05323_/A _05354_/Y vssd1 vssd1 vccd1 vccd1 _13723_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10347__D line[37] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09091_ _09095_/CLK line[103] vssd1 vssd1 vccd1 vccd1 _09092_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[20\].VALID\[8\].FF_D A[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08042_ _08042_/A _08049_/Y vssd1 vssd1 vccd1 vccd1 _13642_/Z sky130_fd_sc_hd__ebufn_2
X_05254_ _05280_/CLK line[27] vssd1 vssd1 vccd1 vccd1 _05255_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13658__D line[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05738__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05185_ _05185_/A _05214_/Y vssd1 vssd1 vccd1 vccd1 _13865_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07656__D line[87] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09993_ _10005_/CLK line[3] vssd1 vssd1 vccd1 vccd1 _09994_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_88_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10082__D line[58] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08944_ _08944_/A _08959_/Y vssd1 vssd1 vccd1 vccd1 _13704_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[9\].CLKBUF\[7\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08875_ _08885_/CLK line[4] vssd1 vssd1 vccd1 vccd1 _08876_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_69_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11906__D line[124] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10810__D line[121] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07826_ _07826_/A _07839_/Y vssd1 vssd1 vccd1 vccd1 _13706_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05904__D line[54] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07391__D line[108] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_04969_ _13931_/Y vssd1 vssd1 vccd1 vccd1 _04969_/Y sky130_fd_sc_hd__inv_2
X_07757_ _07765_/CLK line[5] vssd1 vssd1 vccd1 vccd1 _07758_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_37_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06708_ _06708_/A _06719_/Y vssd1 vssd1 vccd1 vccd1 _13708_/Z sky130_fd_sc_hd__ebufn_2
X_07688_ _07688_/A _07699_/Y vssd1 vssd1 vccd1 vccd1 _13848_/Z sky130_fd_sc_hd__ebufn_2
X_09427_ _09445_/CLK line[15] vssd1 vssd1 vccd1 vccd1 _09428_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[31\].CLKBUF\[0\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06639_ _06645_/CLK line[6] vssd1 vssd1 vccd1 vccd1 _06640_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_100_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09358_ _09358_/A _09379_/Y vssd1 vssd1 vccd1 vccd1 _13838_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10257__D line[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08309_ _08325_/CLK line[1] vssd1 vssd1 vccd1 vccd1 _08310_/A sky130_fd_sc_hd__dfxtp_1
X_09289_ _09305_/CLK line[65] vssd1 vssd1 vccd1 vccd1 _09290_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_126_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11320_ _11320_/A _11339_/Y vssd1 vssd1 vccd1 vccd1 _13840_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[28\].VALID\[10\].FF OVHB\[28\].V/CLK A[17] vssd1 vssd1 vccd1 vccd1 OVHB\[28\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11251_ _11265_/CLK line[66] vssd1 vssd1 vccd1 vccd1 _11252_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_109_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12472__D line[127] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07566__D line[60] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06470__D line[57] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10202_ _10202_/A _10219_/Y vssd1 vssd1 vccd1 vccd1 _13842_/Z sky130_fd_sc_hd__ebufn_2
X_11182_ _11182_/A _11199_/Y vssd1 vssd1 vccd1 vccd1 _13702_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_192_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11088__D line[120] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10133_ _10145_/CLK line[67] vssd1 vssd1 vccd1 vccd1 _10134_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[5\].VALID\[5\].TOBUF OVHB\[5\].VALID\[5\].FF/Q OVHB\[5\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04927_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_0_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09781__D line[34] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10064_ _10064_/A _10079_/Y vssd1 vssd1 vccd1 vccd1 _13704_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[1\].VALID\[3\].FF_D A[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10720__D line[94] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05814__D line[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13823_ _13899_/X wr vssd1 vssd1 vccd1 vccd1 _13823_/X sky130_fd_sc_hd__and2_1
XFILLER_28_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13754_ _13899_/X vssd1 vssd1 vccd1 vccd1 _13754_/Y sky130_fd_sc_hd__inv_2
X_10966_ _10966_/A _10989_/Y vssd1 vssd1 vccd1 vccd1 _13766_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_189_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12705_ _12735_/CLK line[96] vssd1 vssd1 vccd1 vccd1 _12706_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[18\].VALID\[12\].FF OVHB\[18\].V/CLK A[19] vssd1 vssd1 vccd1 vccd1 OVHB\[18\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_16_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12647__D line[79] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13685_ _13715_/CLK line[32] vssd1 vssd1 vccd1 vccd1 _13686_/A sky130_fd_sc_hd__dfxtp_1
X_10897_ _10915_/CLK line[47] vssd1 vssd1 vccd1 vccd1 _10898_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_188_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07103__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06645__D line[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12636_ _12636_/A _12669_/Y vssd1 vssd1 vccd1 vccd1 _13756_/Z sky130_fd_sc_hd__ebufn_2
XPHY_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09021__D line[71] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12567_ _12595_/CLK line[42] vssd1 vssd1 vccd1 vccd1 _12568_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09956__D line[114] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11518_ _11518_/A _11549_/Y vssd1 vssd1 vccd1 vccd1 _13758_/Z sky130_fd_sc_hd__ebufn_2
X_12498_ _12498_/A _12529_/Y vssd1 vssd1 vccd1 vccd1 _13618_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_156_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11449_ _11475_/CLK line[43] vssd1 vssd1 vccd1 vccd1 _11450_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06380__D line[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13119_ _13119_/A _13124_/Y vssd1 vssd1 vccd1 vccd1 _13679_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_98_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06990_ _06990_/A _06999_/Y vssd1 vssd1 vccd1 vccd1 _13710_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_79_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05941_ _05945_/CLK line[71] vssd1 vssd1 vccd1 vccd1 _05942_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_85_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05872_ _05872_/A _05879_/Y vssd1 vssd1 vccd1 vccd1 _13712_/Z sky130_fd_sc_hd__ebufn_2
X_08660_ _08660_/A _08679_/Y vssd1 vssd1 vccd1 vccd1 _13700_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_66_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07611_ _07625_/CLK line[66] vssd1 vssd1 vccd1 vccd1 _07612_/A sky130_fd_sc_hd__dfxtp_1
X_08591_ _08605_/CLK line[2] vssd1 vssd1 vccd1 vccd1 _08592_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_53_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07542_ _07542_/A _07559_/Y vssd1 vssd1 vccd1 vccd1 _13702_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[12\].VALID\[0\].TOBUF OVHB\[12\].VALID\[0\].FF/Q OVHB\[12\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04924_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__04918__A A_h[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07473_ _07485_/CLK line[3] vssd1 vssd1 vccd1 vccd1 _07474_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[16\].VALID\[0\].FF_D A[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XMUX.SEL0BUF\[1\] A[0] vssd1 vssd1 vccd1 vccd1 MUX.SEL0BUF\[1\]/X sky130_fd_sc_hd__clkbuf_2
XFILLER_179_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11461__D line[34] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09212_ _09212_/A _09239_/Y vssd1 vssd1 vccd1 vccd1 _13692_/Z sky130_fd_sc_hd__ebufn_2
X_06424_ _06424_/A _06439_/Y vssd1 vssd1 vccd1 vccd1 _13704_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06555__D line[110] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09143_ _09165_/CLK line[13] vssd1 vssd1 vccd1 vccd1 _09144_/A sky130_fd_sc_hd__dfxtp_1
X_06355_ _06365_/CLK line[4] vssd1 vssd1 vccd1 vccd1 _06356_/A sky130_fd_sc_hd__dfxtp_1
X_05306_ _05306_/A _05319_/Y vssd1 vssd1 vccd1 vccd1 _13706_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08770__D line[84] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09074_ _09074_/A _09099_/Y vssd1 vssd1 vccd1 vccd1 _13834_/Z sky130_fd_sc_hd__ebufn_2
X_06286_ _06286_/A _06299_/Y vssd1 vssd1 vccd1 vccd1 _13846_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13388__D line[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08025_ _08045_/CLK line[14] vssd1 vssd1 vccd1 vccd1 _08026_/A sky130_fd_sc_hd__dfxtp_1
X_05237_ _05245_/CLK line[5] vssd1 vssd1 vccd1 vccd1 _05238_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_162_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05168_ _05168_/A _05179_/Y vssd1 vssd1 vccd1 vccd1 _13848_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[10\].CLKBUF\[0\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09976_ _09976_/A _10009_/Y vssd1 vssd1 vccd1 vccd1 _13616_/Z sky130_fd_sc_hd__ebufn_2
X_05099_ _05105_/CLK line[70] vssd1 vssd1 vccd1 vccd1 _05100_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_39_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08927_ _08955_/CLK line[42] vssd1 vssd1 vccd1 vccd1 _08928_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11636__D line[114] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDATA\[3\].CLKBUF\[7\] clk vssd1 vssd1 vccd1 vccd1 _12212_/CLK sky130_fd_sc_hd__clkbuf_4
X_08858_ _08858_/A _08889_/Y vssd1 vssd1 vccd1 vccd1 _13618_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09106__D line[124] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11933__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[0\].VALID\[10\].FF OVHB\[0\].V/CLK A[17] vssd1 vssd1 vccd1 vccd1 OVHB\[0\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_07809_ _07835_/CLK line[43] vssd1 vssd1 vccd1 vccd1 _07810_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08010__D line[121] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[7\].VALID\[7\].FF_D A[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08789_ _08815_/CLK line[107] vssd1 vssd1 vccd1 vccd1 _08790_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_26_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13851__D line[103] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10820_ _10820_/A _10849_/Y vssd1 vssd1 vccd1 vccd1 _13620_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08945__D line[36] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10751_ _10775_/CLK line[108] vssd1 vssd1 vccd1 vccd1 _10752_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[3\].CLKBUF\[0\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13470_ _13470_/CLK line[57] vssd1 vssd1 vccd1 vccd1 _13471_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_40_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10682_ _10682_/A _10709_/Y vssd1 vssd1 vccd1 vccd1 _13762_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_139_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12421_ _12421_/A _12424_/Y vssd1 vssd1 vccd1 vccd1 _13821_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08680__D line[48] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12352_ _12352_/CLK _12353_/X vssd1 vssd1 vccd1 vccd1 _12350_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_5_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11303_ _13933_/X wr vssd1 vssd1 vccd1 vccd1 _11303_/X sky130_fd_sc_hd__and2_1
X_12283_ _13935_/X wr vssd1 vssd1 vccd1 vccd1 _12283_/X sky130_fd_sc_hd__and2_1
XANTENNA__07296__D line[50] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07874__A _13912_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11234_ _13933_/X vssd1 vssd1 vccd1 vccd1 _11234_/Y sky130_fd_sc_hd__inv_2
XANTENNA__07593__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11165_ _11195_/CLK line[32] vssd1 vssd1 vccd1 vccd1 _11166_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_96_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10116_ _10116_/A _10149_/Y vssd1 vssd1 vccd1 vccd1 _13756_/Z sky130_fd_sc_hd__ebufn_2
X_11096_ _11096_/A _11129_/Y vssd1 vssd1 vccd1 vccd1 _13616_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[8\].VALID\[10\].TOBUF OVHB\[8\].VALID\[10\].FF/Q OVHB\[8\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04932_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_0_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10450__D line[84] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10047_ _10075_/CLK line[42] vssd1 vssd1 vccd1 vccd1 _10048_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[16\].CG clk OVHB\[16\].CGAND/X vssd1 vssd1 vccd1 vccd1 OVHB\[16\].V/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_208_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05544__D line[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_MUX.M\[0\].MUX\[6\]_A3 _13850_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13761__D line[76] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13806_ _13820_/CLK line[82] vssd1 vssd1 vccd1 vccd1 _13807_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[29\].VALID\[0\].FF_D A[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08855__D line[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11998_ _12000_/CLK line[24] vssd1 vssd1 vccd1 vccd1 _11999_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[2\].CLKBUF\[4\] clk vssd1 vssd1 vccd1 vccd1 _11267_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__12377__D line[69] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13737_ _13737_/A _13754_/Y vssd1 vssd1 vccd1 vccd1 _13737_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_44_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10949_ _10949_/A _10954_/Y vssd1 vssd1 vccd1 vccd1 _13749_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_188_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13668_ _13680_/CLK line[19] vssd1 vssd1 vccd1 vccd1 _13669_/A sky130_fd_sc_hd__dfxtp_1
XPHY_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12619_ _12619_/A _12634_/Y vssd1 vssd1 vccd1 vccd1 _13739_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_31_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07768__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13599_ _13599_/A _13614_/Y vssd1 vssd1 vccd1 vccd1 _13879_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09686__D line[119] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06140_ _06140_/A _06159_/Y vssd1 vssd1 vccd1 vccd1 _13700_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_184_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06071_ _06085_/CLK line[2] vssd1 vssd1 vccd1 vccd1 _06072_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10625__D line[36] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13001__D line[98] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05719__D line[97] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05022_ _05022_/A _05039_/Y vssd1 vssd1 vccd1 vccd1 _13702_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[10\].VALID\[5\].TOBUF OVHB\[10\].VALID\[5\].FF/Q OVHB\[10\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04927_/B2 sky130_fd_sc_hd__ebufn_2
XDEC.DEC0.AND2 A[5] A[6] vssd1 vssd1 vccd1 vccd1 _13916_/D sky130_fd_sc_hd__and2b_2
XANTENNA__12840__D line[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09830_ _09830_/CLK line[57] vssd1 vssd1 vccd1 vccd1 _09831_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07934__D line[86] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09761_ _09761_/A _09764_/Y vssd1 vssd1 vccd1 vccd1 _13681_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_100_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06973_ _06995_/CLK line[45] vssd1 vssd1 vccd1 vccd1 _06974_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_39_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XOVHB\[14\].VALID\[10\].FF OVHB\[14\].V/CLK A[17] vssd1 vssd1 vccd1 vccd1 OVHB\[14\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_08712_ _08712_/CLK _08713_/X vssd1 vssd1 vccd1 vccd1 _08710_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__10360__D line[48] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05924_ _05924_/A _05949_/Y vssd1 vssd1 vccd1 vccd1 _13764_/Z sky130_fd_sc_hd__ebufn_2
X_09692_ _09692_/CLK _09693_/X vssd1 vssd1 vccd1 vccd1 _09690_/CLK sky130_fd_sc_hd__dlclkp_1
X_08643_ _13914_/X wr vssd1 vssd1 vccd1 vccd1 _08643_/X sky130_fd_sc_hd__and2_1
X_05855_ _05875_/CLK line[46] vssd1 vssd1 vccd1 vccd1 _05856_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08574_ _13913_/X vssd1 vssd1 vccd1 vccd1 _08574_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05786_ _05786_/A _05809_/Y vssd1 vssd1 vccd1 vccd1 _13626_/Z sky130_fd_sc_hd__ebufn_2
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07525_ _07555_/CLK line[32] vssd1 vssd1 vccd1 vccd1 _07526_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12287__D line[42] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11191__D line[39] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06285__D line[100] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07456_ _07456_/A _07489_/Y vssd1 vssd1 vccd1 vccd1 _13616_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XDATA\[1\].CLKBUF\[1\] clk vssd1 vssd1 vccd1 vccd1 _08082_/CLK sky130_fd_sc_hd__clkbuf_4
X_06407_ _06435_/CLK line[42] vssd1 vssd1 vccd1 vccd1 _06408_/A sky130_fd_sc_hd__dfxtp_1
X_07387_ _07415_/CLK line[106] vssd1 vssd1 vccd1 vccd1 _07388_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09596__D line[92] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[28\].CLKBUF\[3\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09126_ _09130_/CLK line[119] vssd1 vssd1 vccd1 vccd1 _09127_/A sky130_fd_sc_hd__dfxtp_1
X_06338_ _06338_/A _06369_/Y vssd1 vssd1 vccd1 vccd1 _13618_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[21\].V_RESET_B rst_n vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__04932__A2_N _04932_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10535__D line[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09057_ _09057_/A _09064_/Y vssd1 vssd1 vccd1 vccd1 _13817_/Z sky130_fd_sc_hd__ebufn_2
X_06269_ _06295_/CLK line[107] vssd1 vssd1 vccd1 vccd1 _06270_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_135_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08008_ _08010_/CLK line[120] vssd1 vssd1 vccd1 vccd1 _08009_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12750__D line[126] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07844__D line[59] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09959_ _09959_/A _09974_/Y vssd1 vssd1 vccd1 vccd1 _13879_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11366__D line[119] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12970_ _12980_/CLK line[84] vssd1 vssd1 vccd1 vccd1 _12971_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_181_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11921_ _11921_/A _11934_/Y vssd1 vssd1 vccd1 vccd1 _13881_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09414__A _13916_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11852_ _11860_/CLK line[85] vssd1 vssd1 vccd1 vccd1 _11853_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08675__D line[41] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09133__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDATA\[21\].CLKBUF\[5\] clk vssd1 vssd1 vccd1 vccd1 _08782_/CLK sky130_fd_sc_hd__clkbuf_4
X_10803_ _10803_/A _10814_/Y vssd1 vssd1 vccd1 vccd1 _13883_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_60_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11783_ _11783_/A _11794_/Y vssd1 vssd1 vccd1 vccd1 _13743_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_201_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06195__D line[64] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13522_ _13540_/CLK line[95] vssd1 vssd1 vccd1 vccd1 _13523_/A sky130_fd_sc_hd__dfxtp_1
X_10734_ _10740_/CLK line[86] vssd1 vssd1 vccd1 vccd1 _10735_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_41_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[19\].VALID\[0\].TOBUF OVHB\[19\].VALID\[0\].FF/Q OVHB\[19\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04924_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_158_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_DECH.DEC0.AND0_A A_h[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12925__D line[78] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13453_ _13453_/A _13474_/Y vssd1 vssd1 vccd1 vccd1 _13733_/Z sky130_fd_sc_hd__ebufn_2
X_10665_ _10665_/A _10674_/Y vssd1 vssd1 vccd1 vccd1 _13745_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_185_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05389__A _13900_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12404_ _12420_/CLK line[81] vssd1 vssd1 vccd1 vccd1 _12405_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06923__D line[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13384_ _13400_/CLK line[17] vssd1 vssd1 vccd1 vccd1 _13385_/A sky130_fd_sc_hd__dfxtp_1
X_10596_ _10600_/CLK line[23] vssd1 vssd1 vccd1 vccd1 _10597_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_182_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12335_ _12335_/A _12354_/Y vssd1 vssd1 vccd1 vccd1 _13735_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[1\].CLKBUF\[2\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12266_ _12280_/CLK line[18] vssd1 vssd1 vccd1 vccd1 _12267_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_141_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XOVHB\[24\].VALID\[11\].TOBUF OVHB\[24\].VALID\[11\].FF/Q OVHB\[24\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04915_/B2 sky130_fd_sc_hd__ebufn_2
X_11217_ _11217_/A _11234_/Y vssd1 vssd1 vccd1 vccd1 _13737_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09308__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12197_ _12197_/A _12214_/Y vssd1 vssd1 vccd1 vccd1 _13877_/Z sky130_fd_sc_hd__ebufn_2
X_11148_ _11160_/CLK line[19] vssd1 vssd1 vccd1 vccd1 _11149_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_110_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11276__D line[92] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10180__D line[89] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11079_ _11079_/A _11094_/Y vssd1 vssd1 vccd1 vccd1 _13879_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05274__D line[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13491__D line[66] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[9\].VALID\[12\].FF OVHB\[9\].V/CLK A[19] vssd1 vssd1 vccd1 vccd1 OVHB\[9\].VALID\[12\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__08585__D line[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05640_ _05640_/A _05669_/Y vssd1 vssd1 vccd1 vccd1 _13760_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[12\].VALID\[3\].FF_D A[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05571_ _05595_/CLK line[44] vssd1 vssd1 vccd1 vccd1 _05572_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_205_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07310_ _07310_/CLK line[57] vssd1 vssd1 vccd1 vccd1 _07311_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_32_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06683__A _13905_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08290_ _08290_/CLK line[121] vssd1 vssd1 vccd1 vccd1 _08291_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_31_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XDATA\[20\].CLKBUF\[2\] clk vssd1 vssd1 vccd1 vccd1 _08397_/CLK sky130_fd_sc_hd__clkbuf_4
X_07241_ _07241_/A _07244_/Y vssd1 vssd1 vccd1 vccd1 _13681_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_165_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07172_ _07172_/CLK _07173_/X vssd1 vssd1 vccd1 vccd1 _07170_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__06833__D line[109] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06123_ _13903_/X wr vssd1 vssd1 vccd1 vccd1 _06123_/X sky130_fd_sc_hd__and2_1
XANTENNA__10355__D line[41] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05449__D line[102] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06054_ _13902_/X vssd1 vssd1 vccd1 vccd1 _06054_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13666__D line[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05005_ _05035_/CLK line[32] vssd1 vssd1 vccd1 vccd1 _05006_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_160_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09813_ _09813_/A _09834_/Y vssd1 vssd1 vccd1 vccd1 _13733_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_100_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10090__D line[62] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09744_ _09760_/CLK line[17] vssd1 vssd1 vccd1 vccd1 _09745_/A sky130_fd_sc_hd__dfxtp_1
X_06956_ _06960_/CLK line[23] vssd1 vssd1 vccd1 vccd1 _06957_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06858__A _13905_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05184__D line[123] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05907_ _05907_/A _05914_/Y vssd1 vssd1 vccd1 vccd1 _13747_/Z sky130_fd_sc_hd__ebufn_2
X_09675_ _09675_/A _09694_/Y vssd1 vssd1 vccd1 vccd1 _13875_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_39_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06887_ _06887_/A _06894_/Y vssd1 vssd1 vccd1 vccd1 _13887_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11914__D line[113] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08626_ _08640_/CLK line[18] vssd1 vssd1 vccd1 vccd1 _08627_/A sky130_fd_sc_hd__dfxtp_1
X_05838_ _05840_/CLK line[24] vssd1 vssd1 vccd1 vccd1 _05839_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08557_ _08557_/A _08574_/Y vssd1 vssd1 vccd1 vccd1 _13877_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05769_ _05769_/A _05774_/Y vssd1 vssd1 vccd1 vccd1 _13889_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07508_ _07520_/CLK line[19] vssd1 vssd1 vccd1 vccd1 _07509_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08488_ _08500_/CLK line[83] vssd1 vssd1 vccd1 vccd1 _08489_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07439_ _07439_/A _07454_/Y vssd1 vssd1 vccd1 vccd1 _13879_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[4\].VALID\[12\].FF_D A[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XOVHB\[20\].VALID\[1\].FF OVHB\[20\].V/CLK A[8] vssd1 vssd1 vccd1 vccd1 OVHB\[20\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_6_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10450_ _10460_/CLK line[84] vssd1 vssd1 vccd1 vccd1 _10451_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_182_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10265__D line[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09109_ _09109_/A _09134_/Y vssd1 vssd1 vccd1 vccd1 _13869_/Z sky130_fd_sc_hd__ebufn_2
X_10381_ _10381_/A _10394_/Y vssd1 vssd1 vccd1 vccd1 _13741_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05359__D line[75] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12120_ _12140_/CLK line[94] vssd1 vssd1 vccd1 vccd1 _12121_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12480__D line[116] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[26\].CLKBUF\[5\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12051_ _12051_/A _12074_/Y vssd1 vssd1 vccd1 vccd1 _13731_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07574__D line[49] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11002_ _11020_/CLK line[95] vssd1 vssd1 vccd1 vccd1 _11003_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_77_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[17\].VALID\[5\].TOBUF OVHB\[17\].VALID\[5\].FF/Q OVHB\[17\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04927_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_92_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[25\].VALID\[3\].FF_D A[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12953_ _12953_/A _12984_/Y vssd1 vssd1 vccd1 vccd1 _13793_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_85_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11904_ _11930_/CLK line[123] vssd1 vssd1 vccd1 vccd1 _11905_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_18_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12884_ _12910_/CLK line[59] vssd1 vssd1 vccd1 vccd1 _12885_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05822__D line[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11835_ _11835_/A _11864_/Y vssd1 vssd1 vccd1 vccd1 _13795_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09798__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[3\].CGAND_B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[18\].VALID\[7\].FF_D A[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[22\].CGAND_A _13915_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11766_ _11790_/CLK line[60] vssd1 vssd1 vccd1 vccd1 _11767_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13505_ _13505_/CLK line[73] vssd1 vssd1 vccd1 vccd1 _13506_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[19\].VALID\[2\].FF OVHB\[19\].V/CLK A[9] vssd1 vssd1 vccd1 vccd1 OVHB\[19\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_10717_ _10717_/A _10744_/Y vssd1 vssd1 vccd1 vccd1 _13797_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12655__D line[68] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11697_ _11697_/A _11724_/Y vssd1 vssd1 vccd1 vccd1 _13657_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07749__D line[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[7\].CGAND_A _13938_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13436_ _13436_/A _13439_/Y vssd1 vssd1 vccd1 vccd1 _13716_/Z sky130_fd_sc_hd__ebufn_2
X_10648_ _10670_/CLK line[61] vssd1 vssd1 vccd1 vccd1 _10649_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_6_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13367_ _13367_/CLK _13368_/X vssd1 vssd1 vccd1 vccd1 _13365_/CLK sky130_fd_sc_hd__dlclkp_1
X_10579_ _10579_/A _10604_/Y vssd1 vssd1 vccd1 vccd1 _13659_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09964__D line[118] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12318_ _13935_/X wr vssd1 vssd1 vccd1 vccd1 _12318_/X sky130_fd_sc_hd__and2_1
XFILLER_181_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08223__A _13932_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13298_ _13938_/X wr vssd1 vssd1 vccd1 vccd1 _13298_/X sky130_fd_sc_hd__and2_1
XANTENNA__10903__D line[35] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12390__D line[80] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12249_ _13935_/X vssd1 vssd1 vccd1 vccd1 _12249_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11584__A _13926_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06810_ _06820_/CLK line[84] vssd1 vssd1 vccd1 vccd1 _06811_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_68_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07790_ _07800_/CLK line[20] vssd1 vssd1 vccd1 vccd1 _07791_/A sky130_fd_sc_hd__dfxtp_1
X_06741_ _06741_/A _06754_/Y vssd1 vssd1 vccd1 vccd1 _13741_/Z sky130_fd_sc_hd__ebufn_2
X_09460_ _09480_/CLK line[30] vssd1 vssd1 vccd1 vccd1 _09461_/A sky130_fd_sc_hd__dfxtp_1
X_06672_ _06680_/CLK line[21] vssd1 vssd1 vccd1 vccd1 _06673_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_52_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08411_ _08411_/A _08434_/Y vssd1 vssd1 vccd1 vccd1 _13731_/Z sky130_fd_sc_hd__ebufn_2
X_05623_ _05623_/A _05634_/Y vssd1 vssd1 vccd1 vccd1 _13743_/Z sky130_fd_sc_hd__ebufn_2
X_09391_ _09391_/A _09414_/Y vssd1 vssd1 vccd1 vccd1 _13871_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[23\].VALID\[4\].TOBUF OVHB\[23\].VALID\[4\].FF/Q OVHB\[23\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04925_/B2 sky130_fd_sc_hd__ebufn_2
X_08342_ _08360_/CLK line[31] vssd1 vssd1 vccd1 vccd1 _08343_/A sky130_fd_sc_hd__dfxtp_1
X_05554_ _05560_/CLK line[22] vssd1 vssd1 vccd1 vccd1 _05555_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_149_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12565__D line[32] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05485_ _05485_/A _05494_/Y vssd1 vssd1 vccd1 vccd1 _13885_/Z sky130_fd_sc_hd__ebufn_2
X_08273_ _08273_/A _08294_/Y vssd1 vssd1 vccd1 vccd1 _13873_/Z sky130_fd_sc_hd__ebufn_2
X_07224_ _07240_/CLK line[17] vssd1 vssd1 vccd1 vccd1 _07225_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06563__D line[99] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11759__A _13927_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07155_ _07155_/A _07174_/Y vssd1 vssd1 vccd1 vccd1 _13875_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_106_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09874__D line[91] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06106_ _06120_/CLK line[18] vssd1 vssd1 vccd1 vccd1 _06107_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11478__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07086_ _07100_/CLK line[82] vssd1 vssd1 vccd1 vccd1 _07087_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[17\].VALID\[4\].FF OVHB\[17\].V/CLK A[11] vssd1 vssd1 vccd1 vccd1 OVHB\[17\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_160_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13396__D line[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13974__A A_h[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06037_ _06037_/A _06054_/Y vssd1 vssd1 vccd1 vccd1 _13877_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_154_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XOVHB\[5\].VALID\[10\].FF OVHB\[5\].V/CLK A[17] vssd1 vssd1 vccd1 vccd1 OVHB\[5\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_113_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07988_ _08010_/CLK line[125] vssd1 vssd1 vccd1 vccd1 _07989_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_47_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09727_ _09727_/CLK _09728_/X vssd1 vssd1 vccd1 vccd1 _09725_/CLK sky130_fd_sc_hd__dlclkp_1
X_06939_ _06939_/A _06964_/Y vssd1 vssd1 vccd1 vccd1 _13659_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11644__D line[118] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09658_ _13920_/Y wr vssd1 vssd1 vccd1 vccd1 _09658_/X sky130_fd_sc_hd__and2_1
XFILLER_27_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06738__D line[51] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09114__D line[113] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08609_ _13914_/X vssd1 vssd1 vccd1 vccd1 _08609_/Y sky130_fd_sc_hd__inv_2
XPHY_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09589_ _13920_/Y vssd1 vssd1 vccd1 vccd1 _09589_/Y sky130_fd_sc_hd__inv_2
XPHY_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11620_ _11650_/CLK line[112] vssd1 vssd1 vccd1 vccd1 _11621_/A sky130_fd_sc_hd__dfxtp_1
XPHY_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08953__D line[40] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11551_ _11551_/A _11584_/Y vssd1 vssd1 vccd1 vccd1 _13791_/Z sky130_fd_sc_hd__ebufn_2
XPHY_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10502_ _10530_/CLK line[122] vssd1 vssd1 vccd1 vccd1 _10503_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11482_ _11510_/CLK line[58] vssd1 vssd1 vccd1 vccd1 _11483_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13221_ _13225_/CLK line[71] vssd1 vssd1 vccd1 vccd1 _13222_/A sky130_fd_sc_hd__dfxtp_1
X_10433_ _10433_/A _10464_/Y vssd1 vssd1 vccd1 vccd1 _13793_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05089__D line[65] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13152_ _13152_/A _13159_/Y vssd1 vssd1 vccd1 vccd1 _13712_/Z sky130_fd_sc_hd__ebufn_2
X_10364_ _10390_/CLK line[59] vssd1 vssd1 vccd1 vccd1 _10365_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11819__D line[70] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12103_ _12105_/CLK line[72] vssd1 vssd1 vccd1 vccd1 _12104_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_88_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13083_ _13085_/CLK line[8] vssd1 vssd1 vccd1 vccd1 _13084_/A sky130_fd_sc_hd__dfxtp_1
X_10295_ _10295_/A _10324_/Y vssd1 vssd1 vccd1 vccd1 _13655_/Z sky130_fd_sc_hd__ebufn_2
X_12034_ _12034_/A _12039_/Y vssd1 vssd1 vccd1 vccd1 _13714_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_78_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XOVHB\[15\].VALID\[6\].FF OVHB\[15\].V/CLK A[13] vssd1 vssd1 vccd1 vccd1 OVHB\[15\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_DATA\[24\].CLKBUF\[7\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11554__D line[91] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12936_ _12936_/A _12949_/Y vssd1 vssd1 vccd1 vccd1 _13776_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_19_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05552__D line[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12867_ _12875_/CLK line[37] vssd1 vssd1 vccd1 vccd1 _12868_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13124__A _13938_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08863__D line[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11818_ _11818_/A _11829_/Y vssd1 vssd1 vccd1 vccd1 _13778_/Z sky130_fd_sc_hd__ebufn_2
X_12798_ _12798_/A _12809_/Y vssd1 vssd1 vccd1 vccd1 _13638_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12385__D line[73] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11749_ _11755_/CLK line[38] vssd1 vssd1 vccd1 vccd1 _11750_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07479__D line[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05270_ _05280_/CLK line[20] vssd1 vssd1 vccd1 vccd1 _05271_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_128_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13419_ _13435_/CLK line[33] vssd1 vssd1 vccd1 vccd1 _13420_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_127_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XOVHB\[19\].VALID\[10\].FF OVHB\[19\].V/CLK A[17] vssd1 vssd1 vccd1 vccd1 OVHB\[19\].VALID\[10\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11729__D line[43] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10633__D line[40] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08960_ _08990_/CLK line[48] vssd1 vssd1 vccd1 vccd1 _08961_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08888__A _13915_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05727__D line[101] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07911_ _07911_/A _07944_/Y vssd1 vssd1 vccd1 vccd1 _13791_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08103__D line[35] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[21\].VALID\[9\].TOBUF OVHB\[21\].VALID\[9\].FF/Q OVHB\[21\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04914_/B2 sky130_fd_sc_hd__ebufn_2
X_08891_ _08891_/A _08924_/Y vssd1 vssd1 vccd1 vccd1 _13651_/Z sky130_fd_sc_hd__ebufn_2
X_07842_ _07870_/CLK line[58] vssd1 vssd1 vccd1 vccd1 _07843_/A sky130_fd_sc_hd__dfxtp_1
X_07773_ _07773_/A _07804_/Y vssd1 vssd1 vccd1 vccd1 _13653_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13018__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_04985_ _04985_/A _05004_/Y vssd1 vssd1 vccd1 vccd1 _13665_/Z sky130_fd_sc_hd__ebufn_2
X_09512_ _09512_/A _09519_/Y vssd1 vssd1 vccd1 vccd1 _13712_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_17_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06724_ _06750_/CLK line[59] vssd1 vssd1 vccd1 vccd1 _06725_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05462__D line[122] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09443_ _09445_/CLK line[8] vssd1 vssd1 vccd1 vccd1 _09444_/A sky130_fd_sc_hd__dfxtp_1
X_06655_ _06655_/A _06684_/Y vssd1 vssd1 vccd1 vccd1 _13655_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_197_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05606_ _05630_/CLK line[60] vssd1 vssd1 vccd1 vccd1 _05607_/A sky130_fd_sc_hd__dfxtp_1
X_09374_ _09374_/A _09379_/Y vssd1 vssd1 vccd1 vccd1 _13854_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[13\].VALID\[8\].FF OVHB\[13\].V/CLK A[15] vssd1 vssd1 vccd1 vccd1 OVHB\[13\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06586_ _06610_/CLK line[124] vssd1 vssd1 vccd1 vccd1 _06587_/A sky130_fd_sc_hd__dfxtp_1
X_08325_ _08325_/CLK line[9] vssd1 vssd1 vccd1 vccd1 _08326_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12295__D line[46] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10808__D line[120] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05537_ _05537_/A _05564_/Y vssd1 vssd1 vccd1 vccd1 _13657_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07389__D line[107] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06293__D line[104] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08256_ _08256_/A _08259_/Y vssd1 vssd1 vccd1 vccd1 _13856_/Z sky130_fd_sc_hd__ebufn_2
X_05468_ _05490_/CLK line[125] vssd1 vssd1 vccd1 vccd1 _05469_/A sky130_fd_sc_hd__dfxtp_1
X_07207_ _07207_/CLK _07208_/X vssd1 vssd1 vccd1 vccd1 _07205_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__10393__A _13923_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08187_ _08187_/CLK _08188_/X vssd1 vssd1 vccd1 vccd1 _08185_/CLK sky130_fd_sc_hd__dlclkp_1
X_05399_ _05399_/A _05424_/Y vssd1 vssd1 vccd1 vccd1 _13799_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_152_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07138_ _13909_/Y wr vssd1 vssd1 vccd1 vccd1 _07138_/X sky130_fd_sc_hd__and2_1
XFILLER_3_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10543__D line[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07069_ _13909_/Y vssd1 vssd1 vccd1 vccd1 _07069_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05637__D line[74] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10080_ _10110_/CLK line[48] vssd1 vssd1 vccd1 vccd1 _10081_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[21\].VALID\[6\].FF_D A[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07852__D line[63] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13770_ _13770_/A _13789_/Y vssd1 vssd1 vccd1 vccd1 _13770_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06468__D line[56] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10982_ _10982_/A _10989_/Y vssd1 vssd1 vccd1 vccd1 _13782_/Z sky130_fd_sc_hd__ebufn_2
X_12721_ _12735_/CLK line[98] vssd1 vssd1 vccd1 vccd1 _12722_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_204_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10568__A _13924_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09779__D line[33] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12652_ _12652_/A _12669_/Y vssd1 vssd1 vccd1 vccd1 _13772_/Z sky130_fd_sc_hd__ebufn_2
XPHY_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[5\].VALID\[1\].TOBUF OVHB\[5\].VALID\[1\].FF/Q OVHB\[5\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04926_/B2 sky130_fd_sc_hd__ebufn_2
XPHY_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11603_ _11615_/CLK line[99] vssd1 vssd1 vccd1 vccd1 _11604_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10718__D line[93] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12583_ _12595_/CLK line[35] vssd1 vssd1 vccd1 vccd1 _12584_/A sky130_fd_sc_hd__dfxtp_1
XPHY_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11534_ _11534_/A _11549_/Y vssd1 vssd1 vccd1 vccd1 _13774_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12933__D line[67] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11465_ _11475_/CLK line[36] vssd1 vssd1 vccd1 vccd1 _11466_/A sky130_fd_sc_hd__dfxtp_1
X_13204_ _13204_/A _13229_/Y vssd1 vssd1 vccd1 vccd1 _13764_/Z sky130_fd_sc_hd__ebufn_2
X_10416_ _10416_/A _10429_/Y vssd1 vssd1 vccd1 vccd1 _13776_/Z sky130_fd_sc_hd__ebufn_2
X_11396_ _11396_/A _11409_/Y vssd1 vssd1 vccd1 vccd1 _13636_/Z sky130_fd_sc_hd__ebufn_2
X_13135_ _13155_/CLK line[46] vssd1 vssd1 vccd1 vccd1 _13136_/A sky130_fd_sc_hd__dfxtp_1
X_10347_ _10355_/CLK line[37] vssd1 vssd1 vccd1 vccd1 _10348_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[11\].VALID\[14\].FF_D A[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09019__D line[70] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13066_ _13066_/A _13089_/Y vssd1 vssd1 vccd1 vccd1 _13626_/Z sky130_fd_sc_hd__ebufn_2
X_10278_ _10278_/A _10289_/Y vssd1 vssd1 vccd1 vccd1 _13638_/Z sky130_fd_sc_hd__ebufn_2
X_12017_ _12035_/CLK line[47] vssd1 vssd1 vccd1 vccd1 _12018_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[10\].VALID\[14\].TOBUF OVHB\[10\].VALID\[14\].FF/Q OVHB\[10\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_93_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11284__D line[81] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06378__D line[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13968_ _13971_/A _13971_/B _13971_/C _13971_/D vssd1 vssd1 vccd1 vccd1 _13968_/X
+ sky130_fd_sc_hd__and4bb_4
X_12919_ _12945_/CLK line[75] vssd1 vssd1 vccd1 vccd1 _12920_/A sky130_fd_sc_hd__dfxtp_1
X_13899_ _13905_/C _13905_/B _13905_/A _13905_/D vssd1 vssd1 vccd1 vccd1 _13899_/X
+ sky130_fd_sc_hd__and4bb_4
XFILLER_61_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[21\].VALID\[13\].FF_D A[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDATA\[30\].CLKBUF\[7\] clk vssd1 vssd1 vccd1 vccd1 _11652_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__08593__D line[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06440_ _06470_/CLK line[48] vssd1 vssd1 vccd1 vccd1 _06441_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_210_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[2\].VALID\[1\].FF_D A[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13789__A _13899_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06371_ _06371_/A _06404_/Y vssd1 vssd1 vccd1 vccd1 _13651_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08110_ _08110_/A _08119_/Y vssd1 vssd1 vccd1 vccd1 _13710_/Z sky130_fd_sc_hd__ebufn_2
X_05322_ _05350_/CLK line[58] vssd1 vssd1 vccd1 vccd1 _05323_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_119_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09090_ _09090_/A _09099_/Y vssd1 vssd1 vccd1 vccd1 _13850_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07002__D line[58] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08041_ _08045_/CLK line[7] vssd1 vssd1 vccd1 vccd1 _08042_/A sky130_fd_sc_hd__dfxtp_1
X_05253_ _05253_/A _05284_/Y vssd1 vssd1 vccd1 vccd1 _13653_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_162_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06841__D line[98] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05184_ _05210_/CLK line[123] vssd1 vssd1 vccd1 vccd1 _05185_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11459__D line[33] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[31\].VALID\[12\].FF_D A[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09992_ _09992_/A _10009_/Y vssd1 vssd1 vccd1 vccd1 _13632_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_88_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08943_ _08955_/CLK line[35] vssd1 vssd1 vccd1 vccd1 _08944_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13674__D line[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[23\].V_D TIE/HI vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08874_ _08874_/A _08889_/Y vssd1 vssd1 vccd1 vccd1 _13634_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08768__D line[83] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07825_ _07835_/CLK line[36] vssd1 vssd1 vccd1 vccd1 _07826_/A sky130_fd_sc_hd__dfxtp_1
X_07756_ _07756_/A _07769_/Y vssd1 vssd1 vccd1 vccd1 _13636_/Z sky130_fd_sc_hd__ebufn_2
X_04968_ _13931_/Y wr vssd1 vssd1 vccd1 vccd1 _04968_/X sky130_fd_sc_hd__and2_1
XANTENNA__05192__D line[127] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06707_ _06715_/CLK line[37] vssd1 vssd1 vccd1 vccd1 _06708_/A sky130_fd_sc_hd__dfxtp_1
X_07687_ _07695_/CLK line[101] vssd1 vssd1 vccd1 vccd1 _07688_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11922__D line[117] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09426_ _09426_/A _09449_/Y vssd1 vssd1 vccd1 vccd1 _13626_/Z sky130_fd_sc_hd__ebufn_2
X_06638_ _06638_/A _06649_/Y vssd1 vssd1 vccd1 vccd1 _13638_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_40_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_OVHB\[13\].VALID\[10\].FF_D A[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09357_ _09375_/CLK line[111] vssd1 vssd1 vccd1 vccd1 _09358_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_200_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06569_ _06575_/CLK line[102] vssd1 vssd1 vccd1 vccd1 _06570_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[6\].VALID\[1\].FF OVHB\[6\].V/CLK A[8] vssd1 vssd1 vccd1 vccd1 OVHB\[6\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_100_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08308_ _08308_/A _08329_/Y vssd1 vssd1 vccd1 vccd1 _13628_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08008__D line[120] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09288_ _09288_/A _09309_/Y vssd1 vssd1 vccd1 vccd1 _13768_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_60_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13849__D line[102] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08239_ _08255_/CLK line[97] vssd1 vssd1 vccd1 vccd1 _08240_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12108__A _13934_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[30\].VALID\[14\].TOBUF OVHB\[30\].VALID\[14\].FF/Q OVHB\[30\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_119_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11250_ _11250_/A _11269_/Y vssd1 vssd1 vccd1 vccd1 _13770_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_106_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10201_ _10215_/CLK line[98] vssd1 vssd1 vccd1 vccd1 _10202_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10273__D line[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11181_ _11195_/CLK line[34] vssd1 vssd1 vccd1 vccd1 _11182_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_134_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05367__D line[79] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10132_ _10132_/A _10149_/Y vssd1 vssd1 vccd1 vccd1 _13772_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_133_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13584__D line[123] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XOVHB\[3\].VALID\[6\].TOBUF OVHB\[3\].VALID\[6\].FF/Q OVHB\[3\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04923_/A2 sky130_fd_sc_hd__ebufn_2
XFILLER_125_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10063_ _10075_/CLK line[35] vssd1 vssd1 vccd1 vccd1 _10064_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07582__D line[53] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XOVHB\[28\].VALID\[9\].TOBUF OVHB\[28\].VALID\[9\].FF/Q OVHB\[28\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04914_/B2 sky130_fd_sc_hd__ebufn_2
X_13822_ _13822_/CLK _13823_/X vssd1 vssd1 vccd1 vccd1 _13820_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_63_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13753_ _13899_/X wr vssd1 vssd1 vccd1 vccd1 _13753_/X sky130_fd_sc_hd__and2_1
XFILLER_90_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10965_ _10985_/CLK line[78] vssd1 vssd1 vccd1 vccd1 _10966_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11832__D line[90] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12704_ _13936_/X vssd1 vssd1 vccd1 vccd1 _12704_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13684_ _13899_/X vssd1 vssd1 vccd1 vccd1 _13684_/Y sky130_fd_sc_hd__inv_2
XANTENNA__05830__D line[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10896_ _10896_/A _10919_/Y vssd1 vssd1 vccd1 vccd1 _13696_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_31_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12635_ _12665_/CLK line[64] vssd1 vssd1 vccd1 vccd1 _12636_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10448__D line[83] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_DATA\[17\].CLKBUF\[1\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12566_ _12566_/A _12599_/Y vssd1 vssd1 vccd1 vccd1 _13686_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[8\].VALID\[5\].FF_D A[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13759__D line[75] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11517_ _11545_/CLK line[74] vssd1 vssd1 vccd1 vccd1 _11518_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12663__D line[72] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12497_ _12525_/CLK line[10] vssd1 vssd1 vccd1 vccd1 _12498_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07757__D line[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11448_ _11448_/A _11479_/Y vssd1 vssd1 vccd1 vccd1 _13688_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_144_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XOVHB\[4\].VALID\[3\].FF OVHB\[4\].V/CLK A[10] vssd1 vssd1 vccd1 vccd1 OVHB\[4\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_171_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11379_ _11405_/CLK line[11] vssd1 vssd1 vccd1 vccd1 _11380_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_113_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13118_ _13120_/CLK line[24] vssd1 vssd1 vccd1 vccd1 _13119_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_79_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05940_ _05940_/A _05949_/Y vssd1 vssd1 vccd1 vccd1 _13780_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10911__D line[39] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13049_ _13049_/A _13054_/Y vssd1 vssd1 vccd1 vccd1 _13889_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07492__D line[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05871_ _05875_/CLK line[39] vssd1 vssd1 vccd1 vccd1 _05872_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_94_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07610_ _07610_/A _07629_/Y vssd1 vssd1 vccd1 vccd1 _13770_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_93_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08590_ _08590_/A _08609_/Y vssd1 vssd1 vccd1 vccd1 _13630_/Z sky130_fd_sc_hd__ebufn_2
X_07541_ _07555_/CLK line[34] vssd1 vssd1 vccd1 vccd1 _07542_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12838__D line[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[10\].VALID\[1\].TOBUF OVHB\[10\].VALID\[1\].FF/Q OVHB\[10\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04926_/B2 sky130_fd_sc_hd__ebufn_2
X_07472_ _07472_/A _07489_/Y vssd1 vssd1 vccd1 vccd1 _13632_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05740__D line[112] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09211_ _09235_/CLK line[44] vssd1 vssd1 vccd1 vccd1 _09212_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_195_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06423_ _06435_/CLK line[35] vssd1 vssd1 vccd1 vccd1 _06424_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_179_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09142_ _09142_/A _09169_/Y vssd1 vssd1 vccd1 vccd1 _13622_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[8\].V_D TIE/HI vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06354_ _06354_/A _06369_/Y vssd1 vssd1 vccd1 vccd1 _13634_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[20\].V_RESET_B rst_n vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05305_ _05315_/CLK line[36] vssd1 vssd1 vccd1 vccd1 _05306_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12573__D line[45] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09073_ _09095_/CLK line[109] vssd1 vssd1 vccd1 vccd1 _09074_/A sky130_fd_sc_hd__dfxtp_1
X_06285_ _06295_/CLK line[100] vssd1 vssd1 vccd1 vccd1 _06286_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07667__D line[106] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08024_ _08024_/A _08049_/Y vssd1 vssd1 vccd1 vccd1 _13624_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06571__D line[103] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05236_ _05236_/A _05249_/Y vssd1 vssd1 vccd1 vccd1 _13636_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_146_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11189__D line[38] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05167_ _05175_/CLK line[101] vssd1 vssd1 vccd1 vccd1 _05168_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09882__D line[95] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09975_ _10005_/CLK line[0] vssd1 vssd1 vccd1 vccd1 _09976_/A sky130_fd_sc_hd__dfxtp_1
X_05098_ _05098_/A _05109_/Y vssd1 vssd1 vccd1 vccd1 _13778_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_131_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10821__D line[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08926_ _08926_/A _08959_/Y vssd1 vssd1 vccd1 vccd1 _13686_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08498__D line[88] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[18\].VALID\[14\].FF_D A[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05915__D line[64] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08857_ _08885_/CLK line[10] vssd1 vssd1 vccd1 vccd1 _08858_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[2\].VALID\[5\].FF OVHB\[2\].V/CLK A[12] vssd1 vssd1 vccd1 vccd1 OVHB\[2\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12598__A _13936_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07808_ _07808_/A _07839_/Y vssd1 vssd1 vccd1 vccd1 _13688_/Z sky130_fd_sc_hd__ebufn_2
X_08788_ _08788_/A _08819_/Y vssd1 vssd1 vccd1 vccd1 _13828_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_55_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07739_ _07765_/CLK line[11] vssd1 vssd1 vccd1 vccd1 _07740_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12748__D line[125] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__04932__B1 A_h[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10750_ _10750_/A _10779_/Y vssd1 vssd1 vccd1 vccd1 _13830_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06746__D line[55] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09122__D line[117] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09409_ _09409_/A _09414_/Y vssd1 vssd1 vccd1 vccd1 _13889_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_52_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10681_ _10705_/CLK line[76] vssd1 vssd1 vccd1 vccd1 _10682_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_139_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[28\].VALID\[13\].FF_D A[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12420_ _12420_/CLK line[89] vssd1 vssd1 vccd1 vccd1 _12421_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_185_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12351_ _12351_/A _12354_/Y vssd1 vssd1 vccd1 vccd1 _13751_/Z sky130_fd_sc_hd__ebufn_2
X_11302_ _11302_/CLK _11303_/X vssd1 vssd1 vccd1 vccd1 _11300_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__06481__D line[76] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12282_ _12282_/CLK _12283_/X vssd1 vssd1 vccd1 vccd1 _12280_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_4_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[12\].INV _13946_/X vssd1 vssd1 vccd1 vccd1 OVHB\[12\].INV/Y sky130_fd_sc_hd__inv_2
XOVHB\[4\].VALID\[11\].TOBUF OVHB\[4\].VALID\[11\].FF/Q OVHB\[4\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04915_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__11099__D line[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11233_ _13933_/X wr vssd1 vssd1 vccd1 vccd1 _11233_/X sky130_fd_sc_hd__and2_1
XFILLER_153_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05097__D line[69] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11164_ _13933_/X vssd1 vssd1 vccd1 vccd1 _11164_/Y sky130_fd_sc_hd__inv_2
X_10115_ _10145_/CLK line[64] vssd1 vssd1 vccd1 vccd1 _10116_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[27\].INV _13967_/X vssd1 vssd1 vccd1 vccd1 OVHB\[27\].INV/Y sky130_fd_sc_hd__inv_2
XFILLER_110_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11095_ _11125_/CLK line[0] vssd1 vssd1 vccd1 vccd1 _11096_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_88_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10046_ _10046_/A _10079_/Y vssd1 vssd1 vccd1 vccd1 _13686_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_209_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13805_ _13805_/A _13824_/Y vssd1 vssd1 vccd1 vccd1 _13805_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_91_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11562__D line[95] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11997_ _11997_/A _12004_/Y vssd1 vssd1 vccd1 vccd1 _13677_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06656__D line[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13736_ _13750_/CLK line[50] vssd1 vssd1 vccd1 vccd1 _13737_/A sky130_fd_sc_hd__dfxtp_1
X_10948_ _10950_/CLK line[56] vssd1 vssd1 vccd1 vccd1 _10949_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_16_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05560__D line[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[0\].VALID\[7\].FF OVHB\[0\].V/CLK A[14] vssd1 vssd1 vccd1 vccd1 OVHB\[0\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__09032__D line[90] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10178__D line[88] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10879_ _10879_/A _10884_/Y vssd1 vssd1 vccd1 vccd1 _13679_/Z sky130_fd_sc_hd__ebufn_2
X_13667_ _13667_/A _13684_/Y vssd1 vssd1 vccd1 vccd1 _13667_/Z sky130_fd_sc_hd__ebufn_2
XPHY_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08871__D line[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12618_ _12630_/CLK line[51] vssd1 vssd1 vccd1 vccd1 _12619_/A sky130_fd_sc_hd__dfxtp_1
XPHY_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13598_ _13610_/CLK line[115] vssd1 vssd1 vccd1 vccd1 _13599_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13489__D line[65] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12549_ _12549_/A _12564_/Y vssd1 vssd1 vccd1 vccd1 _13669_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_6_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06070_ _06070_/A _06089_/Y vssd1 vssd1 vccd1 vccd1 _13630_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[30\].VALID\[9\].FF_D A[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05021_ _05035_/CLK line[34] vssd1 vssd1 vccd1 vccd1 _05022_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_132_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_DATA\[15\].CLKBUF\[3\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XDEC.DEC0.AND3 A[6] A[5] vssd1 vssd1 vccd1 vccd1 _13927_/D sky130_fd_sc_hd__and2_2
XOVHB\[29\].VALID\[0\].FF OVHB\[29\].V/CLK A[7] vssd1 vssd1 vccd1 vccd1 OVHB\[29\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11737__D line[47] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09760_ _09760_/CLK line[25] vssd1 vssd1 vccd1 vccd1 _09761_/A sky130_fd_sc_hd__dfxtp_1
X_06972_ _06972_/A _06999_/Y vssd1 vssd1 vccd1 vccd1 _13692_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_98_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_MUX.M\[2\].MUX\[0\]_A0 _13651_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09207__D line[42] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05735__D line[105] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08711_ _08711_/A _08714_/Y vssd1 vssd1 vccd1 vccd1 _13751_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_67_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05923_ _05945_/CLK line[77] vssd1 vssd1 vccd1 vccd1 _05924_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08111__D line[39] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09691_ _09691_/A _09694_/Y vssd1 vssd1 vccd1 vccd1 _13891_/Z sky130_fd_sc_hd__ebufn_2
X_08642_ _08642_/CLK _08643_/X vssd1 vssd1 vccd1 vccd1 _08640_/CLK sky130_fd_sc_hd__dlclkp_1
X_05854_ _05854_/A _05879_/Y vssd1 vssd1 vccd1 vccd1 _13694_/Z sky130_fd_sc_hd__ebufn_2
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08573_ _13913_/X wr vssd1 vssd1 vccd1 vccd1 _08573_/X sky130_fd_sc_hd__and2_1
XPHY_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05785_ _05805_/CLK line[14] vssd1 vssd1 vccd1 vccd1 _05786_/A sky130_fd_sc_hd__dfxtp_1
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07524_ _13911_/X vssd1 vssd1 vccd1 vccd1 _07524_/Y sky130_fd_sc_hd__inv_2
XPHY_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05470__D line[126] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_DATA\[8\].CLKBUF\[3\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10088__D line[61] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07455_ _07485_/CLK line[0] vssd1 vssd1 vccd1 vccd1 _07456_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06406_ _06406_/A _06439_/Y vssd1 vssd1 vccd1 vccd1 _13686_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_41_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07386_ _07386_/A _07419_/Y vssd1 vssd1 vccd1 vccd1 _13826_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_182_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09125_ _09125_/A _09134_/Y vssd1 vssd1 vccd1 vccd1 _13885_/Z sky130_fd_sc_hd__ebufn_2
X_06337_ _06365_/CLK line[10] vssd1 vssd1 vccd1 vccd1 _06338_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[13\].VALID\[1\].FF_D A[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07397__D line[111] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09056_ _09060_/CLK line[87] vssd1 vssd1 vccd1 vccd1 _09057_/A sky130_fd_sc_hd__dfxtp_1
X_06268_ _06268_/A _06299_/Y vssd1 vssd1 vccd1 vccd1 _13828_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_163_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08007_ _08007_/A _08014_/Y vssd1 vssd1 vccd1 vccd1 _13887_/Z sky130_fd_sc_hd__ebufn_2
X_05219_ _05245_/CLK line[11] vssd1 vssd1 vccd1 vccd1 _05220_/A sky130_fd_sc_hd__dfxtp_1
X_06199_ _06225_/CLK line[75] vssd1 vssd1 vccd1 vccd1 _06200_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[27\].VALID\[13\].TOBUF OVHB\[27\].VALID\[13\].FF/Q OVHB\[27\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04916_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_131_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10551__D line[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09958_ _09970_/CLK line[115] vssd1 vssd1 vccd1 vccd1 _09959_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05645__D line[78] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08021__D line[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08909_ _08909_/A _08924_/Y vssd1 vssd1 vccd1 vccd1 _13669_/Z sky130_fd_sc_hd__ebufn_2
X_09889_ _09889_/A _09904_/Y vssd1 vssd1 vccd1 vccd1 _13809_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13862__D line[122] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11920_ _11930_/CLK line[116] vssd1 vssd1 vccd1 vccd1 _11921_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07860__D line[52] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XOVHB\[27\].VALID\[2\].FF OVHB\[27\].V/CLK A[9] vssd1 vssd1 vccd1 vccd1 OVHB\[27\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11851_ _11851_/A _11864_/Y vssd1 vssd1 vccd1 vccd1 _13811_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12478__D line[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10802_ _10810_/CLK line[117] vssd1 vssd1 vccd1 vccd1 _10803_/A sky130_fd_sc_hd__dfxtp_1
X_11782_ _11790_/CLK line[53] vssd1 vssd1 vccd1 vccd1 _11783_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_53_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10733_ _10733_/A _10744_/Y vssd1 vssd1 vccd1 vccd1 _13813_/Z sky130_fd_sc_hd__ebufn_2
X_13521_ _13521_/A _13544_/Y vssd1 vssd1 vccd1 vccd1 _13801_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[4\].VALID\[8\].FF_D A[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09787__D line[37] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DECH.DEC0.AND0_B A_h[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13452_ _13470_/CLK line[63] vssd1 vssd1 vccd1 vccd1 _13453_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[17\].VALID\[1\].TOBUF OVHB\[17\].VALID\[1\].FF/Q OVHB\[17\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04926_/B2 sky130_fd_sc_hd__ebufn_2
X_10664_ _10670_/CLK line[54] vssd1 vssd1 vccd1 vccd1 _10665_/A sky130_fd_sc_hd__dfxtp_1
X_12403_ _12403_/A _12424_/Y vssd1 vssd1 vccd1 vccd1 _13803_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10726__D line[82] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[20\].VALID\[12\].TOBUF OVHB\[20\].VALID\[12\].FF/Q OVHB\[20\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04929_/B2 sky130_fd_sc_hd__ebufn_2
X_13383_ _13383_/A _13404_/Y vssd1 vssd1 vccd1 vccd1 _13663_/Z sky130_fd_sc_hd__ebufn_2
X_10595_ _10595_/A _10604_/Y vssd1 vssd1 vccd1 vccd1 _13675_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13102__D line[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12334_ _12350_/CLK line[49] vssd1 vssd1 vccd1 vccd1 _12335_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_31_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07100__D line[89] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12265_ _12265_/A _12284_/Y vssd1 vssd1 vccd1 vccd1 _13665_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12941__D line[71] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11216_ _11230_/CLK line[50] vssd1 vssd1 vccd1 vccd1 _11217_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_107_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12196_ _12210_/CLK line[114] vssd1 vssd1 vccd1 vccd1 _12197_/A sky130_fd_sc_hd__dfxtp_1
X_11147_ _11147_/A _11164_/Y vssd1 vssd1 vccd1 vccd1 _13667_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_95_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11078_ _11090_/CLK line[115] vssd1 vssd1 vccd1 vccd1 _11079_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_48_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10029_ _10029_/A _10044_/Y vssd1 vssd1 vccd1 vccd1 _13669_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_64_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07770__D line[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11292__D line[85] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06386__D line[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05570_ _05570_/A _05599_/Y vssd1 vssd1 vccd1 vccd1 _13690_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_17_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06964__A _13909_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13719_ _13899_/X vssd1 vssd1 vccd1 vccd1 _13719_/Y sky130_fd_sc_hd__inv_2
XANTENNA__06683__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09697__D line[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[26\].VALID\[1\].FF_D A[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07240_ _07240_/CLK line[25] vssd1 vssd1 vccd1 vccd1 _07241_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[25\].VALID\[4\].FF OVHB\[25\].V/CLK A[11] vssd1 vssd1 vccd1 vccd1 OVHB\[25\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_20_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07171_ _07171_/A _07174_/Y vssd1 vssd1 vccd1 vccd1 _13891_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_118_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06122_ _06122_/CLK _06123_/X vssd1 vssd1 vccd1 vccd1 _06120_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_117_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XDATA\[19\].CLKBUF\[0\] clk vssd1 vssd1 vccd1 vccd1 _07767_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__07010__D line[62] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12851__D line[44] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06053_ _13902_/X wr vssd1 vssd1 vccd1 vccd1 _06053_/X sky130_fd_sc_hd__and2_1
XANTENNA_OVHB\[19\].VALID\[5\].FF_D A[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07945__D line[96] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05004_ _13931_/Y vssd1 vssd1 vccd1 vccd1 _05004_/Y sky130_fd_sc_hd__inv_2
XOVHB\[23\].VALID\[0\].TOBUF OVHB\[23\].VALID\[0\].FF/Q OVHB\[23\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04924_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__11467__D line[37] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09812_ _09830_/CLK line[63] vssd1 vssd1 vccd1 vccd1 _09813_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_140_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06955_ _06955_/A _06964_/Y vssd1 vssd1 vccd1 vccd1 _13675_/Z sky130_fd_sc_hd__ebufn_2
X_09743_ _09743_/A _09764_/Y vssd1 vssd1 vccd1 vccd1 _13663_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[13\].CLKBUF\[5\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06858__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05906_ _05910_/CLK line[55] vssd1 vssd1 vccd1 vccd1 _05907_/A sky130_fd_sc_hd__dfxtp_1
X_09674_ _09690_/CLK line[113] vssd1 vssd1 vccd1 vccd1 _09675_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08776__D line[87] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06886_ _06890_/CLK line[119] vssd1 vssd1 vccd1 vccd1 _06887_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08625_ _08625_/A _08644_/Y vssd1 vssd1 vccd1 vccd1 _13665_/Z sky130_fd_sc_hd__ebufn_2
X_05837_ _05837_/A _05844_/Y vssd1 vssd1 vccd1 vccd1 _13677_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08556_ _08570_/CLK line[114] vssd1 vssd1 vccd1 vccd1 _08557_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05768_ _05770_/CLK line[120] vssd1 vssd1 vccd1 vccd1 _05769_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07507_ _07507_/A _07524_/Y vssd1 vssd1 vccd1 vccd1 _13667_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_52_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08487_ _08487_/A _08504_/Y vssd1 vssd1 vccd1 vccd1 _13807_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11930__D line[121] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05699_ _05699_/A _05704_/Y vssd1 vssd1 vccd1 vccd1 _13819_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07438_ _07450_/CLK line[115] vssd1 vssd1 vccd1 vccd1 _07439_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09400__D line[116] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07369_ _07369_/A _07384_/Y vssd1 vssd1 vccd1 vccd1 _13809_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_176_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_DATA\[6\].CLKBUF\[5\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09108_ _09130_/CLK line[125] vssd1 vssd1 vccd1 vccd1 _09109_/A sky130_fd_sc_hd__dfxtp_1
X_10380_ _10390_/CLK line[52] vssd1 vssd1 vccd1 vccd1 _10381_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_136_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09039_ _09039_/A _09064_/Y vssd1 vssd1 vccd1 vccd1 _13799_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[23\].VALID\[6\].FF OVHB\[23\].V/CLK A[13] vssd1 vssd1 vccd1 vccd1 OVHB\[23\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_151_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12050_ _12070_/CLK line[62] vssd1 vssd1 vccd1 vccd1 _12051_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_104_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11377__D line[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11001_ _11001_/A _11024_/Y vssd1 vssd1 vccd1 vccd1 _13801_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10281__D line[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05375__D line[68] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XOVHB\[15\].VALID\[6\].TOBUF OVHB\[15\].VALID\[6\].FF/Q OVHB\[15\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04923_/A2 sky130_fd_sc_hd__ebufn_2
XANTENNA__13592__D line[127] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08686__D line[60] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12952_ _12980_/CLK line[90] vssd1 vssd1 vccd1 vccd1 _12953_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_206_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07590__D line[57] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11903_ _11903_/A _11934_/Y vssd1 vssd1 vccd1 vccd1 _13863_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_206_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12883_ _12883_/A _12914_/Y vssd1 vssd1 vccd1 vccd1 _13723_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_61_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11834_ _11860_/CLK line[91] vssd1 vssd1 vccd1 vccd1 _11835_/A sky130_fd_sc_hd__dfxtp_1
X_11765_ _11765_/A _11794_/Y vssd1 vssd1 vccd1 vccd1 _13725_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11840__D line[94] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[22\].CGAND_B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10716_ _10740_/CLK line[92] vssd1 vssd1 vccd1 vccd1 _10717_/A sky130_fd_sc_hd__dfxtp_1
X_13504_ _13504_/A _13509_/Y vssd1 vssd1 vccd1 vccd1 _13784_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_158_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06934__D line[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11696_ _11720_/CLK line[28] vssd1 vssd1 vccd1 vccd1 _11697_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09310__D line[80] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10456__D line[87] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[26\].CGAND_A _13922_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13435_ _13435_/CLK line[41] vssd1 vssd1 vccd1 vccd1 _13436_/A sky130_fd_sc_hd__dfxtp_1
X_10647_ _10647_/A _10674_/Y vssd1 vssd1 vccd1 vccd1 _13727_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_139_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[7\].CGAND_B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[15\].CG_CLK clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13366_ _13366_/A _13369_/Y vssd1 vssd1 vccd1 vccd1 _13646_/Z sky130_fd_sc_hd__ebufn_2
X_10578_ _10600_/CLK line[29] vssd1 vssd1 vccd1 vccd1 _10579_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08504__A _13913_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13767__D line[79] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12317_ _12317_/CLK _12318_/X vssd1 vssd1 vccd1 vccd1 _12315_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_154_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13297_ _13297_/CLK _13298_/X vssd1 vssd1 vccd1 vccd1 _13295_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__07765__D line[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08223__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12248_ _13935_/X wr vssd1 vssd1 vccd1 vccd1 _12248_/X sky130_fd_sc_hd__and2_1
XANTENNA__10191__D line[108] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12179_ _13934_/X vssd1 vssd1 vccd1 vccd1 _12179_/Y sky130_fd_sc_hd__inv_2
XANTENNA__05285__D line[32] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06740_ _06750_/CLK line[52] vssd1 vssd1 vccd1 vccd1 _06741_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[21\].VALID\[8\].FF OVHB\[21\].V/CLK A[15] vssd1 vssd1 vccd1 vccd1 OVHB\[21\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_92_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__04931__A2_N _04931_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06671_ _06671_/A _06684_/Y vssd1 vssd1 vccd1 vccd1 _13671_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13007__D line[101] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08410_ _08430_/CLK line[62] vssd1 vssd1 vccd1 vccd1 _08411_/A sky130_fd_sc_hd__dfxtp_1
X_05622_ _05630_/CLK line[53] vssd1 vssd1 vccd1 vccd1 _05623_/A sky130_fd_sc_hd__dfxtp_1
X_09390_ _09410_/CLK line[126] vssd1 vssd1 vccd1 vccd1 _09391_/A sky130_fd_sc_hd__dfxtp_1
X_08341_ _08341_/A _08364_/Y vssd1 vssd1 vccd1 vccd1 _13661_/Z sky130_fd_sc_hd__ebufn_2
X_05553_ _05553_/A _05564_/Y vssd1 vssd1 vccd1 vccd1 _13673_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_177_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XOVHB\[21\].VALID\[5\].TOBUF OVHB\[21\].VALID\[5\].FF/Q OVHB\[21\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04927_/B2 sky130_fd_sc_hd__ebufn_2
XOVHB\[29\].CG clk OVHB\[29\].CGAND/X vssd1 vssd1 vccd1 vccd1 OVHB\[29\].V/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_149_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08272_ _08290_/CLK line[127] vssd1 vssd1 vccd1 vccd1 _08273_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_20_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05484_ _05490_/CLK line[118] vssd1 vssd1 vccd1 vccd1 _05485_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_177_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07223_ _07223_/A _07244_/Y vssd1 vssd1 vccd1 vccd1 _13663_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_149_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10366__D line[60] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07154_ _07170_/CLK line[113] vssd1 vssd1 vccd1 vccd1 _07155_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_145_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06105_ _06105_/A _06124_/Y vssd1 vssd1 vccd1 vccd1 _13665_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12581__D line[34] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07085_ _07085_/A _07104_/Y vssd1 vssd1 vccd1 vccd1 _13805_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07675__D line[110] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06036_ _06050_/CLK line[114] vssd1 vssd1 vccd1 vccd1 _06037_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_160_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09890__D line[84] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05773__A _13901_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07987_ _07987_/A _08014_/Y vssd1 vssd1 vccd1 vccd1 _13867_/Z sky130_fd_sc_hd__ebufn_2
X_09726_ _09726_/A _09729_/Y vssd1 vssd1 vccd1 vccd1 _13646_/Z sky130_fd_sc_hd__ebufn_2
X_06938_ _06960_/CLK line[29] vssd1 vssd1 vccd1 vccd1 _06939_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05923__D line[77] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06869_ _06869_/A _06894_/Y vssd1 vssd1 vccd1 vccd1 _13869_/Z sky130_fd_sc_hd__ebufn_2
X_09657_ _09657_/CLK _09658_/X vssd1 vssd1 vccd1 vccd1 _09655_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_55_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08608_ _13914_/X wr vssd1 vssd1 vccd1 vccd1 _08608_/X sky130_fd_sc_hd__and2_1
XFILLER_188_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09588_ _13920_/Y wr vssd1 vssd1 vccd1 vccd1 _09588_/X sky130_fd_sc_hd__and2_1
XPHY_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_DATA\[11\].CLKBUF\[7\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08539_ _13913_/X vssd1 vssd1 vccd1 vccd1 _08539_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12756__D line[114] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11550_ _11580_/CLK line[80] vssd1 vssd1 vccd1 vccd1 _11551_/A sky130_fd_sc_hd__dfxtp_1
XPHY_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09130__D line[121] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10501_ _10501_/A _10534_/Y vssd1 vssd1 vccd1 vccd1 _13861_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11481_ _11481_/A _11514_/Y vssd1 vssd1 vccd1 vccd1 _13721_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13220_ _13220_/A _13229_/Y vssd1 vssd1 vccd1 vccd1 _13780_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05948__A _13902_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10432_ _10460_/CLK line[90] vssd1 vssd1 vccd1 vccd1 _10433_/A sky130_fd_sc_hd__dfxtp_1
X_13151_ _13155_/CLK line[39] vssd1 vssd1 vccd1 vccd1 _13152_/A sky130_fd_sc_hd__dfxtp_1
X_10363_ _10363_/A _10394_/Y vssd1 vssd1 vccd1 vccd1 _13723_/Z sky130_fd_sc_hd__ebufn_2
X_12102_ _12102_/A _12109_/Y vssd1 vssd1 vccd1 vccd1 _13782_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[17\].VALID\[11\].TOBUF OVHB\[17\].VALID\[11\].FF/Q OVHB\[17\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04915_/B2 sky130_fd_sc_hd__ebufn_2
X_13082_ _13082_/A _13089_/Y vssd1 vssd1 vccd1 vccd1 _13642_/Z sky130_fd_sc_hd__ebufn_2
X_10294_ _10320_/CLK line[27] vssd1 vssd1 vccd1 vccd1 _10295_/A sky130_fd_sc_hd__dfxtp_1
X_12033_ _12035_/CLK line[40] vssd1 vssd1 vccd1 vccd1 _12034_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_DATA\[4\].CLKBUF\[7\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08994__A _13915_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09305__D line[73] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12935_ _12945_/CLK line[68] vssd1 vssd1 vccd1 vccd1 _12936_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_18_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12866_ _12866_/A _12879_/Y vssd1 vssd1 vccd1 vccd1 _13706_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[22\].VALID\[4\].FF_D A[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11817_ _11825_/CLK line[69] vssd1 vssd1 vccd1 vccd1 _11818_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_159_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11570__D line[84] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12797_ _12805_/CLK line[5] vssd1 vssd1 vccd1 vccd1 _12798_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06664__D line[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11748_ _11748_/A _11759_/Y vssd1 vssd1 vccd1 vccd1 _13708_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06019__A _13902_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09040__D line[94] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[10\].VALID\[10\].TOBUF OVHB\[10\].VALID\[10\].FF/Q OVHB\[10\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04932_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_159_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11679_ _11685_/CLK line[6] vssd1 vssd1 vccd1 vccd1 _11680_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09975__D line[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13418_ _13418_/A _13439_/Y vssd1 vssd1 vccd1 vccd1 _13698_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[15\].VALID\[8\].FF_D A[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13497__D line[69] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MUX.M\[3\].MUX\[2\]_A0 _13653_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13349_ _13365_/CLK line[1] vssd1 vssd1 vccd1 vccd1 _13350_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08888__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07910_ _07940_/CLK line[80] vssd1 vssd1 vccd1 vccd1 _07911_/A sky130_fd_sc_hd__dfxtp_1
X_08890_ _08920_/CLK line[16] vssd1 vssd1 vccd1 vccd1 _08891_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_69_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07841_ _07841_/A _07874_/Y vssd1 vssd1 vccd1 vccd1 _13721_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_69_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11745__D line[36] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07772_ _07800_/CLK line[26] vssd1 vssd1 vccd1 vccd1 _07773_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06839__D line[97] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_04984_ _05000_/CLK line[17] vssd1 vssd1 vccd1 vccd1 _04985_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_68_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09215__D line[46] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09511_ _09515_/CLK line[39] vssd1 vssd1 vccd1 vccd1 _09512_/A sky130_fd_sc_hd__dfxtp_1
X_06723_ _06723_/A _06754_/Y vssd1 vssd1 vccd1 vccd1 _13723_/Z sky130_fd_sc_hd__ebufn_2
X_09442_ _09442_/A _09449_/Y vssd1 vssd1 vccd1 vccd1 _13642_/Z sky130_fd_sc_hd__ebufn_2
X_06654_ _06680_/CLK line[27] vssd1 vssd1 vccd1 vccd1 _06655_/A sky130_fd_sc_hd__dfxtp_1
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07313__A _13910_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05605_ _05605_/A _05634_/Y vssd1 vssd1 vccd1 vccd1 _13725_/Z sky130_fd_sc_hd__ebufn_2
X_09373_ _09375_/CLK line[104] vssd1 vssd1 vccd1 vccd1 _09374_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_197_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06585_ _06585_/A _06614_/Y vssd1 vssd1 vccd1 vccd1 _13865_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11480__D line[48] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08324_ _08324_/A _08329_/Y vssd1 vssd1 vccd1 vccd1 _13644_/Z sky130_fd_sc_hd__ebufn_2
X_05536_ _05560_/CLK line[28] vssd1 vssd1 vccd1 vccd1 _05537_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_20_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10096__D line[50] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08255_ _08255_/CLK line[105] vssd1 vssd1 vccd1 vccd1 _08256_/A sky130_fd_sc_hd__dfxtp_1
X_05467_ _05467_/A _05494_/Y vssd1 vssd1 vccd1 vccd1 _13867_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10674__A _13924_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07206_ _07206_/A _07209_/Y vssd1 vssd1 vccd1 vccd1 _13646_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[5\].VALID\[13\].FF_D A[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08186_ _08186_/A _08189_/Y vssd1 vssd1 vccd1 vccd1 _13786_/Z sky130_fd_sc_hd__ebufn_2
X_05398_ _05420_/CLK line[93] vssd1 vssd1 vccd1 vccd1 _05399_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_180_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10393__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07137_ _07137_/CLK _07138_/X vssd1 vssd1 vccd1 vccd1 _07135_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_106_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07068_ _13909_/Y wr vssd1 vssd1 vccd1 vccd1 _07068_/X sky130_fd_sc_hd__and2_1
XFILLER_0_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06019_ _13902_/X vssd1 vssd1 vccd1 vccd1 _06019_/Y sky130_fd_sc_hd__inv_2
XANTENNA_MUX.SEL0BUF\[1\]_A A[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11655__D line[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05653__D line[67] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XOVHB\[30\].VALID\[10\].TOBUF OVHB\[30\].VALID\[10\].FF/Q OVHB\[30\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04932_/B2 sky130_fd_sc_hd__ebufn_2
X_09709_ _09725_/CLK line[1] vssd1 vssd1 vccd1 vccd1 _09710_/A sky130_fd_sc_hd__dfxtp_1
X_10981_ _10985_/CLK line[71] vssd1 vssd1 vccd1 vccd1 _10982_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_90_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10849__A _13925_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13870__D line[126] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[25\].CLKBUF\[1\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12720_ _12720_/A _12739_/Y vssd1 vssd1 vccd1 vccd1 _13840_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08964__D line[59] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10568__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12486__D line[119] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12651_ _12665_/CLK line[66] vssd1 vssd1 vccd1 vccd1 _12652_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11602_ _11602_/A _11619_/Y vssd1 vssd1 vccd1 vccd1 _13842_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12582_ _12582_/A _12599_/Y vssd1 vssd1 vccd1 vccd1 _13702_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_168_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XOVHB\[3\].VALID\[2\].TOBUF OVHB\[3\].VALID\[2\].FF/Q OVHB\[3\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04930_/B2 sky130_fd_sc_hd__ebufn_2
XPHY_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[28\].VALID\[8\].FF_D A[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11533_ _11545_/CLK line[67] vssd1 vssd1 vccd1 vccd1 _11534_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[28\].VALID\[5\].TOBUF OVHB\[28\].VALID\[5\].FF/Q OVHB\[28\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04927_/B2 sky130_fd_sc_hd__ebufn_2
XPHY_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09795__D line[41] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11464_ _11464_/A _11479_/Y vssd1 vssd1 vccd1 vccd1 _13704_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_139_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10415_ _10425_/CLK line[68] vssd1 vssd1 vccd1 vccd1 _10416_/A sky130_fd_sc_hd__dfxtp_1
X_13203_ _13225_/CLK line[77] vssd1 vssd1 vccd1 vccd1 _13204_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13895__A A[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10734__D line[86] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11395_ _11405_/CLK line[4] vssd1 vssd1 vccd1 vccd1 _11396_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13110__D line[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05828__D line[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[27\].VOBUF OVHB\[27\].V/Q OVHB\[27\].INV/Y vssd1 vssd1 vccd1 vccd1 _04912_/B1
+ sky130_fd_sc_hd__ebufn_2
XDATA\[9\].CLKBUF\[1\] clk vssd1 vssd1 vccd1 vccd1 _13682_/CLK sky130_fd_sc_hd__clkbuf_4
X_10346_ _10346_/A _10359_/Y vssd1 vssd1 vccd1 vccd1 _13706_/Z sky130_fd_sc_hd__ebufn_2
X_13134_ _13134_/A _13159_/Y vssd1 vssd1 vccd1 vccd1 _13694_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_151_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08204__D line[81] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13065_ _13085_/CLK line[14] vssd1 vssd1 vccd1 vccd1 _13066_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_3_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10277_ _10285_/CLK line[5] vssd1 vssd1 vccd1 vccd1 _10278_/A sky130_fd_sc_hd__dfxtp_1
X_12016_ _12016_/A _12039_/Y vssd1 vssd1 vccd1 vccd1 _13696_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_47_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13967_ _13971_/C _13971_/B _13971_/A _13971_/D vssd1 vssd1 vccd1 vccd1 _13967_/X
+ sky130_fd_sc_hd__and4b_4
XFILLER_62_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12918_ _12918_/A _12949_/Y vssd1 vssd1 vccd1 vccd1 _13758_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_80_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13898_ _13905_/A _13905_/B _13905_/C _13905_/D vssd1 vssd1 vccd1 vccd1 _13898_/Y
+ sky130_fd_sc_hd__nor4b_4
XANTENNA__10909__D line[38] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12396__D line[92] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12849_ _12875_/CLK line[43] vssd1 vssd1 vccd1 vccd1 _12850_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_22_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_OVHB\[30\].CG_CLK clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06394__D line[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06370_ _06400_/CLK line[16] vssd1 vssd1 vccd1 vccd1 _06371_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_202_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05321_ _05321_/A _05354_/Y vssd1 vssd1 vccd1 vccd1 _13721_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[29\].CLKBUF\[5\] clk vssd1 vssd1 vccd1 vccd1 _11022_/CLK sky130_fd_sc_hd__clkbuf_4
X_08040_ _08040_/A _08049_/Y vssd1 vssd1 vccd1 vccd1 _13640_/Z sky130_fd_sc_hd__ebufn_2
X_05252_ _05280_/CLK line[26] vssd1 vssd1 vccd1 vccd1 _05253_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__04916__A1_N A_h[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10644__D line[59] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05183_ _05183_/A _05214_/Y vssd1 vssd1 vccd1 vccd1 _13863_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13020__D line[112] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09991_ _10005_/CLK line[2] vssd1 vssd1 vccd1 vccd1 _09992_/A sky130_fd_sc_hd__dfxtp_1
X_08942_ _08942_/A _08959_/Y vssd1 vssd1 vccd1 vccd1 _13702_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12214__A _13934_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[9\].VALID\[3\].FF_D A[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07953__D line[109] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08873_ _08885_/CLK line[3] vssd1 vssd1 vccd1 vccd1 _08874_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_29_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11475__D line[41] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07824_ _07824_/A _07839_/Y vssd1 vssd1 vccd1 vccd1 _13704_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06569__D line[102] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_04967_ _04967_/CLK _04968_/X vssd1 vssd1 vccd1 vccd1 _04965_/CLK sky130_fd_sc_hd__dlclkp_1
X_07755_ _07765_/CLK line[4] vssd1 vssd1 vccd1 vccd1 _07756_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_25_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06706_ _06706_/A _06719_/Y vssd1 vssd1 vccd1 vccd1 _13706_/Z sky130_fd_sc_hd__ebufn_2
X_07686_ _07686_/A _07699_/Y vssd1 vssd1 vccd1 vccd1 _13846_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09425_ _09445_/CLK line[14] vssd1 vssd1 vccd1 vccd1 _09426_/A sky130_fd_sc_hd__dfxtp_1
X_06637_ _06645_/CLK line[5] vssd1 vssd1 vccd1 vccd1 _06638_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_197_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10819__D line[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07978__A _13912_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09356_ _09356_/A _09379_/Y vssd1 vssd1 vccd1 vccd1 _13836_/Z sky130_fd_sc_hd__ebufn_2
X_06568_ _06568_/A _06579_/Y vssd1 vssd1 vccd1 vccd1 _13848_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_60_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08307_ _08325_/CLK line[15] vssd1 vssd1 vccd1 vccd1 _08308_/A sky130_fd_sc_hd__dfxtp_1
X_05519_ _05525_/CLK line[6] vssd1 vssd1 vccd1 vccd1 _05520_/A sky130_fd_sc_hd__dfxtp_1
X_09287_ _09305_/CLK line[79] vssd1 vssd1 vccd1 vccd1 _09288_/A sky130_fd_sc_hd__dfxtp_1
X_06499_ _06505_/CLK line[70] vssd1 vssd1 vccd1 vccd1 _06500_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_165_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08238_ _08238_/A _08259_/Y vssd1 vssd1 vccd1 vccd1 _13838_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_176_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12108__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08169_ _08185_/CLK line[65] vssd1 vssd1 vccd1 vccd1 _08170_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[9\].VALID\[6\].FF OVHB\[9\].V/CLK A[13] vssd1 vssd1 vccd1 vccd1 OVHB\[9\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_118_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10200_ _10200_/A _10219_/Y vssd1 vssd1 vccd1 vccd1 _13840_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[28\].CLKBUF\[2\] clk vssd1 vssd1 vccd1 vccd1 _10637_/CLK sky130_fd_sc_hd__clkbuf_4
X_11180_ _11180_/A _11199_/Y vssd1 vssd1 vccd1 vccd1 _13700_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_192_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10131_ _10145_/CLK line[66] vssd1 vssd1 vccd1 vccd1 _10132_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_88_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10062_ _10062_/A _10079_/Y vssd1 vssd1 vccd1 vccd1 _13702_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[1\].VALID\[7\].TOBUF OVHB\[1\].VALID\[7\].FF/Q OVHB\[1\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/A2 sky130_fd_sc_hd__ebufn_2
XANTENNA__11385__D line[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06479__D line[75] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05383__D line[72] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13821_ _13821_/A _13824_/Y vssd1 vssd1 vccd1 vccd1 _13821_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_28_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08694__D line[49] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13752_ _13752_/CLK _13753_/X vssd1 vssd1 vccd1 vccd1 _13750_/CLK sky130_fd_sc_hd__dlclkp_1
X_10964_ _10964_/A _10989_/Y vssd1 vssd1 vccd1 vccd1 _13764_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08049__A _13932_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12703_ _13936_/X wr vssd1 vssd1 vccd1 vccd1 _12703_/X sky130_fd_sc_hd__and2_1
XFILLER_204_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13683_ _13899_/X wr vssd1 vssd1 vccd1 vccd1 _13683_/X sky130_fd_sc_hd__and2_1
X_10895_ _10915_/CLK line[46] vssd1 vssd1 vccd1 vccd1 _10896_/A sky130_fd_sc_hd__dfxtp_1
XPHY_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12634_ _13936_/X vssd1 vssd1 vccd1 vccd1 _12634_/Y sky130_fd_sc_hd__inv_2
XPHY_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_DATA\[23\].CLKBUF\[3\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12565_ _12595_/CLK line[32] vssd1 vssd1 vccd1 vccd1 _12566_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06942__D line[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11516_ _11516_/A _11549_/Y vssd1 vssd1 vccd1 vccd1 _13756_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12496_ _12496_/A _12529_/Y vssd1 vssd1 vccd1 vccd1 _13616_/Z sky130_fd_sc_hd__ebufn_2
X_11447_ _11475_/CLK line[42] vssd1 vssd1 vccd1 vccd1 _11448_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05558__D line[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11378_ _11378_/A _11409_/Y vssd1 vssd1 vccd1 vccd1 _13618_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13775__D line[68] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13117_ _13117_/A _13124_/Y vssd1 vssd1 vccd1 vccd1 _13677_/Z sky130_fd_sc_hd__ebufn_2
X_10329_ _10355_/CLK line[43] vssd1 vssd1 vccd1 vccd1 _10330_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_152_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08869__D line[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13048_ _13050_/CLK line[120] vssd1 vssd1 vccd1 vccd1 _13049_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[7\].VALID\[8\].FF OVHB\[7\].V/CLK A[15] vssd1 vssd1 vccd1 vccd1 OVHB\[7\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XMUX.M\[3\].MUX\[0\] _13679_/Z _13749_/Z _13819_/Z _13889_/Z MUX.SEL0BUF\[3\]/X MUX.SEL1BUF\[3\]/X
+ vssd1 vssd1 vccd1 vccd1 Do[24] sky130_fd_sc_hd__mux4_1
XFILLER_39_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05870_ _05870_/A _05879_/Y vssd1 vssd1 vccd1 vccd1 _13710_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05293__D line[45] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09343__A _13916_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDATA\[17\].CLKBUF\[5\] clk vssd1 vssd1 vccd1 vccd1 _07382_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_94_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07540_ _07540_/A _07559_/Y vssd1 vssd1 vccd1 vccd1 _13700_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_207_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07471_ _07485_/CLK line[2] vssd1 vssd1 vccd1 vccd1 _07472_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13015__D line[105] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06422_ _06422_/A _06439_/Y vssd1 vssd1 vccd1 vccd1 _13702_/Z sky130_fd_sc_hd__ebufn_2
X_09210_ _09210_/A _09239_/Y vssd1 vssd1 vccd1 vccd1 _13690_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08109__D line[38] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09141_ _09165_/CLK line[12] vssd1 vssd1 vccd1 vccd1 _09142_/A sky130_fd_sc_hd__dfxtp_1
X_06353_ _06365_/CLK line[3] vssd1 vssd1 vccd1 vccd1 _06354_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[7\].V OVHB\[7\].V/CLK TIE/HI rst_n vssd1 vssd1 vccd1 vccd1 OVHB\[7\].V/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_187_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05304_ _05304_/A _05319_/Y vssd1 vssd1 vccd1 vccd1 _13704_/Z sky130_fd_sc_hd__ebufn_2
X_09072_ _09072_/A _09099_/Y vssd1 vssd1 vccd1 vccd1 _13832_/Z sky130_fd_sc_hd__ebufn_2
X_06284_ _06284_/A _06299_/Y vssd1 vssd1 vccd1 vccd1 _13844_/Z sky130_fd_sc_hd__ebufn_2
X_08023_ _08045_/CLK line[13] vssd1 vssd1 vccd1 vccd1 _08024_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_190_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05235_ _05245_/CLK line[4] vssd1 vssd1 vccd1 vccd1 _05236_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10374__D line[49] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[7\].VALID\[13\].TOBUF OVHB\[7\].VALID\[13\].FF/Q OVHB\[7\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04916_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__05468__D line[125] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09518__A _13920_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05166_ _05166_/A _05179_/Y vssd1 vssd1 vccd1 vccd1 _13846_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_89_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13685__D line[32] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09974_ _13921_/X vssd1 vssd1 vccd1 vccd1 _09974_/Y sky130_fd_sc_hd__inv_2
X_05097_ _05105_/CLK line[69] vssd1 vssd1 vccd1 vccd1 _05098_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_39_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07683__D line[99] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08925_ _08955_/CLK line[32] vssd1 vssd1 vccd1 vccd1 _08926_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12879__A _13937_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08856_ _08856_/A _08889_/Y vssd1 vssd1 vccd1 vccd1 _13616_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[30\].V OVHB\[30\].V/CLK TIE/HI rst_n vssd1 vssd1 vccd1 vccd1 OVHB\[30\].V/Q
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_OVHB\[31\].VALID\[7\].FF_D A[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12598__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07807_ _07835_/CLK line[42] vssd1 vssd1 vccd1 vccd1 _07808_/A sky130_fd_sc_hd__dfxtp_1
X_05999_ _06015_/CLK line[97] vssd1 vssd1 vccd1 vccd1 _06000_/A sky130_fd_sc_hd__dfxtp_1
X_08787_ _08815_/CLK line[106] vssd1 vssd1 vccd1 vccd1 _08788_/A sky130_fd_sc_hd__dfxtp_1
X_07738_ _07738_/A _07769_/Y vssd1 vssd1 vccd1 vccd1 _13618_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__04932__B2 _04932_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05931__D line[66] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10549__D line[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDATA\[16\].CLKBUF\[2\] clk vssd1 vssd1 vccd1 vccd1 _06997_/CLK sky130_fd_sc_hd__clkbuf_4
X_07669_ _07695_/CLK line[107] vssd1 vssd1 vccd1 vccd1 _07670_/A sky130_fd_sc_hd__dfxtp_1
X_09408_ _09410_/CLK line[120] vssd1 vssd1 vccd1 vccd1 _09409_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[0\].VALID\[12\].TOBUF OVHB\[0\].VALID\[12\].FF/Q OVHB\[0\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04929_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__08019__D line[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10680_ _10680_/A _10709_/Y vssd1 vssd1 vccd1 vccd1 _13760_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_71_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XMUX.M\[2\].MUX\[2\] _13667_/Z _13737_/Z _13807_/Z _13877_/Z MUX.SEL0BUF\[2\]/X MUX.SEL1BUF\[2\]/X
+ vssd1 vssd1 vccd1 vccd1 Do[18] sky130_fd_sc_hd__mux4_1
X_09339_ _09339_/A _09344_/Y vssd1 vssd1 vccd1 vccd1 _13819_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12764__D line[118] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07858__D line[51] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11023__A _13925_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12350_ _12350_/CLK line[57] vssd1 vssd1 vccd1 vccd1 _12351_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_138_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11301_ _11301_/A _11304_/Y vssd1 vssd1 vccd1 vccd1 _13821_/Z sky130_fd_sc_hd__ebufn_2
X_12281_ _12281_/A _12284_/Y vssd1 vssd1 vccd1 vccd1 _13681_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_119_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11232_ _11232_/CLK _11233_/X vssd1 vssd1 vccd1 vccd1 _11230_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_153_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[23\].VALID\[13\].FF OVHB\[23\].V/CLK A[20] vssd1 vssd1 vccd1 vccd1 OVHB\[23\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_11163_ _13933_/X wr vssd1 vssd1 vccd1 vccd1 _11163_/X sky130_fd_sc_hd__and2_1
XFILLER_122_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10114_ _13922_/X vssd1 vssd1 vccd1 vccd1 _10114_/Y sky130_fd_sc_hd__inv_2
XFILLER_122_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11094_ _13925_/X vssd1 vssd1 vccd1 vccd1 _11094_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10045_ _10075_/CLK line[32] vssd1 vssd1 vccd1 vccd1 _10046_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_75_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XOVHB\[21\].V OVHB\[21\].V/CLK TIE/HI rst_n vssd1 vssd1 vccd1 vccd1 OVHB\[21\].V/Q
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_48_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XOVHB\[16\].VALID\[0\].FF OVHB\[16\].V/CLK A[7] vssd1 vssd1 vccd1 vccd1 OVHB\[16\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__12939__D line[70] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13804_ _13820_/CLK line[81] vssd1 vssd1 vccd1 vccd1 _13805_/A sky130_fd_sc_hd__dfxtp_1
X_11996_ _12000_/CLK line[23] vssd1 vssd1 vccd1 vccd1 _11997_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_45_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13735_ _13735_/A _13754_/Y vssd1 vssd1 vccd1 vccd1 _13735_/Z sky130_fd_sc_hd__ebufn_2
X_10947_ _10947_/A _10954_/Y vssd1 vssd1 vccd1 vccd1 _13747_/Z sky130_fd_sc_hd__ebufn_2
X_13666_ _13680_/CLK line[18] vssd1 vssd1 vccd1 vccd1 _13667_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[22\].VALID\[14\].FF_D A[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10878_ _10880_/CLK line[24] vssd1 vssd1 vccd1 vccd1 _10879_/A sky130_fd_sc_hd__dfxtp_1
XPHY_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12674__D line[91] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12617_ _12617_/A _12634_/Y vssd1 vssd1 vccd1 vccd1 _13737_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[22\].V_D TIE/HI vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13597_ _13597_/A _13614_/Y vssd1 vssd1 vccd1 vccd1 _13877_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_8_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06672__D line[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12548_ _12560_/CLK line[19] vssd1 vssd1 vccd1 vccd1 _12549_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_157_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12479_ _12479_/A _12494_/Y vssd1 vssd1 vccd1 vccd1 _13879_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09983__D line[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05020_ _05020_/A _05039_/Y vssd1 vssd1 vccd1 vccd1 _13700_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[5\].VALID\[6\].FF_D A[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[21\].CLKBUF\[5\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10922__D line[58] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08599__D line[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06971_ _06995_/CLK line[44] vssd1 vssd1 vccd1 vccd1 _06972_/A sky130_fd_sc_hd__dfxtp_1
XMUX.M\[1\].MUX\[4\] _13622_/Z _13692_/Z _13762_/Z _13832_/Z MUX.SEL0BUF\[1\]/X MUX.SEL1BUF\[1\]/X
+ vssd1 vssd1 vccd1 vccd1 Do[12] sky130_fd_sc_hd__mux4_1
XFILLER_140_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_MUX.M\[2\].MUX\[0\]_A1 _13721_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08710_ _08710_/CLK line[57] vssd1 vssd1 vccd1 vccd1 _08711_/A sky130_fd_sc_hd__dfxtp_1
X_05922_ _05922_/A _05949_/Y vssd1 vssd1 vccd1 vccd1 _13762_/Z sky130_fd_sc_hd__ebufn_2
X_09690_ _09690_/CLK line[121] vssd1 vssd1 vccd1 vccd1 _09691_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[12\].V OVHB\[12\].V/CLK TIE/HI rst_n vssd1 vssd1 vccd1 vccd1 OVHB\[12\].V/Q
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07008__D line[61] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08641_ _08641_/A _08644_/Y vssd1 vssd1 vccd1 vccd1 _13681_/Z sky130_fd_sc_hd__ebufn_2
X_05853_ _05875_/CLK line[45] vssd1 vssd1 vccd1 vccd1 _05854_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12849__D line[43] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11753__D line[40] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[8\].VALID\[7\].TOBUF OVHB\[8\].VALID\[7\].FF/Q OVHB\[8\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/A2 sky130_fd_sc_hd__ebufn_2
XANTENNA__06847__D line[101] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05784_ _05784_/A _05809_/Y vssd1 vssd1 vccd1 vccd1 _13624_/Z sky130_fd_sc_hd__ebufn_2
X_08572_ _08572_/CLK _08573_/X vssd1 vssd1 vccd1 vccd1 _08570_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__04914__B2 _04914_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09223__D line[35] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07523_ _13911_/X wr vssd1 vssd1 vccd1 vccd1 _07523_/X sky130_fd_sc_hd__and2_1
XFILLER_179_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07454_ _13910_/X vssd1 vssd1 vccd1 vccd1 _07454_/Y sky130_fd_sc_hd__inv_2
XPHY_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[14\].VALID\[2\].FF OVHB\[14\].V/CLK A[9] vssd1 vssd1 vccd1 vccd1 OVHB\[14\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_195_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06405_ _06435_/CLK line[32] vssd1 vssd1 vccd1 vccd1 _06406_/A sky130_fd_sc_hd__dfxtp_1
X_07385_ _07415_/CLK line[96] vssd1 vssd1 vccd1 vccd1 _07386_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_176_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_OVHB\[14\].VALID\[11\].FF_D A[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[31\].VALID\[6\].FF OVHB\[31\].V/CLK A[13] vssd1 vssd1 vccd1 vccd1 OVHB\[31\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_41_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06336_ _06336_/A _06369_/Y vssd1 vssd1 vccd1 vccd1 _13616_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06582__D line[122] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09124_ _09130_/CLK line[118] vssd1 vssd1 vccd1 vccd1 _09125_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[23\].VALID\[14\].TOBUF OVHB\[23\].VALID\[14\].FF/Q OVHB\[23\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_163_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09055_ _09055_/A _09064_/Y vssd1 vssd1 vccd1 vccd1 _13815_/Z sky130_fd_sc_hd__ebufn_2
X_06267_ _06295_/CLK line[106] vssd1 vssd1 vccd1 vccd1 _06268_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05198__D line[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05218_ _05218_/A _05249_/Y vssd1 vssd1 vccd1 vccd1 _13618_/Z sky130_fd_sc_hd__ebufn_2
X_08006_ _08010_/CLK line[119] vssd1 vssd1 vccd1 vccd1 _08007_/A sky130_fd_sc_hd__dfxtp_1
X_06198_ _06198_/A _06229_/Y vssd1 vssd1 vccd1 vccd1 _13758_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_163_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11928__D line[120] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05149_ _05175_/CLK line[107] vssd1 vssd1 vccd1 vccd1 _05150_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_150_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09957_ _09957_/A _09974_/Y vssd1 vssd1 vccd1 vccd1 _13877_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_106_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[24\].VALID\[10\].FF_D A[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08908_ _08920_/CLK line[19] vssd1 vssd1 vccd1 vccd1 _08909_/A sky130_fd_sc_hd__dfxtp_1
X_09888_ _09900_/CLK line[83] vssd1 vssd1 vccd1 vccd1 _09889_/A sky130_fd_sc_hd__dfxtp_1
X_08839_ _08839_/A _08854_/Y vssd1 vssd1 vccd1 vccd1 _13879_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_17_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11663__D line[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11850_ _11860_/CLK line[84] vssd1 vssd1 vccd1 vccd1 _11851_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_17_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06757__D line[74] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05661__D line[71] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10801_ _10801_/A _10814_/Y vssd1 vssd1 vccd1 vccd1 _13881_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10279__D line[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11781_ _11781_/A _11794_/Y vssd1 vssd1 vccd1 vccd1 _13741_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_159_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13520_ _13540_/CLK line[94] vssd1 vssd1 vccd1 vccd1 _13521_/A sky130_fd_sc_hd__dfxtp_1
X_10732_ _10740_/CLK line[85] vssd1 vssd1 vccd1 vccd1 _10733_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08972__D line[63] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XMUX.M\[0\].MUX\[6\] _13640_/Z _13710_/Z _13780_/Z _13850_/Z MUX.SEL0BUF\[0\]/X MUX.SEL1BUF\[0\]/X
+ vssd1 vssd1 vccd1 vccd1 Do[6] sky130_fd_sc_hd__mux4_1
X_13451_ _13451_/A _13474_/Y vssd1 vssd1 vccd1 vccd1 _13731_/Z sky130_fd_sc_hd__ebufn_2
X_10663_ _10663_/A _10674_/Y vssd1 vssd1 vccd1 vccd1 _13743_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_139_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07588__D line[56] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[15\].VALID\[2\].TOBUF OVHB\[15\].VALID\[2\].FF/Q OVHB\[15\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04930_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_139_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12402_ _12420_/CLK line[95] vssd1 vssd1 vccd1 vccd1 _12403_/A sky130_fd_sc_hd__dfxtp_1
X_10594_ _10600_/CLK line[22] vssd1 vssd1 vccd1 vccd1 _10595_/A sky130_fd_sc_hd__dfxtp_1
X_13382_ _13400_/CLK line[31] vssd1 vssd1 vccd1 vccd1 _13383_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11688__A _13927_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12333_ _12333_/A _12354_/Y vssd1 vssd1 vccd1 vccd1 _13733_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_31_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XOVHB\[12\].VALID\[4\].FF OVHB\[12\].V/CLK A[11] vssd1 vssd1 vccd1 vccd1 OVHB\[12\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_5_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12264_ _12280_/CLK line[17] vssd1 vssd1 vccd1 vccd1 _12265_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11838__D line[93] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11215_ _11215_/A _11234_/Y vssd1 vssd1 vccd1 vccd1 _13735_/Z sky130_fd_sc_hd__ebufn_2
X_12195_ _12195_/A _12214_/Y vssd1 vssd1 vccd1 vccd1 _13875_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_150_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05836__D line[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08212__D line[85] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11146_ _11160_/CLK line[18] vssd1 vssd1 vccd1 vccd1 _11147_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_122_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11077_ _11077_/A _11094_/Y vssd1 vssd1 vccd1 vccd1 _13877_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[7\].V_D TIE/HI vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10028_ _10040_/CLK line[19] vssd1 vssd1 vccd1 vccd1 _10029_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_64_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05571__D line[44] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10189__D line[107] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11979_ _11979_/A _12004_/Y vssd1 vssd1 vccd1 vccd1 _13659_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_44_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13718_ _13899_/X wr vssd1 vssd1 vccd1 vccd1 _13718_/X sky130_fd_sc_hd__and2_1
XFILLER_177_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13649_ _13899_/X vssd1 vssd1 vccd1 vccd1 _13649_/Y sky130_fd_sc_hd__inv_2
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07498__D line[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07170_ _07170_/CLK line[121] vssd1 vssd1 vccd1 vccd1 _07171_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_118_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06121_ _06121_/A _06124_/Y vssd1 vssd1 vccd1 vccd1 _13681_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_172_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06052_ _06052_/CLK _06053_/X vssd1 vssd1 vccd1 vccd1 _06050_/CLK sky130_fd_sc_hd__dlclkp_1
XOVHB\[28\].VALID\[9\].FF OVHB\[28\].V/CLK A[16] vssd1 vssd1 vccd1 vccd1 OVHB\[28\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_05003_ _13931_/Y wr vssd1 vssd1 vccd1 vccd1 _05003_/X sky130_fd_sc_hd__and2_1
XANTENNA__10652__D line[63] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_OVHB\[4\].CG_CLK clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05746__D line[124] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09811_ _09811_/A _09834_/Y vssd1 vssd1 vccd1 vccd1 _13731_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[21\].VALID\[1\].TOBUF OVHB\[21\].VALID\[1\].FF/Q OVHB\[21\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04926_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__08122__D line[58] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09742_ _09760_/CLK line[31] vssd1 vssd1 vccd1 vccd1 _09743_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_86_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06954_ _06960_/CLK line[22] vssd1 vssd1 vccd1 vccd1 _06955_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_101_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[10\].VALID\[6\].FF OVHB\[10\].V/CLK A[13] vssd1 vssd1 vccd1 vccd1 OVHB\[10\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__07961__D line[98] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05905_ _05905_/A _05914_/Y vssd1 vssd1 vccd1 vccd1 _13745_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12579__D line[33] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09673_ _09673_/A _09694_/Y vssd1 vssd1 vccd1 vccd1 _13873_/Z sky130_fd_sc_hd__ebufn_2
X_06885_ _06885_/A _06894_/Y vssd1 vssd1 vccd1 vccd1 _13885_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_39_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08624_ _08640_/CLK line[17] vssd1 vssd1 vccd1 vccd1 _08625_/A sky130_fd_sc_hd__dfxtp_1
X_05836_ _05840_/CLK line[23] vssd1 vssd1 vccd1 vccd1 _05837_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_54_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XOVHB\[11\].INV _13945_/X vssd1 vssd1 vccd1 vccd1 OVHB\[11\].INV/Y sky130_fd_sc_hd__inv_2
XPHY_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08555_ _08555_/A _08574_/Y vssd1 vssd1 vccd1 vccd1 _13875_/Z sky130_fd_sc_hd__ebufn_2
X_05767_ _05767_/A _05774_/Y vssd1 vssd1 vccd1 vccd1 _13887_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09888__D line[83] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13053__A _13937_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07506_ _07520_/CLK line[18] vssd1 vssd1 vccd1 vccd1 _07507_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08486_ _08500_/CLK line[82] vssd1 vssd1 vccd1 vccd1 _08487_/A sky130_fd_sc_hd__dfxtp_1
X_05698_ _05700_/CLK line[88] vssd1 vssd1 vccd1 vccd1 _05699_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10827__D line[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07437_ _07437_/A _07454_/Y vssd1 vssd1 vccd1 vccd1 _13877_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_50_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XOVHB\[26\].INV _13966_/X vssd1 vssd1 vccd1 vccd1 OVHB\[26\].INV/Y sky130_fd_sc_hd__inv_2
XPHY_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13203__D line[77] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_OVHB\[29\].VALID\[14\].FF_D A[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07368_ _07380_/CLK line[83] vssd1 vssd1 vccd1 vccd1 _07369_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07201__D line[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09107_ _09107_/A _09134_/Y vssd1 vssd1 vccd1 vccd1 _13867_/Z sky130_fd_sc_hd__ebufn_2
X_06319_ _06319_/A _06334_/Y vssd1 vssd1 vccd1 vccd1 _13879_/Z sky130_fd_sc_hd__ebufn_2
X_07299_ _07299_/A _07314_/Y vssd1 vssd1 vccd1 vccd1 _13739_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_163_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09038_ _09060_/CLK line[93] vssd1 vssd1 vccd1 vccd1 _09039_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[10\].VALID\[2\].FF_D A[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09128__D line[120] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11000_ _11020_/CLK line[94] vssd1 vssd1 vccd1 vccd1 _11001_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_132_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13228__A _13938_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[13\].VALID\[7\].TOBUF OVHB\[13\].VALID\[7\].FF/Q OVHB\[13\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/A2 sky130_fd_sc_hd__ebufn_2
X_12951_ _12951_/A _12984_/Y vssd1 vssd1 vccd1 vccd1 _13791_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11393__D line[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11902_ _11930_/CLK line[122] vssd1 vssd1 vccd1 vccd1 _11903_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06487__D line[79] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12882_ _12910_/CLK line[58] vssd1 vssd1 vccd1 vccd1 _12883_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[7\].CLKBUF\[6\] clk vssd1 vssd1 vccd1 vccd1 _13297_/CLK sky130_fd_sc_hd__clkbuf_4
X_11833_ _11833_/A _11864_/Y vssd1 vssd1 vccd1 vccd1 _13793_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_61_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11764_ _11790_/CLK line[59] vssd1 vssd1 vccd1 vccd1 _11765_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_202_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13503_ _13505_/CLK line[72] vssd1 vssd1 vccd1 vccd1 _13504_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10715_ _10715_/A _10744_/Y vssd1 vssd1 vccd1 vccd1 _13795_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11695_ _11695_/A _11724_/Y vssd1 vssd1 vccd1 vccd1 _13655_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13434_ _13434_/A _13439_/Y vssd1 vssd1 vccd1 vccd1 _13714_/Z sky130_fd_sc_hd__ebufn_2
X_10646_ _10670_/CLK line[60] vssd1 vssd1 vccd1 vccd1 _10647_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07111__D line[108] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[26\].CGAND_B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12952__D line[90] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[1\].VALID\[9\].FF_D A[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13365_ _13365_/CLK line[9] vssd1 vssd1 vccd1 vccd1 _13366_/A sky130_fd_sc_hd__dfxtp_1
X_10577_ _10577_/A _10604_/Y vssd1 vssd1 vccd1 vccd1 _13657_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06950__D line[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12316_ _12316_/A _12319_/Y vssd1 vssd1 vccd1 vccd1 _13716_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_181_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13296_ _13296_/A _13299_/Y vssd1 vssd1 vccd1 vccd1 _13856_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11568__D line[83] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12247_ _12247_/CLK _12248_/X vssd1 vssd1 vccd1 vccd1 _12245_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__09038__D line[93] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12178_ _13934_/X wr vssd1 vssd1 vccd1 vccd1 _12178_/X sky130_fd_sc_hd__and2_1
XANTENNA__13783__D line[72] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11129_ _13933_/X vssd1 vssd1 vccd1 vccd1 _11129_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08877__D line[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06670_ _06680_/CLK line[20] vssd1 vssd1 vccd1 vccd1 _06671_/A sky130_fd_sc_hd__dfxtp_1
X_05621_ _05621_/A _05634_/Y vssd1 vssd1 vccd1 vccd1 _13741_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_24_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05552_ _05560_/CLK line[21] vssd1 vssd1 vccd1 vccd1 _05553_/A sky130_fd_sc_hd__dfxtp_1
X_08340_ _08360_/CLK line[30] vssd1 vssd1 vccd1 vccd1 _08341_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_205_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09501__D line[34] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDATA\[6\].CLKBUF\[3\] clk vssd1 vssd1 vccd1 vccd1 _12912_/CLK sky130_fd_sc_hd__clkbuf_4
X_08271_ _08271_/A _08294_/Y vssd1 vssd1 vccd1 vccd1 _13871_/Z sky130_fd_sc_hd__ebufn_2
X_05483_ _05483_/A _05494_/Y vssd1 vssd1 vccd1 vccd1 _13883_/Z sky130_fd_sc_hd__ebufn_2
X_07222_ _07240_/CLK line[31] vssd1 vssd1 vccd1 vccd1 _07223_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_146_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07153_ _07153_/A _07174_/Y vssd1 vssd1 vccd1 vccd1 _13873_/Z sky130_fd_sc_hd__ebufn_2
X_06104_ _06120_/CLK line[17] vssd1 vssd1 vccd1 vccd1 _06105_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06860__D line[112] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[23\].VALID\[2\].FF_D A[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07084_ _07100_/CLK line[81] vssd1 vssd1 vccd1 vccd1 _07085_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10382__D line[53] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06035_ _06035_/A _06054_/Y vssd1 vssd1 vccd1 vccd1 _13875_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05476__D line[114] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13693__D line[45] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05773__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[16\].VALID\[6\].FF_D A[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08787__D line[106] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07691__D line[103] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07986_ _08010_/CLK line[124] vssd1 vssd1 vccd1 vccd1 _07987_/A sky130_fd_sc_hd__dfxtp_1
X_09725_ _09725_/CLK line[9] vssd1 vssd1 vccd1 vccd1 _09726_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_86_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06937_ _06937_/A _06964_/Y vssd1 vssd1 vccd1 vccd1 _13657_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_170_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09656_ _09656_/A _09659_/Y vssd1 vssd1 vccd1 vccd1 _13856_/Z sky130_fd_sc_hd__ebufn_2
X_06868_ _06890_/CLK line[125] vssd1 vssd1 vccd1 vccd1 _06869_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[26\].CLKBUF\[7\] clk vssd1 vssd1 vccd1 vccd1 _10252_/CLK sky130_fd_sc_hd__clkbuf_4
X_08607_ _08607_/CLK _08608_/X vssd1 vssd1 vccd1 vccd1 _08605_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__06100__D line[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05819_ _05819_/A _05844_/Y vssd1 vssd1 vccd1 vccd1 _13659_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_43_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09587_ _09587_/CLK _09588_/X vssd1 vssd1 vccd1 vccd1 _09585_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA__11941__D line[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06799_ _06799_/A _06824_/Y vssd1 vssd1 vccd1 vccd1 _13799_/Z sky130_fd_sc_hd__ebufn_2
XPHY_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08538_ _13913_/X wr vssd1 vssd1 vccd1 vccd1 _08538_/X sky130_fd_sc_hd__and2_1
XPHY_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10557__D line[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08469_ _13913_/X vssd1 vssd1 vccd1 vccd1 _08469_/Y sky130_fd_sc_hd__inv_2
XPHY_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[13\].VALID\[12\].TOBUF OVHB\[13\].VALID\[12\].FF/Q OVHB\[13\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04929_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_10_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10500_ _10530_/CLK line[112] vssd1 vssd1 vccd1 vccd1 _10501_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08027__D line[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[28\].VALID\[13\].FF OVHB\[28\].V/CLK A[20] vssd1 vssd1 vccd1 vccd1 OVHB\[28\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_11480_ _11510_/CLK line[48] vssd1 vssd1 vccd1 vccd1 _11481_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13868__D line[125] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10431_ _10431_/A _10464_/Y vssd1 vssd1 vccd1 vccd1 _13791_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_195_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05948__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDATA\[5\].CLKBUF\[0\] clk vssd1 vssd1 vccd1 vccd1 _12527_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__07866__D line[55] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13150_ _13150_/A _13159_/Y vssd1 vssd1 vccd1 vccd1 _13710_/Z sky130_fd_sc_hd__ebufn_2
X_10362_ _10390_/CLK line[58] vssd1 vssd1 vccd1 vccd1 _10363_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_163_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10292__D line[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12101_ _12105_/CLK line[71] vssd1 vssd1 vccd1 vccd1 _12102_/A sky130_fd_sc_hd__dfxtp_1
X_13081_ _13085_/CLK line[7] vssd1 vssd1 vccd1 vccd1 _13082_/A sky130_fd_sc_hd__dfxtp_1
X_10293_ _10293_/A _10324_/Y vssd1 vssd1 vccd1 vccd1 _13653_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_105_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12032_ _12032_/A _12039_/Y vssd1 vssd1 vccd1 vccd1 _13712_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_77_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XOVHB\[28\].VALID\[1\].TOBUF OVHB\[28\].VALID\[1\].FF/Q OVHB\[28\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04926_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_77_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13108__D line[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12934_ _12934_/A _12949_/Y vssd1 vssd1 vccd1 vccd1 _13774_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_37_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12865_ _12875_/CLK line[36] vssd1 vssd1 vccd1 vccd1 _12866_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[23\].VOBUF OVHB\[23\].V/Q OVHB\[23\].INV/Y vssd1 vssd1 vccd1 vccd1 _04912_/B1
+ sky130_fd_sc_hd__ebufn_2
X_11816_ _11816_/A _11829_/Y vssd1 vssd1 vccd1 vccd1 _13776_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_61_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12796_ _12796_/A _12809_/Y vssd1 vssd1 vccd1 vccd1 _13636_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XDATA\[25\].CLKBUF\[4\] clk vssd1 vssd1 vccd1 vccd1 _09867_/CLK sky130_fd_sc_hd__clkbuf_4
XOVHB\[1\].VALID\[1\].FF OVHB\[1\].V/CLK A[8] vssd1 vssd1 vccd1 vccd1 OVHB\[1\].VALID\[1\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10467__D line[106] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11747_ _11755_/CLK line[37] vssd1 vssd1 vccd1 vccd1 _11748_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_159_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11678_ _11678_/A _11689_/Y vssd1 vssd1 vccd1 vccd1 _13638_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12682__D line[95] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13417_ _13435_/CLK line[47] vssd1 vssd1 vccd1 vccd1 _13418_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_146_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10629_ _10635_/CLK line[38] vssd1 vssd1 vccd1 vccd1 _10630_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_127_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07776__D line[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06680__D line[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13348_ _13348_/A _13369_/Y vssd1 vssd1 vccd1 vccd1 _13628_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.M\[3\].MUX\[2\]_A1 _13723_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11298__D line[88] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13279_ _13295_/CLK line[97] vssd1 vssd1 vccd1 vccd1 _13280_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09991__D line[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[29\].VALID\[6\].FF_D A[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10930__D line[62] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07840_ _07870_/CLK line[48] vssd1 vssd1 vccd1 vccd1 _07841_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_110_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08400__D line[48] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07771_ _07771_/A _07804_/Y vssd1 vssd1 vccd1 vccd1 _13651_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_83_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_04983_ _04983_/A _05004_/Y vssd1 vssd1 vccd1 vccd1 _13663_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_84_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09510_ _09510_/A _09519_/Y vssd1 vssd1 vccd1 vccd1 _13710_/Z sky130_fd_sc_hd__ebufn_2
X_06722_ _06750_/CLK line[58] vssd1 vssd1 vccd1 vccd1 _06723_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07016__D line[50] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09441_ _09445_/CLK line[7] vssd1 vssd1 vccd1 vccd1 _09442_/A sky130_fd_sc_hd__dfxtp_1
X_06653_ _06653_/A _06684_/Y vssd1 vssd1 vccd1 vccd1 _13653_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12857__D line[47] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05604_ _05630_/CLK line[59] vssd1 vssd1 vccd1 vccd1 _05605_/A sky130_fd_sc_hd__dfxtp_1
X_09372_ _09372_/A _09379_/Y vssd1 vssd1 vccd1 vccd1 _13852_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07313__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06855__D line[105] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06584_ _06610_/CLK line[123] vssd1 vssd1 vccd1 vccd1 _06585_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09231__D line[39] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08323_ _08325_/CLK line[8] vssd1 vssd1 vccd1 vccd1 _08324_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_33_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_DATA\[12\].CLKBUF\[1\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05535_ _05535_/A _05564_/Y vssd1 vssd1 vccd1 vccd1 _13655_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_32_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05466_ _05490_/CLK line[124] vssd1 vssd1 vccd1 vccd1 _05467_/A sky130_fd_sc_hd__dfxtp_1
X_08254_ _08254_/A _08259_/Y vssd1 vssd1 vccd1 vccd1 _13854_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_192_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07205_ _07205_/CLK line[9] vssd1 vssd1 vccd1 vccd1 _07206_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_165_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XDATA\[24\].CLKBUF\[1\] clk vssd1 vssd1 vccd1 vccd1 _09482_/CLK sky130_fd_sc_hd__clkbuf_4
X_08185_ _08185_/CLK line[73] vssd1 vssd1 vccd1 vccd1 _08186_/A sky130_fd_sc_hd__dfxtp_1
X_05397_ _05397_/A _05424_/Y vssd1 vssd1 vccd1 vccd1 _13797_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06590__D line[126] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07136_ _07136_/A _07139_/Y vssd1 vssd1 vccd1 vccd1 _13856_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[14\].CLKBUF\[7\] clk vssd1 vssd1 vccd1 vccd1 _06612_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_161_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07067_ _07067_/CLK _07068_/X vssd1 vssd1 vccd1 vccd1 _07065_/CLK sky130_fd_sc_hd__dlclkp_1
X_06018_ _13902_/X wr vssd1 vssd1 vccd1 vccd1 _06018_/X sky130_fd_sc_hd__and2_1
XFILLER_58_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09406__D line[119] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[5\].CLKBUF\[1\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XOVHB\[0\].VALID\[13\].FF OVHB\[0\].V/CLK A[20] vssd1 vssd1 vccd1 vccd1 OVHB\[0\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_87_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07969_ _07975_/CLK line[102] vssd1 vssd1 vccd1 vccd1 _07970_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_101_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09708_ _09708_/A _09729_/Y vssd1 vssd1 vccd1 vccd1 _13628_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_114_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10980_ _10980_/A _10989_/Y vssd1 vssd1 vccd1 vccd1 _13780_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[31\].CLKBUF\[3\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09639_ _09655_/CLK line[97] vssd1 vssd1 vccd1 vccd1 _09640_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_83_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11671__D line[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12650_ _12650_/A _12669_/Y vssd1 vssd1 vccd1 vccd1 _13770_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06765__D line[78] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09141__D line[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11601_ _11615_/CLK line[98] vssd1 vssd1 vccd1 vccd1 _11602_/A sky130_fd_sc_hd__dfxtp_1
XPHY_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12581_ _12595_/CLK line[34] vssd1 vssd1 vccd1 vccd1 _12582_/A sky130_fd_sc_hd__dfxtp_1
XPHY_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[1\].VALID\[3\].TOBUF OVHB\[1\].VALID\[3\].FF/Q OVHB\[1\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04919_/B2 sky130_fd_sc_hd__ebufn_2
XPHY_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08980__D line[52] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11532_ _11532_/A _11549_/Y vssd1 vssd1 vccd1 vccd1 _13772_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13598__D line[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XOVHB\[26\].VALID\[6\].TOBUF OVHB\[26\].VALID\[6\].FF/Q OVHB\[26\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04923_/A2 sky130_fd_sc_hd__ebufn_2
X_11463_ _11475_/CLK line[35] vssd1 vssd1 vccd1 vccd1 _11464_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13202_ _13202_/A _13229_/Y vssd1 vssd1 vccd1 vccd1 _13762_/Z sky130_fd_sc_hd__ebufn_2
X_10414_ _10414_/A _10429_/Y vssd1 vssd1 vccd1 vccd1 _13774_/Z sky130_fd_sc_hd__ebufn_2
X_11394_ _11394_/A _11409_/Y vssd1 vssd1 vccd1 vccd1 _13634_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__04930__A2_N _04930_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13133_ _13155_/CLK line[45] vssd1 vssd1 vccd1 vccd1 _13134_/A sky130_fd_sc_hd__dfxtp_1
X_10345_ _10355_/CLK line[36] vssd1 vssd1 vccd1 vccd1 _10346_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12007__D line[42] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06005__D line[100] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13064_ _13064_/A _13089_/Y vssd1 vssd1 vccd1 vccd1 _13624_/Z sky130_fd_sc_hd__ebufn_2
X_10276_ _10276_/A _10289_/Y vssd1 vssd1 vccd1 vccd1 _13636_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11846__D line[82] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12015_ _12035_/CLK line[46] vssd1 vssd1 vccd1 vccd1 _12016_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[19\].CG clk OVHB\[19\].CGAND/X vssd1 vssd1 vccd1 vccd1 OVHB\[19\].V/CLK sky130_fd_sc_hd__dlclkp_1
XDATA\[13\].CLKBUF\[4\] clk vssd1 vssd1 vccd1 vccd1 _06227_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_120_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09316__D line[92] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08220__D line[89] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13966_ _13971_/C _13971_/A _13971_/B _13971_/D vssd1 vssd1 vccd1 vccd1 _13966_/X
+ sky130_fd_sc_hd__and4bb_4
X_12917_ _12945_/CLK line[74] vssd1 vssd1 vccd1 vccd1 _12918_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[24\].VALID\[11\].FF OVHB\[24\].V/CLK A[18] vssd1 vssd1 vccd1 vccd1 OVHB\[24\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_80_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13897_ A[4] vssd1 vssd1 vccd1 vccd1 _13905_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_0_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12848_ _12848_/A _12879_/Y vssd1 vssd1 vccd1 vccd1 _13688_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_15_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10197__D line[111] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12779_ _12805_/CLK line[11] vssd1 vssd1 vccd1 vccd1 _12780_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05320_ _05350_/CLK line[48] vssd1 vssd1 vccd1 vccd1 _05321_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08890__D line[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05251_ _05251_/A _05284_/Y vssd1 vssd1 vccd1 vccd1 _13651_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_175_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05182_ _05210_/CLK line[122] vssd1 vssd1 vccd1 vccd1 _05183_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_127_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09990_ _09990_/A _10009_/Y vssd1 vssd1 vccd1 vccd1 _13630_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_170_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[12\].VALID\[9\].FF_D A[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08941_ _08955_/CLK line[34] vssd1 vssd1 vccd1 vccd1 _08942_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_130_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10660__D line[52] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[14\].VALID\[13\].FF OVHB\[14\].V/CLK A[20] vssd1 vssd1 vccd1 vccd1 OVHB\[14\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_08872_ _08872_/A _08889_/Y vssd1 vssd1 vccd1 vccd1 _13632_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05754__D line[113] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08130__D line[62] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07823_ _07835_/CLK line[35] vssd1 vssd1 vccd1 vccd1 _07824_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05109__A _13931_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07754_ _07754_/A _07769_/Y vssd1 vssd1 vccd1 vccd1 _13634_/Z sky130_fd_sc_hd__ebufn_2
X_04966_ _04966_/A _04969_/Y vssd1 vssd1 vccd1 vccd1 _13646_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[1\].VALID\[10\].FF_D A[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDATA\[12\].CLKBUF\[1\] clk vssd1 vssd1 vccd1 vccd1 _05842_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_37_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06705_ _06715_/CLK line[36] vssd1 vssd1 vccd1 vccd1 _06706_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12587__D line[37] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07685_ _07695_/CLK line[100] vssd1 vssd1 vccd1 vccd1 _07686_/A sky130_fd_sc_hd__dfxtp_1
X_09424_ _09424_/A _09449_/Y vssd1 vssd1 vccd1 vccd1 _13624_/Z sky130_fd_sc_hd__ebufn_2
X_06636_ _06636_/A _06649_/Y vssd1 vssd1 vccd1 vccd1 _13636_/Z sky130_fd_sc_hd__ebufn_2
X_09355_ _09375_/CLK line[110] vssd1 vssd1 vccd1 vccd1 _09356_/A sky130_fd_sc_hd__dfxtp_1
X_06567_ _06575_/CLK line[101] vssd1 vssd1 vccd1 vccd1 _06568_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07978__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09896__D line[87] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08306_ _08306_/A _08329_/Y vssd1 vssd1 vccd1 vccd1 _13626_/Z sky130_fd_sc_hd__ebufn_2
X_05518_ _05518_/A _05529_/Y vssd1 vssd1 vccd1 vccd1 _13638_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09286_ _09286_/A _09309_/Y vssd1 vssd1 vccd1 vccd1 _13766_/Z sky130_fd_sc_hd__ebufn_2
X_06498_ _06498_/A _06509_/Y vssd1 vssd1 vccd1 vccd1 _13778_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_21_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10835__D line[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08237_ _08255_/CLK line[111] vssd1 vssd1 vccd1 vccd1 _08238_/A sky130_fd_sc_hd__dfxtp_1
X_05449_ _05455_/CLK line[102] vssd1 vssd1 vccd1 vccd1 _05450_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13211__D line[66] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05929__D line[65] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08305__D line[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08168_ _08168_/A _08189_/Y vssd1 vssd1 vccd1 vccd1 _13768_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[10\].CLKBUF\[3\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07119_ _07135_/CLK line[97] vssd1 vssd1 vccd1 vccd1 _07120_/A sky130_fd_sc_hd__dfxtp_1
X_08099_ _08115_/CLK line[33] vssd1 vssd1 vccd1 vccd1 _08100_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_133_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XOVHB\[24\].VALID\[0\].FF OVHB\[24\].V/CLK A[7] vssd1 vssd1 vccd1 vccd1 OVHB\[24\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_69_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10130_ _10130_/A _10149_/Y vssd1 vssd1 vccd1 vccd1 _13770_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06403__A _13904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10570__D line[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10061_ _10075_/CLK line[34] vssd1 vssd1 vccd1 vccd1 _10062_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[0\].VALID\[0\].FF_D A[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13820_ _13820_/CLK line[89] vssd1 vssd1 vccd1 vccd1 _13821_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_28_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12497__D line[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13751_ _13751_/A _13754_/Y vssd1 vssd1 vccd1 vccd1 _13751_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_16_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10963_ _10985_/CLK line[77] vssd1 vssd1 vccd1 vccd1 _10964_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[31\].CGAND _13927_/X wr vssd1 vssd1 vccd1 vccd1 OVHB\[31\].CGAND/X sky130_fd_sc_hd__and2_4
X_12702_ _12702_/CLK _12703_/X vssd1 vssd1 vccd1 vccd1 _12700_/CLK sky130_fd_sc_hd__dlclkp_1
XANTENNA_DATA\[3\].CLKBUF\[3\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06495__D line[68] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13682_ _13682_/CLK _13683_/X vssd1 vssd1 vccd1 vccd1 _13680_/CLK sky130_fd_sc_hd__dlclkp_1
X_10894_ _10894_/A _10919_/Y vssd1 vssd1 vccd1 vccd1 _13694_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_71_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12633_ _13936_/X wr vssd1 vssd1 vccd1 vccd1 _12633_/X sky130_fd_sc_hd__and2_1
XPHY_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12564_ _13936_/X vssd1 vssd1 vccd1 vccd1 _12564_/Y sky130_fd_sc_hd__inv_2
XPHY_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10745__D line[96] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11515_ _11545_/CLK line[64] vssd1 vssd1 vccd1 vccd1 _11516_/A sky130_fd_sc_hd__dfxtp_1
XPHY_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12495_ _12525_/CLK line[0] vssd1 vssd1 vccd1 vccd1 _12496_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_156_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11446_ _11446_/A _11479_/Y vssd1 vssd1 vccd1 vccd1 _13686_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_144_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_OVHB\[25\].VALID\[9\].FF_D A[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12960__D line[94] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11377_ _11405_/CLK line[10] vssd1 vssd1 vccd1 vccd1 _11378_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_125_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13116_ _13120_/CLK line[23] vssd1 vssd1 vccd1 vccd1 _13117_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_125_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10328_ _10328_/A _10359_/Y vssd1 vssd1 vccd1 vccd1 _13688_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_112_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11576__D line[87] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13047_ _13047_/A _13054_/Y vssd1 vssd1 vccd1 vccd1 _13887_/Z sky130_fd_sc_hd__ebufn_2
X_10259_ _10285_/CLK line[11] vssd1 vssd1 vccd1 vccd1 _10260_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_79_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09046__D line[82] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09624__A _13920_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08885__D line[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09343__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[22\].VALID\[2\].FF OVHB\[22\].V/CLK A[9] vssd1 vssd1 vccd1 vccd1 OVHB\[22\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_19_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13949_ _13949_/A _13949_/B _13949_/C _13949_/D vssd1 vssd1 vccd1 vccd1 _13949_/X
+ sky130_fd_sc_hd__and4_4
XANTENNA__12200__D line[116] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07470_ _07470_/A _07489_/Y vssd1 vssd1 vccd1 vccd1 _13630_/Z sky130_fd_sc_hd__ebufn_2
X_06421_ _06435_/CLK line[34] vssd1 vssd1 vccd1 vccd1 _06422_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_201_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[3\].VALID\[14\].TOBUF OVHB\[3\].VALID\[14\].FF/Q OVHB\[3\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_201_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09140_ _09140_/A _09169_/Y vssd1 vssd1 vccd1 vccd1 _13620_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05599__A _13901_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06352_ _06352_/A _06369_/Y vssd1 vssd1 vccd1 vccd1 _13632_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_30_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05303_ _05315_/CLK line[35] vssd1 vssd1 vccd1 vccd1 _05304_/A sky130_fd_sc_hd__dfxtp_1
X_09071_ _09095_/CLK line[108] vssd1 vssd1 vccd1 vccd1 _09072_/A sky130_fd_sc_hd__dfxtp_1
X_06283_ _06295_/CLK line[99] vssd1 vssd1 vccd1 vccd1 _06284_/A sky130_fd_sc_hd__dfxtp_1
X_08022_ _08022_/A _08049_/Y vssd1 vssd1 vccd1 vccd1 _13622_/Z sky130_fd_sc_hd__ebufn_2
X_05234_ _05234_/A _05249_/Y vssd1 vssd1 vccd1 vccd1 _13634_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[8\].VALID\[3\].TOBUF OVHB\[8\].VALID\[3\].FF/Q OVHB\[8\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04919_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_190_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05165_ _05175_/CLK line[100] vssd1 vssd1 vccd1 vccd1 _05166_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[6\].VALID\[14\].FF_D A[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09518__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09973_ _13921_/X wr vssd1 vssd1 vccd1 vccd1 _09973_/X sky130_fd_sc_hd__and2_1
X_05096_ _05096_/A _05109_/Y vssd1 vssd1 vccd1 vccd1 _13776_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11486__D line[60] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10390__D line[57] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08924_ _13915_/X vssd1 vssd1 vccd1 vccd1 _08924_/Y sky130_fd_sc_hd__inv_2
XANTENNA__05484__D line[118] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08855_ _08885_/CLK line[0] vssd1 vssd1 vccd1 vccd1 _08856_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_69_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[23\].VALID\[10\].TOBUF OVHB\[23\].VALID\[10\].FF/Q OVHB\[23\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04932_/B2 sky130_fd_sc_hd__ebufn_2
X_07806_ _07806_/A _07839_/Y vssd1 vssd1 vccd1 vccd1 _13686_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08795__D line[110] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08786_ _08786_/A _08819_/Y vssd1 vssd1 vccd1 vccd1 _13826_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_55_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05998_ _05998_/A _06019_/Y vssd1 vssd1 vccd1 vccd1 _13838_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[6\].VALID\[4\].FF_D A[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07737_ _07765_/CLK line[10] vssd1 vssd1 vccd1 vccd1 _07738_/A sky130_fd_sc_hd__dfxtp_1
X_04949_ _04965_/CLK line[1] vssd1 vssd1 vccd1 vccd1 _04950_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12110__D line[80] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06893__A _13905_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07668_ _07668_/A _07699_/Y vssd1 vssd1 vccd1 vccd1 _13828_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_52_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09407_ _09407_/A _09414_/Y vssd1 vssd1 vccd1 vccd1 _13887_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_40_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06619_ _06645_/CLK line[11] vssd1 vssd1 vccd1 vccd1 _06620_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_25_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_DATA\[28\].CLKBUF\[6\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07599_ _07625_/CLK line[75] vssd1 vssd1 vccd1 vccd1 _07600_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[20\].VALID\[4\].FF OVHB\[20\].V/CLK A[11] vssd1 vssd1 vccd1 vccd1 OVHB\[20\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__11304__A _13933_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09338_ _09340_/CLK line[88] vssd1 vssd1 vccd1 vccd1 _09339_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_21_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10565__D line[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11023__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09269_ _09269_/A _09274_/Y vssd1 vssd1 vccd1 vccd1 _13749_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_5_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05659__D line[70] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[10\].VALID\[11\].FF OVHB\[10\].V/CLK A[18] vssd1 vssd1 vccd1 vccd1 OVHB\[10\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_11300_ _11300_/CLK line[89] vssd1 vssd1 vccd1 vccd1 _11301_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08035__D line[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12280_ _12280_/CLK line[25] vssd1 vssd1 vccd1 vccd1 _12281_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_112_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13876__D line[114] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11231_ _11231_/A _11234_/Y vssd1 vssd1 vccd1 vccd1 _13751_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_181_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11162_ _11162_/CLK _11163_/X vssd1 vssd1 vccd1 vccd1 _11160_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_136_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10113_ _13922_/X wr vssd1 vssd1 vccd1 vccd1 _10113_/X sky130_fd_sc_hd__and2_1
X_11093_ _13925_/X wr vssd1 vssd1 vccd1 vccd1 _11093_/X sky130_fd_sc_hd__and2_1
XANTENNA__05394__D line[91] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10044_ _13922_/X vssd1 vssd1 vccd1 vccd1 _10044_/Y sky130_fd_sc_hd__inv_2
XFILLER_102_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__04915__A1_N A_h[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13803_ _13803_/A _13824_/Y vssd1 vssd1 vccd1 vccd1 _13803_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__04923__A2 _04923_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11995_ _11995_/A _12004_/Y vssd1 vssd1 vccd1 vccd1 _13675_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13116__D line[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13734_ _13750_/CLK line[49] vssd1 vssd1 vccd1 vccd1 _13735_/A sky130_fd_sc_hd__dfxtp_1
X_10946_ _10950_/CLK line[55] vssd1 vssd1 vccd1 vccd1 _10947_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_32_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_OVHB\[8\].VALID\[10\].FF_D A[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[19\].VALID\[5\].FF OVHB\[19\].V/CLK A[12] vssd1 vssd1 vccd1 vccd1 OVHB\[19\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_13665_ _13665_/A _13684_/Y vssd1 vssd1 vccd1 vccd1 _13665_/Z sky130_fd_sc_hd__ebufn_2
X_10877_ _10877_/A _10884_/Y vssd1 vssd1 vccd1 vccd1 _13677_/Z sky130_fd_sc_hd__ebufn_2
X_12616_ _12630_/CLK line[50] vssd1 vssd1 vccd1 vccd1 _12617_/A sky130_fd_sc_hd__dfxtp_1
XPHY_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13596_ _13610_/CLK line[114] vssd1 vssd1 vccd1 vccd1 _13597_/A sky130_fd_sc_hd__dfxtp_1
XPHY_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10475__D line[110] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12547_ _12547_/A _12564_/Y vssd1 vssd1 vccd1 vccd1 _13667_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[1\].CLKBUF\[5\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05569__D line[43] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12478_ _12490_/CLK line[115] vssd1 vssd1 vccd1 vccd1 _12479_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12690__D line[84] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11429_ _11429_/A _11444_/Y vssd1 vssd1 vccd1 vccd1 _13669_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_172_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07784__D line[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07139__A _13909_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06970_ _06970_/A _06999_/Y vssd1 vssd1 vccd1 vccd1 _13690_/Z sky130_fd_sc_hd__ebufn_2
X_05921_ _05945_/CLK line[76] vssd1 vssd1 vccd1 vccd1 _05922_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_MUX.M\[2\].MUX\[0\]_A2 _13791_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08640_ _08640_/CLK line[25] vssd1 vssd1 vccd1 vccd1 _08641_/A sky130_fd_sc_hd__dfxtp_1
X_05852_ _05852_/A _05879_/Y vssd1 vssd1 vccd1 vccd1 _13692_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_94_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08571_ _08571_/A _08574_/Y vssd1 vssd1 vccd1 vccd1 _13891_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__04914__A2 _04922_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05783_ _05805_/CLK line[13] vssd1 vssd1 vccd1 vccd1 _05784_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_54_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[6\].VALID\[8\].TOBUF OVHB\[6\].VALID\[8\].FF/Q OVHB\[6\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04931_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__13026__D line[124] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07522_ _07522_/CLK _07523_/X vssd1 vssd1 vccd1 vccd1 _07520_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_35_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07024__D line[54] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12865__D line[36] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07453_ _13910_/X wr vssd1 vssd1 vccd1 vccd1 _07453_/X sky130_fd_sc_hd__and2_1
XFILLER_195_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07959__D line[97] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06404_ _13904_/X vssd1 vssd1 vccd1 vccd1 _06404_/Y sky130_fd_sc_hd__inv_2
X_07384_ _13910_/X vssd1 vssd1 vccd1 vccd1 _07384_/Y sky130_fd_sc_hd__inv_2
XFILLER_176_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09123_ _09123_/A _09134_/Y vssd1 vssd1 vccd1 vccd1 _13883_/Z sky130_fd_sc_hd__ebufn_2
X_06335_ _06365_/CLK line[0] vssd1 vssd1 vccd1 vccd1 _06336_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_175_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09054_ _09060_/CLK line[86] vssd1 vssd1 vccd1 vccd1 _09055_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[17\].VALID\[7\].FF OVHB\[17\].V/CLK A[14] vssd1 vssd1 vccd1 vccd1 OVHB\[17\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_06266_ _06266_/A _06299_/Y vssd1 vssd1 vccd1 vccd1 _13826_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08433__A _13913_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08005_ _08005_/A _08014_/Y vssd1 vssd1 vccd1 vccd1 _13885_/Z sky130_fd_sc_hd__ebufn_2
X_05217_ _05245_/CLK line[10] vssd1 vssd1 vccd1 vccd1 _05218_/A sky130_fd_sc_hd__dfxtp_1
X_06197_ _06225_/CLK line[74] vssd1 vssd1 vccd1 vccd1 _06198_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[5\].VALID\[13\].FF OVHB\[5\].V/CLK A[20] vssd1 vssd1 vccd1 vccd1 OVHB\[5\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_2_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05148_ _05148_/A _05179_/Y vssd1 vssd1 vccd1 vccd1 _13828_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_104_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11794__A _13927_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12105__D line[73] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09956_ _09970_/CLK line[114] vssd1 vssd1 vccd1 vccd1 _09957_/A sky130_fd_sc_hd__dfxtp_1
X_05079_ _05105_/CLK line[75] vssd1 vssd1 vccd1 vccd1 _05080_/A sky130_fd_sc_hd__dfxtp_1
X_08907_ _08907_/A _08924_/Y vssd1 vssd1 vccd1 vccd1 _13667_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_66_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09887_ _09887_/A _09904_/Y vssd1 vssd1 vccd1 vccd1 _13807_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_100_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XDATA\[3\].CLKBUF\[5\] clk vssd1 vssd1 vccd1 vccd1 _12142_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_85_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08838_ _08850_/CLK line[115] vssd1 vssd1 vccd1 vccd1 _08839_/A sky130_fd_sc_hd__dfxtp_1
X_08769_ _08769_/A _08784_/Y vssd1 vssd1 vccd1 vccd1 _13809_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_122_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10800_ _10810_/CLK line[116] vssd1 vssd1 vccd1 vccd1 _10801_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_122_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11780_ _11790_/CLK line[52] vssd1 vssd1 vccd1 vccd1 _11781_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08608__A _13914_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10731_ _10731_/A _10744_/Y vssd1 vssd1 vccd1 vccd1 _13811_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12775__D line[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13450_ _13470_/CLK line[62] vssd1 vssd1 vccd1 vccd1 _13451_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06773__D line[67] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10662_ _10670_/CLK line[53] vssd1 vssd1 vccd1 vccd1 _10663_/A sky130_fd_sc_hd__dfxtp_1
X_12401_ _12401_/A _12424_/Y vssd1 vssd1 vccd1 vccd1 _13801_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11969__A _13934_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13381_ _13381_/A _13404_/Y vssd1 vssd1 vccd1 vccd1 _13661_/Z sky130_fd_sc_hd__ebufn_2
X_10593_ _10593_/A _10604_/Y vssd1 vssd1 vccd1 vccd1 _13673_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[13\].VALID\[3\].TOBUF OVHB\[13\].VALID\[3\].FF/Q OVHB\[13\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04919_/B2 sky130_fd_sc_hd__ebufn_2
X_12332_ _12350_/CLK line[63] vssd1 vssd1 vccd1 vccd1 _12333_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11688__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12263_ _12263_/A _12284_/Y vssd1 vssd1 vccd1 vccd1 _13663_/Z sky130_fd_sc_hd__ebufn_2
X_11214_ _11230_/CLK line[49] vssd1 vssd1 vccd1 vccd1 _11215_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_122_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12194_ _12210_/CLK line[113] vssd1 vssd1 vccd1 vccd1 _12195_/A sky130_fd_sc_hd__dfxtp_1
X_11145_ _11145_/A _11164_/Y vssd1 vssd1 vccd1 vccd1 _13665_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12015__D line[46] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07109__D line[107] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[15\].VALID\[9\].FF OVHB\[15\].V/CLK A[16] vssd1 vssd1 vccd1 vccd1 OVHB\[15\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XOVHB\[29\].VALID\[11\].FF OVHB\[29\].V/CLK A[18] vssd1 vssd1 vccd1 vccd1 OVHB\[29\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_110_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06013__D line[104] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11076_ _11090_/CLK line[114] vssd1 vssd1 vccd1 vccd1 _11077_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_48_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11854__D line[86] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10027_ _10027_/A _10044_/Y vssd1 vssd1 vccd1 vccd1 _13667_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06948__D line[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10113__A _13922_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09324__D line[81] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[11\].VALID\[0\].FF_D A[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11978_ _12000_/CLK line[29] vssd1 vssd1 vccd1 vccd1 _11979_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[2\].CLKBUF\[2\] clk vssd1 vssd1 vccd1 vccd1 _11197_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_16_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13717_ _13717_/CLK _13718_/X vssd1 vssd1 vccd1 vccd1 _13715_/CLK sky130_fd_sc_hd__dlclkp_1
X_10929_ _10929_/A _10954_/Y vssd1 vssd1 vccd1 vccd1 _13729_/Z sky130_fd_sc_hd__ebufn_2
X_13648_ _13899_/X wr vssd1 vssd1 vccd1 vccd1 _13648_/X sky130_fd_sc_hd__and2_1
XFILLER_158_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13579_ _13898_/Y vssd1 vssd1 vccd1 vccd1 _13579_/Y sky130_fd_sc_hd__inv_2
XOVHB\[1\].CG clk OVHB\[1\].CGAND/X vssd1 vssd1 vccd1 vccd1 OVHB\[1\].V/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05299__D line[33] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06120_ _06120_/CLK line[25] vssd1 vssd1 vccd1 vccd1 _06121_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_118_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XOVHB\[19\].VALID\[13\].FF OVHB\[19\].V/CLK A[20] vssd1 vssd1 vccd1 vccd1 OVHB\[19\].VALID\[13\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_145_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06051_ _06051_/A _06054_/Y vssd1 vssd1 vccd1 vccd1 _13891_/Z sky130_fd_sc_hd__ebufn_2
X_05002_ _05002_/CLK _05003_/X vssd1 vssd1 vccd1 vccd1 _05000_/CLK sky130_fd_sc_hd__dlclkp_1
XOVHB\[18\].VOBUF OVHB\[18\].V/Q OVHB\[18\].INV/Y vssd1 vssd1 vccd1 vccd1 _04912_/B1
+ sky130_fd_sc_hd__ebufn_2
X_09810_ _09830_/CLK line[62] vssd1 vssd1 vccd1 vccd1 _09811_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_141_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09741_ _09741_/A _09764_/Y vssd1 vssd1 vccd1 vccd1 _13661_/Z sky130_fd_sc_hd__ebufn_2
X_06953_ _06953_/A _06964_/Y vssd1 vssd1 vccd1 vccd1 _13673_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[2\].VALID\[7\].FF_D A[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11764__D line[59] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDATA\[22\].CLKBUF\[6\] clk vssd1 vssd1 vccd1 vccd1 _09097_/CLK sky130_fd_sc_hd__clkbuf_4
X_05904_ _05910_/CLK line[54] vssd1 vssd1 vccd1 vccd1 _05905_/A sky130_fd_sc_hd__dfxtp_1
X_09672_ _09690_/CLK line[127] vssd1 vssd1 vccd1 vccd1 _09673_/A sky130_fd_sc_hd__dfxtp_1
X_06884_ _06890_/CLK line[118] vssd1 vssd1 vccd1 vccd1 _06885_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05762__D line[117] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08623_ _08623_/A _08644_/Y vssd1 vssd1 vccd1 vccd1 _13663_/Z sky130_fd_sc_hd__ebufn_2
X_05835_ _05835_/A _05844_/Y vssd1 vssd1 vccd1 vccd1 _13675_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_MUX.M\[1\].MUX\[1\]_A0 _13646_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13334__A _13938_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08554_ _08570_/CLK line[113] vssd1 vssd1 vccd1 vccd1 _08555_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05766_ _05770_/CLK line[119] vssd1 vssd1 vccd1 vccd1 _05767_/A sky130_fd_sc_hd__dfxtp_1
X_07505_ _07505_/A _07524_/Y vssd1 vssd1 vccd1 vccd1 _13665_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12595__D line[41] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13053__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08485_ _08485_/A _08504_/Y vssd1 vssd1 vccd1 vccd1 _13805_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05697_ _05697_/A _05704_/Y vssd1 vssd1 vccd1 vccd1 _13817_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07689__D line[102] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07436_ _07450_/CLK line[114] vssd1 vssd1 vccd1 vccd1 _07437_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_167_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07367_ _07367_/A _07384_/Y vssd1 vssd1 vccd1 vccd1 _13807_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11004__D line[81] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09106_ _09130_/CLK line[124] vssd1 vssd1 vccd1 vccd1 _09107_/A sky130_fd_sc_hd__dfxtp_1
X_06318_ _06330_/CLK line[115] vssd1 vssd1 vccd1 vccd1 _06319_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_148_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07298_ _07310_/CLK line[51] vssd1 vssd1 vccd1 vccd1 _07299_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11939__D line[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10843__D line[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09037_ _09037_/A _09064_/Y vssd1 vssd1 vccd1 vccd1 _13797_/Z sky130_fd_sc_hd__ebufn_2
X_06249_ _06249_/A _06264_/Y vssd1 vssd1 vccd1 vccd1 _13809_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__05937__D line[69] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08313__D line[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13509__A _13898_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13228__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09939_ _13921_/X vssd1 vssd1 vccd1 vccd1 _09939_/Y sky130_fd_sc_hd__inv_2
XANTENNA_OVHB\[21\].V_D TIE/HI vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[24\].VALID\[0\].FF_D A[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12950_ _12980_/CLK line[80] vssd1 vssd1 vccd1 vccd1 _12951_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_133_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05672__D line[90] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[11\].VALID\[8\].TOBUF OVHB\[11\].VALID\[8\].FF/Q OVHB\[11\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04931_/B2 sky130_fd_sc_hd__ebufn_2
X_11901_ _11901_/A _11934_/Y vssd1 vssd1 vccd1 vccd1 _13861_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_45_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12881_ _12881_/A _12914_/Y vssd1 vssd1 vccd1 vccd1 _13721_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_133_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11832_ _11860_/CLK line[90] vssd1 vssd1 vccd1 vccd1 _11833_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[21\].CLKBUF\[3\] clk vssd1 vssd1 vccd1 vccd1 _08712_/CLK sky130_fd_sc_hd__clkbuf_4
XFILLER_54_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11763_ _11763_/A _11794_/Y vssd1 vssd1 vccd1 vccd1 _13723_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_159_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_OVHB\[17\].VALID\[4\].FF_D A[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07599__D line[75] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10714_ _10740_/CLK line[91] vssd1 vssd1 vccd1 vccd1 _10715_/A sky130_fd_sc_hd__dfxtp_1
X_13502_ _13502_/A _13509_/Y vssd1 vssd1 vccd1 vccd1 _13782_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11694_ _11720_/CLK line[27] vssd1 vssd1 vccd1 vccd1 _11695_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[1\].VALID\[11\].FF OVHB\[1\].V/CLK A[18] vssd1 vssd1 vccd1 vccd1 OVHB\[1\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_13433_ _13435_/CLK line[40] vssd1 vssd1 vccd1 vccd1 _13434_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10645_ _10645_/A _10674_/Y vssd1 vssd1 vccd1 vccd1 _13725_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09169__A _13916_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13364_ _13364_/A _13369_/Y vssd1 vssd1 vccd1 vccd1 _13644_/Z sky130_fd_sc_hd__ebufn_2
X_10576_ _10600_/CLK line[28] vssd1 vssd1 vccd1 vccd1 _10577_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_139_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10753__D line[109] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12315_ _12315_/CLK line[41] vssd1 vssd1 vccd1 vccd1 _12316_/A sky130_fd_sc_hd__dfxtp_1
X_13295_ _13295_/CLK line[105] vssd1 vssd1 vccd1 vccd1 _13296_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05847__D line[42] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12246_ _12246_/A _12249_/Y vssd1 vssd1 vccd1 vccd1 _13646_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_142_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12177_ _12177_/CLK _12178_/X vssd1 vssd1 vccd1 vccd1 _12175_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_96_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11128_ _13933_/X wr vssd1 vssd1 vccd1 vccd1 _11128_/X sky130_fd_sc_hd__and2_1
XFILLER_68_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[8\].VALID\[2\].FF OVHB\[8\].V/CLK A[9] vssd1 vssd1 vccd1 vccd1 OVHB\[8\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[24\].CG_CLK clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06678__D line[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11059_ _13925_/X vssd1 vssd1 vccd1 vccd1 _11059_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09054__D line[86] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[20\].CLKBUF\[1\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10778__A _13924_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09989__D line[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05620_ _05630_/CLK line[52] vssd1 vssd1 vccd1 vccd1 _05621_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_91_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05551_ _05551_/A _05564_/Y vssd1 vssd1 vccd1 vccd1 _13671_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10928__D line[61] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13304__D line[123] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08270_ _08290_/CLK line[126] vssd1 vssd1 vccd1 vccd1 _08271_/A sky130_fd_sc_hd__dfxtp_1
X_05482_ _05490_/CLK line[117] vssd1 vssd1 vccd1 vccd1 _05483_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07302__D line[53] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07221_ _07221_/A _07244_/Y vssd1 vssd1 vccd1 vccd1 _13661_/Z sky130_fd_sc_hd__ebufn_2
XDATA\[20\].CLKBUF\[0\] clk vssd1 vssd1 vccd1 vccd1 _08327_/CLK sky130_fd_sc_hd__clkbuf_4
XOVHB\[16\].VALID\[14\].TOBUF OVHB\[16\].VALID\[14\].FF/Q OVHB\[16\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_192_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07152_ _07170_/CLK line[127] vssd1 vssd1 vccd1 vccd1 _07153_/A sky130_fd_sc_hd__dfxtp_1
XDATA\[10\].CLKBUF\[6\] clk vssd1 vssd1 vccd1 vccd1 _05457_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA_OVHB\[15\].VALID\[12\].FF_D A[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06103_ _06103_/A _06124_/Y vssd1 vssd1 vccd1 vccd1 _13663_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_145_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07083_ _07083_/A _07104_/Y vssd1 vssd1 vccd1 vccd1 _13803_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09229__D line[38] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06034_ _06050_/CLK line[113] vssd1 vssd1 vccd1 vccd1 _06035_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_141_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07985_ _07985_/A _08014_/Y vssd1 vssd1 vccd1 vccd1 _13865_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11494__D line[49] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09724_ _09724_/A _09729_/Y vssd1 vssd1 vccd1 vccd1 _13644_/Z sky130_fd_sc_hd__ebufn_2
X_06936_ _06960_/CLK line[28] vssd1 vssd1 vccd1 vccd1 _06937_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06588__D line[125] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[25\].VALID\[11\].FF_D A[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09655_ _09655_/CLK line[105] vssd1 vssd1 vccd1 vccd1 _09656_/A sky130_fd_sc_hd__dfxtp_1
X_06867_ _06867_/A _06894_/Y vssd1 vssd1 vccd1 vccd1 _13867_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_28_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08606_ _08606_/A _08609_/Y vssd1 vssd1 vccd1 vccd1 _13646_/Z sky130_fd_sc_hd__ebufn_2
X_05818_ _05840_/CLK line[29] vssd1 vssd1 vccd1 vccd1 _05819_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_43_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09586_ _09586_/A _09589_/Y vssd1 vssd1 vccd1 vccd1 _13786_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_63_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06798_ _06820_/CLK line[93] vssd1 vssd1 vccd1 vccd1 _06799_/A sky130_fd_sc_hd__dfxtp_1
XPHY_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08537_ _08537_/CLK _08538_/X vssd1 vssd1 vccd1 vccd1 _08535_/CLK sky130_fd_sc_hd__dlclkp_1
XPHY_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05749_ _05749_/A _05774_/Y vssd1 vssd1 vccd1 vccd1 _13869_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[6\].VALID\[4\].FF OVHB\[6\].V/CLK A[11] vssd1 vssd1 vccd1 vccd1 OVHB\[6\].VALID\[4\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XOVHB\[15\].VALID\[11\].FF OVHB\[15\].V/CLK A[18] vssd1 vssd1 vccd1 vccd1 OVHB\[15\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XPHY_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08468_ _13913_/X wr vssd1 vssd1 vccd1 vccd1 _08468_/X sky130_fd_sc_hd__and2_1
XPHY_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07212__D line[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07419_ _13910_/X vssd1 vssd1 vccd1 vccd1 _07419_/Y sky130_fd_sc_hd__inv_2
XFILLER_50_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08399_ _13913_/X vssd1 vssd1 vccd1 vccd1 _08399_/Y sky130_fd_sc_hd__inv_2
XPHY_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[6\].V_D TIE/HI vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10430_ _10460_/CLK line[80] vssd1 vssd1 vccd1 vccd1 _10431_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_12_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11669__D line[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10361_ _10361_/A _10394_/Y vssd1 vssd1 vccd1 vccd1 _13721_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_128_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09139__D line[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12100_ _12100_/A _12109_/Y vssd1 vssd1 vccd1 vccd1 _13780_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_124_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08043__D line[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13080_ _13080_/A _13089_/Y vssd1 vssd1 vccd1 vccd1 _13640_/Z sky130_fd_sc_hd__ebufn_2
X_10292_ _10320_/CLK line[26] vssd1 vssd1 vccd1 vccd1 _10293_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13884__D line[118] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12031_ _12035_/CLK line[39] vssd1 vssd1 vccd1 vccd1 _12032_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12143__A _13934_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08978__D line[51] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_DATA\[19\].CLKBUF\[2\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13982_ _13982_/A _13982_/B _13982_/C _13982_/D vssd1 vssd1 vccd1 vccd1 _13982_/X
+ sky130_fd_sc_hd__and4_4
XFILLER_46_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[26\].VALID\[2\].TOBUF OVHB\[26\].VALID\[2\].FF/Q OVHB\[26\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04930_/B2 sky130_fd_sc_hd__ebufn_2
X_12933_ _12945_/CLK line[67] vssd1 vssd1 vccd1 vccd1 _12934_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_73_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12864_ _12864_/A _12879_/Y vssd1 vssd1 vccd1 vccd1 _13704_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09602__D line[95] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11815_ _11825_/CLK line[68] vssd1 vssd1 vccd1 vccd1 _11816_/A sky130_fd_sc_hd__dfxtp_1
X_12795_ _12805_/CLK line[4] vssd1 vssd1 vccd1 vccd1 _12796_/A sky130_fd_sc_hd__dfxtp_1
XPHY_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11746_ _11746_/A _11759_/Y vssd1 vssd1 vccd1 vccd1 _13706_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08218__D line[88] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11677_ _11685_/CLK line[5] vssd1 vssd1 vccd1 vccd1 _11678_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12318__A _13935_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10628_ _10628_/A _10639_/Y vssd1 vssd1 vccd1 vccd1 _13708_/Z sky130_fd_sc_hd__ebufn_2
X_13416_ _13416_/A _13439_/Y vssd1 vssd1 vccd1 vccd1 _13696_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[4\].VALID\[6\].FF OVHB\[4\].V/CLK A[13] vssd1 vssd1 vccd1 vccd1 OVHB\[4\].VALID\[6\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__10483__D line[99] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13347_ _13365_/CLK line[15] vssd1 vssd1 vccd1 vccd1 _13348_/A sky130_fd_sc_hd__dfxtp_1
X_10559_ _10565_/CLK line[6] vssd1 vssd1 vccd1 vccd1 _10560_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_170_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MUX.M\[3\].MUX\[2\]_A2 _13793_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05577__D line[47] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[10\].INV _13944_/X vssd1 vssd1 vccd1 vccd1 OVHB\[10\].INV/Y sky130_fd_sc_hd__inv_2
X_13278_ _13278_/A _13299_/Y vssd1 vssd1 vccd1 vccd1 _13838_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[26\].CGAND _13922_/X wr vssd1 vssd1 vccd1 vccd1 OVHB\[26\].CGAND/X sky130_fd_sc_hd__and2_4
XANTENNA__13794__D line[91] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12229_ _12245_/CLK line[1] vssd1 vssd1 vccd1 vccd1 _12230_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_69_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07792__D line[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XOVHB\[25\].INV _13965_/X vssd1 vssd1 vccd1 vccd1 OVHB\[25\].INV/Y sky130_fd_sc_hd__inv_2
X_07770_ _07800_/CLK line[16] vssd1 vssd1 vccd1 vccd1 _07771_/A sky130_fd_sc_hd__dfxtp_1
X_04982_ _05000_/CLK line[31] vssd1 vssd1 vccd1 vccd1 _04983_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_37_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06201__D line[76] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06721_ _06721_/A _06754_/Y vssd1 vssd1 vccd1 vccd1 _13721_/Z sky130_fd_sc_hd__ebufn_2
X_09440_ _09440_/A _09449_/Y vssd1 vssd1 vccd1 vccd1 _13640_/Z sky130_fd_sc_hd__ebufn_2
X_06652_ _06680_/CLK line[26] vssd1 vssd1 vccd1 vccd1 _06653_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[18\].VALID\[8\].TOBUF OVHB\[18\].VALID\[8\].FF/Q OVHB\[18\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04931_/B2 sky130_fd_sc_hd__ebufn_2
X_05603_ _05603_/A _05634_/Y vssd1 vssd1 vccd1 vccd1 _13723_/Z sky130_fd_sc_hd__ebufn_2
X_09371_ _09375_/CLK line[103] vssd1 vssd1 vccd1 vccd1 _09372_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10658__D line[51] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06583_ _06583_/A _06614_/Y vssd1 vssd1 vccd1 vccd1 _13863_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_52_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13034__D line[113] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08322_ _08322_/A _08329_/Y vssd1 vssd1 vccd1 vccd1 _13642_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_178_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05534_ _05560_/CLK line[27] vssd1 vssd1 vccd1 vccd1 _05535_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08128__D line[61] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12873__D line[40] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08253_ _08255_/CLK line[104] vssd1 vssd1 vccd1 vccd1 _08254_/A sky130_fd_sc_hd__dfxtp_1
X_05465_ _05465_/A _05494_/Y vssd1 vssd1 vccd1 vccd1 _13865_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07967__D line[101] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07204_ _07204_/A _07209_/Y vssd1 vssd1 vccd1 vccd1 _13644_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_192_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08184_ _08184_/A _08189_/Y vssd1 vssd1 vccd1 vccd1 _13784_/Z sky130_fd_sc_hd__ebufn_2
X_05396_ _05420_/CLK line[92] vssd1 vssd1 vccd1 vccd1 _05397_/A sky130_fd_sc_hd__dfxtp_1
X_07135_ _07135_/CLK line[105] vssd1 vssd1 vccd1 vccd1 _07136_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_133_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07066_ _07066_/A _07069_/Y vssd1 vssd1 vccd1 vccd1 _13786_/Z sky130_fd_sc_hd__ebufn_2
X_06017_ _06017_/CLK _06018_/X vssd1 vssd1 vccd1 vccd1 _06015_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_99_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_OVHB\[12\].CGAND_A _13902_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[20\].VALID\[3\].FF_D A[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[2\].VALID\[8\].FF OVHB\[2\].V/CLK A[15] vssd1 vssd1 vccd1 vccd1 OVHB\[2\].VALID\[8\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__13209__D line[65] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07968_ _07968_/A _07979_/Y vssd1 vssd1 vccd1 vccd1 _13848_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_114_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09707_ _09725_/CLK line[15] vssd1 vssd1 vccd1 vccd1 _09708_/A sky130_fd_sc_hd__dfxtp_1
X_06919_ _06925_/CLK line[6] vssd1 vssd1 vccd1 vccd1 _06920_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_74_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07899_ _07905_/CLK line[70] vssd1 vssd1 vccd1 vccd1 _07900_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_55_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_OVHB\[13\].VALID\[7\].FF_D A[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09638_ _09638_/A _09659_/Y vssd1 vssd1 vccd1 vccd1 _13838_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_204_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05950__D line[80] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09569_ _09585_/CLK line[65] vssd1 vssd1 vccd1 vccd1 _09570_/A sky130_fd_sc_hd__dfxtp_1
XPHY_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11600_ _11600_/A _11619_/Y vssd1 vssd1 vccd1 vccd1 _13840_/Z sky130_fd_sc_hd__ebufn_2
XPHY_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12580_ _12580_/A _12599_/Y vssd1 vssd1 vccd1 vccd1 _13700_/Z sky130_fd_sc_hd__ebufn_2
XPHY_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12783__D line[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11531_ _11545_/CLK line[66] vssd1 vssd1 vccd1 vccd1 _11532_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_184_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07877__D line[74] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06781__D line[71] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11462_ _11462_/A _11479_/Y vssd1 vssd1 vccd1 vccd1 _13702_/Z sky130_fd_sc_hd__ebufn_2
XPHY_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11399__D line[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13201_ _13225_/CLK line[76] vssd1 vssd1 vccd1 vccd1 _13202_/A sky130_fd_sc_hd__dfxtp_1
X_10413_ _10425_/CLK line[67] vssd1 vssd1 vccd1 vccd1 _10414_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[24\].VALID\[7\].TOBUF OVHB\[24\].VALID\[7\].FF/Q OVHB\[24\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04922_/A2 sky130_fd_sc_hd__ebufn_2
X_11393_ _11405_/CLK line[3] vssd1 vssd1 vccd1 vccd1 _11394_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_152_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13132_ _13132_/A _13159_/Y vssd1 vssd1 vccd1 vccd1 _13692_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_109_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10344_ _10344_/A _10359_/Y vssd1 vssd1 vccd1 vccd1 _13704_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_124_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13063_ _13085_/CLK line[13] vssd1 vssd1 vccd1 vccd1 _13064_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_140_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[30\].VALID\[2\].FF OVHB\[30\].V/CLK A[9] vssd1 vssd1 vccd1 vccd1 OVHB\[30\].VALID\[2\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_10275_ _10285_/CLK line[4] vssd1 vssd1 vccd1 vccd1 _10276_/A sky130_fd_sc_hd__dfxtp_1
X_12014_ _12014_/A _12039_/Y vssd1 vssd1 vccd1 vccd1 _13694_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_66_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12023__D line[35] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07117__D line[111] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12958__D line[93] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13965_ _13971_/C _13971_/B _13971_/A _13971_/D vssd1 vssd1 vccd1 vccd1 _13965_/X
+ sky130_fd_sc_hd__and4bb_4
XANTENNA__06956__D line[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12916_ _12916_/A _12949_/Y vssd1 vssd1 vccd1 vccd1 _13756_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09332__D line[85] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13896_ A[3] vssd1 vssd1 vccd1 vccd1 _13905_/B sky130_fd_sc_hd__clkbuf_2
X_12847_ _12875_/CLK line[42] vssd1 vssd1 vccd1 vccd1 _12848_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_206_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_DATA\[17\].CLKBUF\[4\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12778_ _12778_/A _12809_/Y vssd1 vssd1 vccd1 vccd1 _13618_/Z sky130_fd_sc_hd__ebufn_2
XPHY_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11729_ _11755_/CLK line[43] vssd1 vssd1 vccd1 vccd1 _11730_/A sky130_fd_sc_hd__dfxtp_1
XPHY_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05250_ _05280_/CLK line[16] vssd1 vssd1 vccd1 vccd1 _05251_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06691__D line[44] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05181_ _05181_/A _05214_/Y vssd1 vssd1 vccd1 vccd1 _13861_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_143_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[29\].VALID\[3\].FF OVHB\[29\].V/CLK A[10] vssd1 vssd1 vccd1 vccd1 OVHB\[29\].VALID\[3\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_08940_ _08940_/A _08959_/Y vssd1 vssd1 vccd1 vccd1 _13700_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_170_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_MUX.M\[2\].MUX\[3\]_A0 _13669_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[3\].VALID\[10\].TOBUF OVHB\[3\].VALID\[10\].FF/Q OVHB\[3\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04932_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__09507__D line[37] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08871_ _08885_/CLK line[2] vssd1 vssd1 vccd1 vccd1 _08872_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_97_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07822_ _07822_/A _07839_/Y vssd1 vssd1 vccd1 vccd1 _13702_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[30\].VALID\[6\].TOBUF OVHB\[30\].VALID\[6\].FF/Q OVHB\[30\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04923_/A2 sky130_fd_sc_hd__ebufn_2
XOVHB\[11\].VALID\[0\].FF OVHB\[11\].V/CLK A[7] vssd1 vssd1 vccd1 vccd1 OVHB\[11\].VALID\[0\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_OVHB\[26\].VALID\[7\].FF_D A[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07753_ _07765_/CLK line[3] vssd1 vssd1 vccd1 vccd1 _07754_/A sky130_fd_sc_hd__dfxtp_1
X_04965_ _04965_/CLK line[9] vssd1 vssd1 vccd1 vccd1 _04966_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11772__D line[63] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06704_ _06704_/A _06719_/Y vssd1 vssd1 vccd1 vccd1 _13704_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06866__D line[124] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07684_ _07684_/A _07699_/Y vssd1 vssd1 vccd1 vccd1 _13844_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09242__D line[58] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05770__D line[121] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09423_ _09445_/CLK line[13] vssd1 vssd1 vccd1 vccd1 _09424_/A sky130_fd_sc_hd__dfxtp_1
X_06635_ _06645_/CLK line[4] vssd1 vssd1 vccd1 vccd1 _06636_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10388__D line[56] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09354_ _09354_/A _09379_/Y vssd1 vssd1 vccd1 vccd1 _13834_/Z sky130_fd_sc_hd__ebufn_2
X_06566_ _06566_/A _06579_/Y vssd1 vssd1 vccd1 vccd1 _13846_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13699__D line[33] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08305_ _08325_/CLK line[14] vssd1 vssd1 vccd1 vccd1 _08306_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_21_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05517_ _05525_/CLK line[5] vssd1 vssd1 vccd1 vccd1 _05518_/A sky130_fd_sc_hd__dfxtp_1
X_09285_ _09305_/CLK line[78] vssd1 vssd1 vccd1 vccd1 _09286_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_166_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06497_ _06505_/CLK line[69] vssd1 vssd1 vccd1 vccd1 _06498_/A sky130_fd_sc_hd__dfxtp_1
X_08236_ _08236_/A _08259_/Y vssd1 vssd1 vccd1 vccd1 _13836_/Z sky130_fd_sc_hd__ebufn_2
X_05448_ _05448_/A _05459_/Y vssd1 vssd1 vccd1 vccd1 _13848_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_20_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08167_ _08185_/CLK line[79] vssd1 vssd1 vccd1 vccd1 _08168_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_134_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05379_ _05385_/CLK line[70] vssd1 vssd1 vccd1 vccd1 _05380_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_119_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11012__D line[85] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07118_ _07118_/A _07139_/Y vssd1 vssd1 vccd1 vccd1 _13838_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06106__D line[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08098_ _08098_/A _08119_/Y vssd1 vssd1 vccd1 vccd1 _13698_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11947__D line[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07049_ _07065_/CLK line[65] vssd1 vssd1 vccd1 vccd1 _07050_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_122_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05945__D line[73] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09417__D line[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06403__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08321__D line[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10060_ _10060_/A _10079_/Y vssd1 vssd1 vccd1 vccd1 _13700_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_47_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XOVHB\[27\].VALID\[5\].FF OVHB\[27\].V/CLK A[12] vssd1 vssd1 vccd1 vccd1 OVHB\[27\].VALID\[5\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_85_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10962_ _10962_/A _10989_/Y vssd1 vssd1 vccd1 vccd1 _13762_/Z sky130_fd_sc_hd__ebufn_2
X_13750_ _13750_/CLK line[57] vssd1 vssd1 vccd1 vccd1 _13751_/A sky130_fd_sc_hd__dfxtp_1
XOVHB\[6\].VALID\[11\].FF OVHB\[6\].V/CLK A[18] vssd1 vssd1 vccd1 vccd1 OVHB\[6\].VALID\[11\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__05680__D line[94] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12701_ _12701_/A _12704_/Y vssd1 vssd1 vccd1 vccd1 _13821_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__10298__D line[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13681_ _13681_/A _13684_/Y vssd1 vssd1 vccd1 vccd1 _13681_/Z sky130_fd_sc_hd__ebufn_2
X_10893_ _10915_/CLK line[45] vssd1 vssd1 vccd1 vccd1 _10894_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12632_ _12632_/CLK _12633_/X vssd1 vssd1 vccd1 vccd1 _12630_/CLK sky130_fd_sc_hd__dlclkp_1
XPHY_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12563_ _13936_/X wr vssd1 vssd1 vccd1 vccd1 _12563_/X sky130_fd_sc_hd__and2_1
XPHY_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_OVHB\[7\].VALID\[2\].FF_D A[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11514_ _13926_/X vssd1 vssd1 vccd1 vccd1 _11514_/Y sky130_fd_sc_hd__inv_2
XPHY_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12494_ _13935_/X vssd1 vssd1 vccd1 vccd1 _12494_/Y sky130_fd_sc_hd__inv_2
XPHY_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11445_ _11475_/CLK line[32] vssd1 vssd1 vccd1 vccd1 _11446_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_171_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XDATA\[0\].CLKBUF\[7\] clk vssd1 vssd1 vccd1 vccd1 _05212_/CLK sky130_fd_sc_hd__clkbuf_4
X_11376_ _11376_/A _11409_/Y vssd1 vssd1 vccd1 vccd1 _13616_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_98_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10761__D line[98] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13115_ _13115_/A _13124_/Y vssd1 vssd1 vccd1 vccd1 _13675_/Z sky130_fd_sc_hd__ebufn_2
X_10327_ _10355_/CLK line[42] vssd1 vssd1 vccd1 vccd1 _10328_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05855__D line[46] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08231__D line[108] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13046_ _13050_/CLK line[119] vssd1 vssd1 vccd1 vccd1 _13047_/A sky130_fd_sc_hd__dfxtp_1
X_10258_ _10258_/A _10289_/Y vssd1 vssd1 vccd1 vccd1 _13618_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_78_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10189_ _10215_/CLK line[107] vssd1 vssd1 vccd1 vccd1 _10190_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_93_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XOVHB\[26\].VALID\[12\].TOBUF OVHB\[26\].VALID\[12\].FF/Q OVHB\[26\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04929_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__12688__D line[83] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__04926__B1 A_h[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13948_ _13949_/A _13949_/B _13949_/C _13949_/D vssd1 vssd1 vccd1 vccd1 _13948_/X
+ sky130_fd_sc_hd__and4b_4
XFILLER_47_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13879_ _13879_/A _13894_/Y vssd1 vssd1 vccd1 vccd1 _13879_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09997__D line[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XDATA\[30\].CLKBUF\[5\] clk vssd1 vssd1 vccd1 vccd1 _11582_/CLK sky130_fd_sc_hd__clkbuf_4
XANTENNA__10001__D line[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06420_ _06420_/A _06439_/Y vssd1 vssd1 vccd1 vccd1 _13700_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_61_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XOVHB\[25\].VALID\[7\].FF OVHB\[25\].V/CLK A[14] vssd1 vssd1 vccd1 vccd1 OVHB\[25\].VALID\[7\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_22_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06351_ _06365_/CLK line[2] vssd1 vssd1 vccd1 vccd1 _06352_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10936__D line[50] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13312__D line[127] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05302_ _05302_/A _05319_/Y vssd1 vssd1 vccd1 vccd1 _13702_/Z sky130_fd_sc_hd__ebufn_2
X_09070_ _09070_/A _09099_/Y vssd1 vssd1 vccd1 vccd1 _13830_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_147_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08406__D line[60] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06282_ _06282_/A _06299_/Y vssd1 vssd1 vccd1 vccd1 _13842_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__07310__D line[57] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08021_ _08045_/CLK line[12] vssd1 vssd1 vccd1 vccd1 _08022_/A sky130_fd_sc_hd__dfxtp_1
X_05233_ _05245_/CLK line[3] vssd1 vssd1 vccd1 vccd1 _05234_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_116_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_DATA\[15\].CLKBUF\[6\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[6\].VALID\[4\].TOBUF OVHB\[6\].VALID\[4\].FF/Q OVHB\[6\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04925_/B2 sky130_fd_sc_hd__ebufn_2
XFILLER_115_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05164_ _05164_/A _05179_/Y vssd1 vssd1 vccd1 vccd1 _13844_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_116_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_MUX.SEL1BUF\[0\]_A A[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09972_ _09972_/CLK _09973_/X vssd1 vssd1 vccd1 vccd1 _09970_/CLK sky130_fd_sc_hd__dlclkp_1
X_05095_ _05105_/CLK line[68] vssd1 vssd1 vccd1 vccd1 _05096_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_170_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08923_ _13915_/X wr vssd1 vssd1 vccd1 vccd1 _08923_/X sky130_fd_sc_hd__and2_1
X_08854_ _13914_/X vssd1 vssd1 vccd1 vccd1 _08854_/Y sky130_fd_sc_hd__inv_2
XANTENNA__07980__D line[112] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07805_ _07835_/CLK line[32] vssd1 vssd1 vccd1 vccd1 _07806_/A sky130_fd_sc_hd__dfxtp_1
X_08785_ _08815_/CLK line[96] vssd1 vssd1 vccd1 vccd1 _08786_/A sky130_fd_sc_hd__dfxtp_1
X_05997_ _06015_/CLK line[111] vssd1 vssd1 vccd1 vccd1 _05998_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_55_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07736_ _07736_/A _07769_/Y vssd1 vssd1 vccd1 vccd1 _13616_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__06596__D line[114] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_04948_ _04948_/A _04969_/Y vssd1 vssd1 vccd1 vccd1 _13628_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA_DATA\[8\].CLKBUF\[6\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07667_ _07695_/CLK line[106] vssd1 vssd1 vccd1 vccd1 _07668_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06893__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09406_ _09410_/CLK line[119] vssd1 vssd1 vccd1 vccd1 _09407_/A sky130_fd_sc_hd__dfxtp_1
X_06618_ _06618_/A _06649_/Y vssd1 vssd1 vccd1 vccd1 _13618_/Z sky130_fd_sc_hd__ebufn_2
X_07598_ _07598_/A _07629_/Y vssd1 vssd1 vccd1 vccd1 _13758_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_71_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05005__D line[32] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09337_ _09337_/A _09344_/Y vssd1 vssd1 vccd1 vccd1 _13817_/Z sky130_fd_sc_hd__ebufn_2
X_06549_ _06575_/CLK line[107] vssd1 vssd1 vccd1 vccd1 _06550_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_187_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09268_ _09270_/CLK line[56] vssd1 vssd1 vccd1 vccd1 _09269_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07220__D line[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08219_ _08219_/A _08224_/Y vssd1 vssd1 vccd1 vccd1 _13819_/Z sky130_fd_sc_hd__ebufn_2
X_09199_ _09199_/A _09204_/Y vssd1 vssd1 vccd1 vccd1 _13679_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_193_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XOVHB\[23\].VALID\[9\].FF OVHB\[23\].V/CLK A[16] vssd1 vssd1 vccd1 vccd1 OVHB\[23\].VALID\[9\].FF/Q
+ sky130_fd_sc_hd__dfxtp_1
X_11230_ _11230_/CLK line[57] vssd1 vssd1 vccd1 vccd1 _11231_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_20_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11677__D line[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11161_ _11161_/A _11164_/Y vssd1 vssd1 vccd1 vccd1 _13681_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__09147__D line[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10112_ _10112_/CLK _10113_/X vssd1 vssd1 vccd1 vccd1 _10110_/CLK sky130_fd_sc_hd__dlclkp_1
X_11092_ _11092_/CLK _11093_/X vssd1 vssd1 vccd1 vccd1 _11090_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_88_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10043_ _13922_/X wr vssd1 vssd1 vccd1 vccd1 _10043_/X sky130_fd_sc_hd__and2_1
XFILLER_0_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08986__D line[55] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12301__D line[34] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13802_ _13820_/CLK line[95] vssd1 vssd1 vccd1 vccd1 _13803_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_152_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11994_ _12000_/CLK line[22] vssd1 vssd1 vccd1 vccd1 _11995_/A sky130_fd_sc_hd__dfxtp_1
X_13733_ _13733_/A _13754_/Y vssd1 vssd1 vccd1 vccd1 _13733_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_189_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10945_ _10945_/A _10954_/Y vssd1 vssd1 vccd1 vccd1 _13745_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_45_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13664_ _13680_/CLK line[17] vssd1 vssd1 vccd1 vccd1 _13665_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09610__D line[84] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10876_ _10880_/CLK line[23] vssd1 vssd1 vccd1 vccd1 _10877_/A sky130_fd_sc_hd__dfxtp_1
X_12615_ _12615_/A _12634_/Y vssd1 vssd1 vccd1 vccd1 _13735_/Z sky130_fd_sc_hd__ebufn_2
XPHY_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13595_ _13595_/A _13614_/Y vssd1 vssd1 vccd1 vccd1 _13875_/Z sky130_fd_sc_hd__ebufn_2
XPHY_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12546_ _12560_/CLK line[18] vssd1 vssd1 vccd1 vccd1 _12547_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_12_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12477_ _12477_/A _12494_/Y vssd1 vssd1 vccd1 vccd1 _13877_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_8_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11428_ _11440_/CLK line[19] vssd1 vssd1 vccd1 vccd1 _11429_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11587__D line[106] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10491__D line[103] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11359_ _11359_/A _11374_/Y vssd1 vssd1 vccd1 vccd1 _13879_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_4_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05585__D line[36] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05920_ _05920_/A _05949_/Y vssd1 vssd1 vccd1 vccd1 _13760_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08896__D line[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_MUX.M\[2\].MUX\[0\]_A3 _13861_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13029_ _13029_/A _13054_/Y vssd1 vssd1 vccd1 vccd1 _13869_/Z sky130_fd_sc_hd__ebufn_2
X_05851_ _05875_/CLK line[44] vssd1 vssd1 vccd1 vccd1 _05852_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_66_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08570_ _08570_/CLK line[121] vssd1 vssd1 vccd1 vccd1 _08571_/A sky130_fd_sc_hd__dfxtp_1
X_05782_ _05782_/A _05809_/Y vssd1 vssd1 vccd1 vccd1 _13622_/Z sky130_fd_sc_hd__ebufn_2
X_07521_ _07521_/A _07524_/Y vssd1 vssd1 vccd1 vccd1 _13681_/Z sky130_fd_sc_hd__ebufn_2
XOVHB\[4\].VALID\[9\].TOBUF OVHB\[4\].VALID\[9\].FF/Q OVHB\[4\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04914_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA_OVHB\[2\].VALID\[11\].FF_D A[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XOVHB\[14\].VOBUF OVHB\[14\].V/Q OVHB\[14\].INV/Y vssd1 vssd1 vccd1 vccd1 _04912_/B1
+ sky130_fd_sc_hd__ebufn_2
XFILLER_34_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07452_ _07452_/CLK _07453_/X vssd1 vssd1 vccd1 vccd1 _07450_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_35_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09520__D line[48] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06403_ _13904_/X wr vssd1 vssd1 vccd1 vccd1 _06403_/X sky130_fd_sc_hd__and2_1
XFILLER_210_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10666__D line[55] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07383_ _13910_/X wr vssd1 vssd1 vccd1 vccd1 _07383_/X sky130_fd_sc_hd__and2_1
XANTENNA__13042__D line[117] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_DATA\[29\].CLKBUF\[0\]_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09122_ _09130_/CLK line[117] vssd1 vssd1 vccd1 vccd1 _09123_/A sky130_fd_sc_hd__dfxtp_1
X_06334_ _13903_/X vssd1 vssd1 vccd1 vccd1 _06334_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08136__D line[50] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08714__A _13914_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09053_ _09053_/A _09064_/Y vssd1 vssd1 vccd1 vccd1 _13813_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_163_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06265_ _06295_/CLK line[96] vssd1 vssd1 vccd1 vccd1 _06266_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07975__D line[105] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08433__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08004_ _08010_/CLK line[118] vssd1 vssd1 vccd1 vccd1 _08005_/A sky130_fd_sc_hd__dfxtp_1
X_05216_ _05216_/A _05249_/Y vssd1 vssd1 vccd1 vccd1 _13616_/Z sky130_fd_sc_hd__ebufn_2
X_06196_ _06196_/A _06229_/Y vssd1 vssd1 vccd1 vccd1 _13756_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_131_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05147_ _05175_/CLK line[106] vssd1 vssd1 vccd1 vccd1 _05148_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__05495__D line[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09955_ _09955_/A _09974_/Y vssd1 vssd1 vccd1 vccd1 _13875_/Z sky130_fd_sc_hd__ebufn_2
X_05078_ _05078_/A _05109_/Y vssd1 vssd1 vccd1 vccd1 _13758_/Z sky130_fd_sc_hd__ebufn_2
X_08906_ _08920_/CLK line[18] vssd1 vssd1 vccd1 vccd1 _08907_/A sky130_fd_sc_hd__dfxtp_1
X_09886_ _09900_/CLK line[82] vssd1 vssd1 vccd1 vccd1 _09887_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08837_ _08837_/A _08854_/Y vssd1 vssd1 vccd1 vccd1 _13877_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__13217__D line[69] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08768_ _08780_/CLK line[83] vssd1 vssd1 vccd1 vccd1 _08769_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_82_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07719_ _07719_/A _07734_/Y vssd1 vssd1 vccd1 vccd1 _13879_/Z sky130_fd_sc_hd__ebufn_2
X_08699_ _08699_/A _08714_/Y vssd1 vssd1 vccd1 vccd1 _13739_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__08608__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10730_ _10740_/CLK line[84] vssd1 vssd1 vccd1 vccd1 _10731_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_25_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_OVHB\[3\].VALID\[5\].FF_D A[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10576__D line[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10661_ _10661_/A _10674_/Y vssd1 vssd1 vccd1 vccd1 _13741_/Z sky130_fd_sc_hd__ebufn_2
X_12400_ _12420_/CLK line[94] vssd1 vssd1 vccd1 vccd1 _12401_/A sky130_fd_sc_hd__dfxtp_1
X_13380_ _13400_/CLK line[30] vssd1 vssd1 vccd1 vccd1 _13381_/A sky130_fd_sc_hd__dfxtp_1
X_10592_ _10600_/CLK line[21] vssd1 vssd1 vccd1 vccd1 _10593_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12791__D line[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12331_ _12331_/A _12354_/Y vssd1 vssd1 vccd1 vccd1 _13731_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_126_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XOVHB\[11\].VALID\[4\].TOBUF OVHB\[11\].VALID\[4\].FF/Q OVHB\[11\].INV/Y vssd1 vssd1
+ vccd1 vccd1 _04925_/B2 sky130_fd_sc_hd__ebufn_2
XANTENNA__07885__D line[78] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12262_ _12280_/CLK line[31] vssd1 vssd1 vccd1 vccd1 _12263_/A sky130_fd_sc_hd__dfxtp_1
X_11213_ _11213_/A _11234_/Y vssd1 vssd1 vccd1 vccd1 _13733_/Z sky130_fd_sc_hd__ebufn_2
X_12193_ _12193_/A _12214_/Y vssd1 vssd1 vccd1 vccd1 _13873_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__11200__D line[48] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05983__A _13902_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11144_ _11160_/CLK line[17] vssd1 vssd1 vccd1 vccd1 _11145_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11075_ _11075_/A _11094_/Y vssd1 vssd1 vccd1 vccd1 _13875_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_0_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10026_ _10040_/CLK line[18] vssd1 vssd1 vccd1 vccd1 _10027_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_48_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10113__B wr vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13127__D line[42] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12031__D line[39] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07125__D line[100] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12966__D line[82] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11977_ _11977_/A _12004_/Y vssd1 vssd1 vccd1 vccd1 _13657_/Z sky130_fd_sc_hd__ebufn_2
X_13716_ _13716_/A _13719_/Y vssd1 vssd1 vccd1 vccd1 _13716_/Z sky130_fd_sc_hd__ebufn_2
XFILLER_189_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10928_ _10950_/CLK line[61] vssd1 vssd1 vccd1 vccd1 _10929_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_205_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09340__D line[89] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13647_ _13647_/CLK _13648_/X vssd1 vssd1 vccd1 vccd1 _13645_/CLK sky130_fd_sc_hd__dlclkp_1
XFILLER_177_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10859_ _10859_/A _10884_/Y vssd1 vssd1 vccd1 vccd1 _13659_/Z sky130_fd_sc_hd__ebufn_2
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13578_ _13898_/Y wr vssd1 vssd1 vccd1 vccd1 _13578_/X sky130_fd_sc_hd__and2_1
XFILLER_12_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_MUX.M\[3\].MUX\[5\]_A0 _13659_/Z vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12529_ _13936_/X vssd1 vssd1 vccd1 vccd1 _12529_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06050_ _06050_/CLK line[121] vssd1 vssd1 vccd1 vccd1 _06051_/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06054__A _13902_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_OVHB\[18\].VALID\[2\].FF_D A[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05001_ _05001_/A _05004_/Y vssd1 vssd1 vccd1 vccd1 _13681_/Z sky130_fd_sc_hd__ebufn_2
XANTENNA__12206__D line[119] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06952_ _06960_/CLK line[21] vssd1 vssd1 vccd1 vccd1 _06953_/A sky130_fd_sc_hd__dfxtp_1
X_09740_ _09760_/CLK line[30] vssd1 vssd1 vccd1 vccd1 _09741_/A sky130_fd_sc_hd__dfxtp_1
.ends

