VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO apb_sys_0
  CLASS BLOCK ;
  FOREIGN apb_sys_0 ;
  ORIGIN 0.000 0.000 ;
  SIZE 450.000 BY 700.000 ;
  PIN HADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 0.000 2.210 4.000 ;
    END
  END HADDR[0]
  PIN HADDR[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 0.000 45.910 4.000 ;
    END
  END HADDR[10]
  PIN HADDR[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.230 0.000 50.510 4.000 ;
    END
  END HADDR[11]
  PIN HADDR[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END HADDR[12]
  PIN HADDR[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 4.000 ;
    END
  END HADDR[13]
  PIN HADDR[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.570 0.000 63.850 4.000 ;
    END
  END HADDR[14]
  PIN HADDR[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END HADDR[15]
  PIN HADDR[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 0.000 72.590 4.000 ;
    END
  END HADDR[16]
  PIN HADDR[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.910 0.000 77.190 4.000 ;
    END
  END HADDR[17]
  PIN HADDR[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 0.000 81.330 4.000 ;
    END
  END HADDR[18]
  PIN HADDR[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 4.000 ;
    END
  END HADDR[19]
  PIN HADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 0.000 6.350 4.000 ;
    END
  END HADDR[1]
  PIN HADDR[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 0.000 90.070 4.000 ;
    END
  END HADDR[20]
  PIN HADDR[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 0.000 94.670 4.000 ;
    END
  END HADDR[21]
  PIN HADDR[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 0.000 98.810 4.000 ;
    END
  END HADDR[22]
  PIN HADDR[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END HADDR[23]
  PIN HADDR[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 0.000 108.010 4.000 ;
    END
  END HADDR[24]
  PIN HADDR[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 0.000 112.150 4.000 ;
    END
  END HADDR[25]
  PIN HADDR[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.470 0.000 116.750 4.000 ;
    END
  END HADDR[26]
  PIN HADDR[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 0.000 120.890 4.000 ;
    END
  END HADDR[27]
  PIN HADDR[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.210 0.000 125.490 4.000 ;
    END
  END HADDR[28]
  PIN HADDR[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 4.000 ;
    END
  END HADDR[29]
  PIN HADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.670 0.000 10.950 4.000 ;
    END
  END HADDR[2]
  PIN HADDR[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.950 0.000 134.230 4.000 ;
    END
  END HADDR[30]
  PIN HADDR[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END HADDR[31]
  PIN HADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 0.000 15.090 4.000 ;
    END
  END HADDR[3]
  PIN HADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END HADDR[4]
  PIN HADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 0.000 23.830 4.000 ;
    END
  END HADDR[5]
  PIN HADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 0.000 28.430 4.000 ;
    END
  END HADDR[6]
  PIN HADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.750 0.000 33.030 4.000 ;
    END
  END HADDR[7]
  PIN HADDR[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 4.000 ;
    END
  END HADDR[8]
  PIN HADDR[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.490 0.000 41.770 4.000 ;
    END
  END HADDR[9]
  PIN HCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 19.080 450.000 19.680 ;
    END
  END HCLK
  PIN HRDATA[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 4.000 ;
    END
  END HRDATA[0]
  PIN HRDATA[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END HRDATA[10]
  PIN HRDATA[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.450 0.000 191.730 4.000 ;
    END
  END HRDATA[11]
  PIN HRDATA[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.590 0.000 195.870 4.000 ;
    END
  END HRDATA[12]
  PIN HRDATA[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 0.000 200.470 4.000 ;
    END
  END HRDATA[13]
  PIN HRDATA[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.790 0.000 205.070 4.000 ;
    END
  END HRDATA[14]
  PIN HRDATA[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.930 0.000 209.210 4.000 ;
    END
  END HRDATA[15]
  PIN HRDATA[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.530 0.000 213.810 4.000 ;
    END
  END HRDATA[16]
  PIN HRDATA[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.670 0.000 217.950 4.000 ;
    END
  END HRDATA[17]
  PIN HRDATA[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 4.000 ;
    END
  END HRDATA[18]
  PIN HRDATA[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.870 0.000 227.150 4.000 ;
    END
  END HRDATA[19]
  PIN HRDATA[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 0.000 147.570 4.000 ;
    END
  END HRDATA[1]
  PIN HRDATA[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.010 0.000 231.290 4.000 ;
    END
  END HRDATA[20]
  PIN HRDATA[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.610 0.000 235.890 4.000 ;
    END
  END HRDATA[21]
  PIN HRDATA[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.750 0.000 240.030 4.000 ;
    END
  END HRDATA[22]
  PIN HRDATA[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.350 0.000 244.630 4.000 ;
    END
  END HRDATA[23]
  PIN HRDATA[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.490 0.000 248.770 4.000 ;
    END
  END HRDATA[24]
  PIN HRDATA[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.090 0.000 253.370 4.000 ;
    END
  END HRDATA[25]
  PIN HRDATA[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END HRDATA[26]
  PIN HRDATA[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.830 0.000 262.110 4.000 ;
    END
  END HRDATA[27]
  PIN HRDATA[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.430 0.000 266.710 4.000 ;
    END
  END HRDATA[28]
  PIN HRDATA[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 0.000 270.850 4.000 ;
    END
  END HRDATA[29]
  PIN HRDATA[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 0.000 152.170 4.000 ;
    END
  END HRDATA[2]
  PIN HRDATA[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.170 0.000 275.450 4.000 ;
    END
  END HRDATA[30]
  PIN HRDATA[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.770 0.000 280.050 4.000 ;
    END
  END HRDATA[31]
  PIN HRDATA[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.030 0.000 156.310 4.000 ;
    END
  END HRDATA[3]
  PIN HRDATA[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.630 0.000 160.910 4.000 ;
    END
  END HRDATA[4]
  PIN HRDATA[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.770 0.000 165.050 4.000 ;
    END
  END HRDATA[5]
  PIN HRDATA[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.370 0.000 169.650 4.000 ;
    END
  END HRDATA[6]
  PIN HRDATA[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.510 0.000 173.790 4.000 ;
    END
  END HRDATA[7]
  PIN HRDATA[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.110 0.000 178.390 4.000 ;
    END
  END HRDATA[8]
  PIN HRDATA[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.710 0.000 182.990 4.000 ;
    END
  END HRDATA[9]
  PIN HREADY
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.470 0.000 438.750 4.000 ;
    END
  END HREADY
  PIN HREADYOUT
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.210 0.000 447.490 4.000 ;
    END
  END HREADYOUT
  PIN HRESETn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 57.840 450.000 58.440 ;
    END
  END HRESETn
  PIN HSEL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.610 0.000 442.890 4.000 ;
    END
  END HSEL
  PIN HTRANS[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 0.000 425.410 4.000 ;
    END
  END HTRANS[0]
  PIN HTRANS[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.730 0.000 430.010 4.000 ;
    END
  END HTRANS[1]
  PIN HWDATA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.910 0.000 284.190 4.000 ;
    END
  END HWDATA[0]
  PIN HWDATA[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.070 0.000 328.350 4.000 ;
    END
  END HWDATA[10]
  PIN HWDATA[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.670 0.000 332.950 4.000 ;
    END
  END HWDATA[11]
  PIN HWDATA[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.810 0.000 337.090 4.000 ;
    END
  END HWDATA[12]
  PIN HWDATA[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 0.000 341.690 4.000 ;
    END
  END HWDATA[13]
  PIN HWDATA[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.550 0.000 345.830 4.000 ;
    END
  END HWDATA[14]
  PIN HWDATA[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.150 0.000 350.430 4.000 ;
    END
  END HWDATA[15]
  PIN HWDATA[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.750 0.000 355.030 4.000 ;
    END
  END HWDATA[16]
  PIN HWDATA[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.890 0.000 359.170 4.000 ;
    END
  END HWDATA[17]
  PIN HWDATA[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.490 0.000 363.770 4.000 ;
    END
  END HWDATA[18]
  PIN HWDATA[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.630 0.000 367.910 4.000 ;
    END
  END HWDATA[19]
  PIN HWDATA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.510 0.000 288.790 4.000 ;
    END
  END HWDATA[1]
  PIN HWDATA[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.230 0.000 372.510 4.000 ;
    END
  END HWDATA[20]
  PIN HWDATA[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 0.000 377.110 4.000 ;
    END
  END HWDATA[21]
  PIN HWDATA[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.970 0.000 381.250 4.000 ;
    END
  END HWDATA[22]
  PIN HWDATA[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.570 0.000 385.850 4.000 ;
    END
  END HWDATA[23]
  PIN HWDATA[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 0.000 389.990 4.000 ;
    END
  END HWDATA[24]
  PIN HWDATA[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.310 0.000 394.590 4.000 ;
    END
  END HWDATA[25]
  PIN HWDATA[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.450 0.000 398.730 4.000 ;
    END
  END HWDATA[26]
  PIN HWDATA[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.050 0.000 403.330 4.000 ;
    END
  END HWDATA[27]
  PIN HWDATA[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.650 0.000 407.930 4.000 ;
    END
  END HWDATA[28]
  PIN HWDATA[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.790 0.000 412.070 4.000 ;
    END
  END HWDATA[29]
  PIN HWDATA[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.650 0.000 292.930 4.000 ;
    END
  END HWDATA[2]
  PIN HWDATA[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.390 0.000 416.670 4.000 ;
    END
  END HWDATA[30]
  PIN HWDATA[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.530 0.000 420.810 4.000 ;
    END
  END HWDATA[31]
  PIN HWDATA[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.250 0.000 297.530 4.000 ;
    END
  END HWDATA[3]
  PIN HWDATA[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.850 0.000 302.130 4.000 ;
    END
  END HWDATA[4]
  PIN HWDATA[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 0.000 306.270 4.000 ;
    END
  END HWDATA[5]
  PIN HWDATA[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.590 0.000 310.870 4.000 ;
    END
  END HWDATA[6]
  PIN HWDATA[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.730 0.000 315.010 4.000 ;
    END
  END HWDATA[7]
  PIN HWDATA[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.330 0.000 319.610 4.000 ;
    END
  END HWDATA[8]
  PIN HWDATA[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.470 0.000 323.750 4.000 ;
    END
  END HWDATA[9]
  PIN HWRITE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.870 0.000 434.150 4.000 ;
    END
  END HWRITE
  PIN IRQ[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 96.600 450.000 97.200 ;
    END
  END IRQ[0]
  PIN IRQ[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 485.560 450.000 486.160 ;
    END
  END IRQ[10]
  PIN IRQ[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 524.320 450.000 524.920 ;
    END
  END IRQ[11]
  PIN IRQ[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 563.080 450.000 563.680 ;
    END
  END IRQ[12]
  PIN IRQ[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 601.840 450.000 602.440 ;
    END
  END IRQ[13]
  PIN IRQ[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 640.600 450.000 641.200 ;
    END
  END IRQ[14]
  PIN IRQ[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 679.360 450.000 679.960 ;
    END
  END IRQ[15]
  PIN IRQ[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 135.360 450.000 135.960 ;
    END
  END IRQ[1]
  PIN IRQ[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 174.120 450.000 174.720 ;
    END
  END IRQ[2]
  PIN IRQ[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 212.880 450.000 213.480 ;
    END
  END IRQ[3]
  PIN IRQ[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 252.320 450.000 252.920 ;
    END
  END IRQ[4]
  PIN IRQ[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 291.080 450.000 291.680 ;
    END
  END IRQ[5]
  PIN IRQ[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 329.840 450.000 330.440 ;
    END
  END IRQ[6]
  PIN IRQ[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 368.600 450.000 369.200 ;
    END
  END IRQ[7]
  PIN IRQ[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 407.360 450.000 407.960 ;
    END
  END IRQ[8]
  PIN IRQ[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 446.120 450.000 446.720 ;
    END
  END IRQ[9]
  PIN MSI_S2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 696.000 77.650 700.000 ;
    END
  END MSI_S2
  PIN MSI_S3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.370 696.000 146.650 700.000 ;
    END
  END MSI_S3
  PIN MSO_S2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 696.000 95.130 700.000 ;
    END
  END MSO_S2
  PIN MSO_S3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.850 696.000 164.130 700.000 ;
    END
  END MSO_S3
  PIN RsRx_S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 696.000 8.650 700.000 ;
    END
  END RsRx_S0
  PIN RsRx_S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 696.000 43.150 700.000 ;
    END
  END RsRx_S1
  PIN RsTx_S0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 696.000 25.670 700.000 ;
    END
  END RsTx_S0
  PIN RsTx_S1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 696.000 60.170 700.000 ;
    END
  END RsTx_S1
  PIN SCLK_S2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.350 696.000 129.630 700.000 ;
    END
  END SCLK_S2
  PIN SCLK_S3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.350 696.000 198.630 700.000 ;
    END
  END SCLK_S3
  PIN SSn_S2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 696.000 112.150 700.000 ;
    END
  END SSn_S2
  PIN SSn_S3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.330 696.000 181.610 700.000 ;
    END
  END SSn_S3
  PIN pwm_S6
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.290 696.000 423.570 700.000 ;
    END
  END pwm_S6
  PIN pwm_S7
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.770 696.000 441.050 700.000 ;
    END
  END pwm_S7
  PIN scl_i_S4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 696.000 216.110 700.000 ;
    END
  END scl_i_S4
  PIN scl_i_S5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.790 696.000 320.070 700.000 ;
    END
  END scl_i_S5
  PIN scl_o_S4
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.310 696.000 233.590 700.000 ;
    END
  END scl_o_S4
  PIN scl_o_S5
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.810 696.000 337.090 700.000 ;
    END
  END scl_o_S5
  PIN scl_oen_o_S4
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.330 696.000 250.610 700.000 ;
    END
  END scl_oen_o_S4
  PIN scl_oen_o_S5
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 696.000 354.570 700.000 ;
    END
  END scl_oen_o_S5
  PIN sda_i_S4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.810 696.000 268.090 700.000 ;
    END
  END sda_i_S4
  PIN sda_i_S5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.310 696.000 371.590 700.000 ;
    END
  END sda_i_S5
  PIN sda_o_S4
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.830 696.000 285.110 700.000 ;
    END
  END sda_o_S4
  PIN sda_o_S5
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.790 696.000 389.070 700.000 ;
    END
  END sda_o_S5
  PIN sda_oen_o_S4
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.310 696.000 302.590 700.000 ;
    END
  END sda_oen_o_S4
  PIN sda_oen_o_S5
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.270 696.000 406.550 700.000 ;
    END
  END sda_oen_o_S5
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 688.400 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 688.400 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 688.400 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 688.400 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 688.400 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 688.400 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 8.245 445.135 688.245 ;
      LAYER met1 ;
        RECT 1.910 6.840 447.510 688.400 ;
      LAYER met2 ;
        RECT 1.940 695.720 8.090 696.000 ;
        RECT 8.930 695.720 25.110 696.000 ;
        RECT 25.950 695.720 42.590 696.000 ;
        RECT 43.430 695.720 59.610 696.000 ;
        RECT 60.450 695.720 77.090 696.000 ;
        RECT 77.930 695.720 94.570 696.000 ;
        RECT 95.410 695.720 111.590 696.000 ;
        RECT 112.430 695.720 129.070 696.000 ;
        RECT 129.910 695.720 146.090 696.000 ;
        RECT 146.930 695.720 163.570 696.000 ;
        RECT 164.410 695.720 181.050 696.000 ;
        RECT 181.890 695.720 198.070 696.000 ;
        RECT 198.910 695.720 215.550 696.000 ;
        RECT 216.390 695.720 233.030 696.000 ;
        RECT 233.870 695.720 250.050 696.000 ;
        RECT 250.890 695.720 267.530 696.000 ;
        RECT 268.370 695.720 284.550 696.000 ;
        RECT 285.390 695.720 302.030 696.000 ;
        RECT 302.870 695.720 319.510 696.000 ;
        RECT 320.350 695.720 336.530 696.000 ;
        RECT 337.370 695.720 354.010 696.000 ;
        RECT 354.850 695.720 371.030 696.000 ;
        RECT 371.870 695.720 388.510 696.000 ;
        RECT 389.350 695.720 405.990 696.000 ;
        RECT 406.830 695.720 423.010 696.000 ;
        RECT 423.850 695.720 440.490 696.000 ;
        RECT 441.330 695.720 447.480 696.000 ;
        RECT 1.940 4.280 447.480 695.720 ;
        RECT 2.490 4.000 5.790 4.280 ;
        RECT 6.630 4.000 10.390 4.280 ;
        RECT 11.230 4.000 14.530 4.280 ;
        RECT 15.370 4.000 19.130 4.280 ;
        RECT 19.970 4.000 23.270 4.280 ;
        RECT 24.110 4.000 27.870 4.280 ;
        RECT 28.710 4.000 32.470 4.280 ;
        RECT 33.310 4.000 36.610 4.280 ;
        RECT 37.450 4.000 41.210 4.280 ;
        RECT 42.050 4.000 45.350 4.280 ;
        RECT 46.190 4.000 49.950 4.280 ;
        RECT 50.790 4.000 54.550 4.280 ;
        RECT 55.390 4.000 58.690 4.280 ;
        RECT 59.530 4.000 63.290 4.280 ;
        RECT 64.130 4.000 67.430 4.280 ;
        RECT 68.270 4.000 72.030 4.280 ;
        RECT 72.870 4.000 76.630 4.280 ;
        RECT 77.470 4.000 80.770 4.280 ;
        RECT 81.610 4.000 85.370 4.280 ;
        RECT 86.210 4.000 89.510 4.280 ;
        RECT 90.350 4.000 94.110 4.280 ;
        RECT 94.950 4.000 98.250 4.280 ;
        RECT 99.090 4.000 102.850 4.280 ;
        RECT 103.690 4.000 107.450 4.280 ;
        RECT 108.290 4.000 111.590 4.280 ;
        RECT 112.430 4.000 116.190 4.280 ;
        RECT 117.030 4.000 120.330 4.280 ;
        RECT 121.170 4.000 124.930 4.280 ;
        RECT 125.770 4.000 129.530 4.280 ;
        RECT 130.370 4.000 133.670 4.280 ;
        RECT 134.510 4.000 138.270 4.280 ;
        RECT 139.110 4.000 142.410 4.280 ;
        RECT 143.250 4.000 147.010 4.280 ;
        RECT 147.850 4.000 151.610 4.280 ;
        RECT 152.450 4.000 155.750 4.280 ;
        RECT 156.590 4.000 160.350 4.280 ;
        RECT 161.190 4.000 164.490 4.280 ;
        RECT 165.330 4.000 169.090 4.280 ;
        RECT 169.930 4.000 173.230 4.280 ;
        RECT 174.070 4.000 177.830 4.280 ;
        RECT 178.670 4.000 182.430 4.280 ;
        RECT 183.270 4.000 186.570 4.280 ;
        RECT 187.410 4.000 191.170 4.280 ;
        RECT 192.010 4.000 195.310 4.280 ;
        RECT 196.150 4.000 199.910 4.280 ;
        RECT 200.750 4.000 204.510 4.280 ;
        RECT 205.350 4.000 208.650 4.280 ;
        RECT 209.490 4.000 213.250 4.280 ;
        RECT 214.090 4.000 217.390 4.280 ;
        RECT 218.230 4.000 221.990 4.280 ;
        RECT 222.830 4.000 226.590 4.280 ;
        RECT 227.430 4.000 230.730 4.280 ;
        RECT 231.570 4.000 235.330 4.280 ;
        RECT 236.170 4.000 239.470 4.280 ;
        RECT 240.310 4.000 244.070 4.280 ;
        RECT 244.910 4.000 248.210 4.280 ;
        RECT 249.050 4.000 252.810 4.280 ;
        RECT 253.650 4.000 257.410 4.280 ;
        RECT 258.250 4.000 261.550 4.280 ;
        RECT 262.390 4.000 266.150 4.280 ;
        RECT 266.990 4.000 270.290 4.280 ;
        RECT 271.130 4.000 274.890 4.280 ;
        RECT 275.730 4.000 279.490 4.280 ;
        RECT 280.330 4.000 283.630 4.280 ;
        RECT 284.470 4.000 288.230 4.280 ;
        RECT 289.070 4.000 292.370 4.280 ;
        RECT 293.210 4.000 296.970 4.280 ;
        RECT 297.810 4.000 301.570 4.280 ;
        RECT 302.410 4.000 305.710 4.280 ;
        RECT 306.550 4.000 310.310 4.280 ;
        RECT 311.150 4.000 314.450 4.280 ;
        RECT 315.290 4.000 319.050 4.280 ;
        RECT 319.890 4.000 323.190 4.280 ;
        RECT 324.030 4.000 327.790 4.280 ;
        RECT 328.630 4.000 332.390 4.280 ;
        RECT 333.230 4.000 336.530 4.280 ;
        RECT 337.370 4.000 341.130 4.280 ;
        RECT 341.970 4.000 345.270 4.280 ;
        RECT 346.110 4.000 349.870 4.280 ;
        RECT 350.710 4.000 354.470 4.280 ;
        RECT 355.310 4.000 358.610 4.280 ;
        RECT 359.450 4.000 363.210 4.280 ;
        RECT 364.050 4.000 367.350 4.280 ;
        RECT 368.190 4.000 371.950 4.280 ;
        RECT 372.790 4.000 376.550 4.280 ;
        RECT 377.390 4.000 380.690 4.280 ;
        RECT 381.530 4.000 385.290 4.280 ;
        RECT 386.130 4.000 389.430 4.280 ;
        RECT 390.270 4.000 394.030 4.280 ;
        RECT 394.870 4.000 398.170 4.280 ;
        RECT 399.010 4.000 402.770 4.280 ;
        RECT 403.610 4.000 407.370 4.280 ;
        RECT 408.210 4.000 411.510 4.280 ;
        RECT 412.350 4.000 416.110 4.280 ;
        RECT 416.950 4.000 420.250 4.280 ;
        RECT 421.090 4.000 424.850 4.280 ;
        RECT 425.690 4.000 429.450 4.280 ;
        RECT 430.290 4.000 433.590 4.280 ;
        RECT 434.430 4.000 438.190 4.280 ;
        RECT 439.030 4.000 442.330 4.280 ;
        RECT 443.170 4.000 446.930 4.280 ;
      LAYER met3 ;
        RECT 18.465 680.360 446.000 688.325 ;
        RECT 18.465 678.960 445.600 680.360 ;
        RECT 18.465 641.600 446.000 678.960 ;
        RECT 18.465 640.200 445.600 641.600 ;
        RECT 18.465 602.840 446.000 640.200 ;
        RECT 18.465 601.440 445.600 602.840 ;
        RECT 18.465 564.080 446.000 601.440 ;
        RECT 18.465 562.680 445.600 564.080 ;
        RECT 18.465 525.320 446.000 562.680 ;
        RECT 18.465 523.920 445.600 525.320 ;
        RECT 18.465 486.560 446.000 523.920 ;
        RECT 18.465 485.160 445.600 486.560 ;
        RECT 18.465 447.120 446.000 485.160 ;
        RECT 18.465 445.720 445.600 447.120 ;
        RECT 18.465 408.360 446.000 445.720 ;
        RECT 18.465 406.960 445.600 408.360 ;
        RECT 18.465 369.600 446.000 406.960 ;
        RECT 18.465 368.200 445.600 369.600 ;
        RECT 18.465 330.840 446.000 368.200 ;
        RECT 18.465 329.440 445.600 330.840 ;
        RECT 18.465 292.080 446.000 329.440 ;
        RECT 18.465 290.680 445.600 292.080 ;
        RECT 18.465 253.320 446.000 290.680 ;
        RECT 18.465 251.920 445.600 253.320 ;
        RECT 18.465 213.880 446.000 251.920 ;
        RECT 18.465 212.480 445.600 213.880 ;
        RECT 18.465 175.120 446.000 212.480 ;
        RECT 18.465 173.720 445.600 175.120 ;
        RECT 18.465 136.360 446.000 173.720 ;
        RECT 18.465 134.960 445.600 136.360 ;
        RECT 18.465 97.600 446.000 134.960 ;
        RECT 18.465 96.200 445.600 97.600 ;
        RECT 18.465 58.840 446.000 96.200 ;
        RECT 18.465 57.440 445.600 58.840 ;
        RECT 18.465 20.080 446.000 57.440 ;
        RECT 18.465 18.680 445.600 20.080 ;
        RECT 18.465 10.715 446.000 18.680 ;
      LAYER met4 ;
        RECT 37.095 12.415 97.440 686.625 ;
        RECT 99.840 12.415 174.240 686.625 ;
        RECT 176.640 12.415 251.040 686.625 ;
        RECT 253.440 12.415 327.840 686.625 ;
        RECT 330.240 12.415 404.640 686.625 ;
        RECT 407.040 12.415 415.545 686.625 ;
  END
END apb_sys_0
END LIBRARY

