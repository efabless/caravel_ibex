* NGSPICE file created from apb_sys_0.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd1_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_16 abstract view
.subckt sky130_fd_sc_hd__clkinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_16 abstract view
.subckt sky130_fd_sc_hd__inv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_2 abstract view
.subckt sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

.subckt apb_sys_0 HADDR[0] HADDR[10] HADDR[11] HADDR[12] HADDR[13] HADDR[14] HADDR[15]
+ HADDR[16] HADDR[17] HADDR[18] HADDR[19] HADDR[1] HADDR[20] HADDR[21] HADDR[22] HADDR[23]
+ HADDR[24] HADDR[25] HADDR[26] HADDR[27] HADDR[28] HADDR[29] HADDR[2] HADDR[30] HADDR[31]
+ HADDR[3] HADDR[4] HADDR[5] HADDR[6] HADDR[7] HADDR[8] HADDR[9] HCLK HRDATA[0] HRDATA[10]
+ HRDATA[11] HRDATA[12] HRDATA[13] HRDATA[14] HRDATA[15] HRDATA[16] HRDATA[17] HRDATA[18]
+ HRDATA[19] HRDATA[1] HRDATA[20] HRDATA[21] HRDATA[22] HRDATA[23] HRDATA[24] HRDATA[25]
+ HRDATA[26] HRDATA[27] HRDATA[28] HRDATA[29] HRDATA[2] HRDATA[30] HRDATA[31] HRDATA[3]
+ HRDATA[4] HRDATA[5] HRDATA[6] HRDATA[7] HRDATA[8] HRDATA[9] HREADY HREADYOUT HRESETn
+ HSEL HTRANS[0] HTRANS[1] HWDATA[0] HWDATA[10] HWDATA[11] HWDATA[12] HWDATA[13] HWDATA[14]
+ HWDATA[15] HWDATA[16] HWDATA[17] HWDATA[18] HWDATA[19] HWDATA[1] HWDATA[20] HWDATA[21]
+ HWDATA[22] HWDATA[23] HWDATA[24] HWDATA[25] HWDATA[26] HWDATA[27] HWDATA[28] HWDATA[29]
+ HWDATA[2] HWDATA[30] HWDATA[31] HWDATA[3] HWDATA[4] HWDATA[5] HWDATA[6] HWDATA[7]
+ HWDATA[8] HWDATA[9] HWRITE IRQ[0] IRQ[10] IRQ[11] IRQ[12] IRQ[13] IRQ[14] IRQ[15]
+ IRQ[1] IRQ[2] IRQ[3] IRQ[4] IRQ[5] IRQ[6] IRQ[7] IRQ[8] IRQ[9] MSI_S2 MSI_S3 MSO_S2
+ MSO_S3 RsRx_S0 RsRx_S1 RsTx_S0 RsTx_S1 SCLK_S2 SCLK_S3 SSn_S2 SSn_S3 pwm_S6 pwm_S7
+ scl_i_S4 scl_i_S5 scl_o_S4 scl_o_S5 scl_oen_o_S4 scl_oen_o_S5 sda_i_S4 sda_i_S5
+ sda_o_S4 sda_o_S5 sda_oen_o_S4 sda_oen_o_S5 vccd1 vssd1
XANTENNA__21280__CLK _21342_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09671_ _21470_/Q _09657_/X _09670_/X _09660_/X vssd1 vssd1 vccd1 vccd1 _21470_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_55_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18869_ _18868_/X _10985_/Y _18929_/S vssd1 vssd1 vccd1 vccd1 _18869_/X sky130_fd_sc_hd__mux2_1
XFILLER_227_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20900_ _21147_/CLK _20900_/D repeater212/X vssd1 vssd1 vccd1 vccd1 _20900_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_199_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20831_ _21372_/CLK _20831_/D repeater269/X vssd1 vssd1 vccd1 vccd1 _20831_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_242_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18617__S _18617_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20762_ _21342_/CLK _20762_/D repeater211/X vssd1 vssd1 vccd1 vccd1 _20762_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20693_ _20693_/CLK _20693_/D repeater196/X vssd1 vssd1 vccd1 vccd1 _20693_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10974__A _20890_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14446__A _20028_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20762__RESET_B repeater211/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13791__B1 _20614_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18352__S _18875_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21314_ _21321_/CLK _21314_/D repeater222/X vssd1 vssd1 vccd1 vccd1 _21314_/Q sky130_fd_sc_hd__dfrtp_1
X_21245_ _21431_/CLK _21245_/D repeater238/X vssd1 vssd1 vccd1 vccd1 _21245_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_104_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21176_ _21183_/CLK _21176_/D repeater216/X vssd1 vssd1 vccd1 vccd1 _21176_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_77_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20127_ _21273_/CLK _20127_/D repeater245/X vssd1 vssd1 vccd1 vccd1 _20127_/Q sky130_fd_sc_hd__dfrtp_1
X_09938_ _13188_/A _10859_/B _13188_/C vssd1 vssd1 vccd1 vccd1 _17231_/A sky130_fd_sc_hd__or3_4
XFILLER_219_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20058_ _20480_/CLK _20058_/D repeater281/X vssd1 vssd1 vccd1 vccd1 _20058_/Q sky130_fd_sc_hd__dfrtp_1
X_09869_ _18966_/X _09869_/B vssd1 vssd1 vccd1 vccd1 _09872_/A sky130_fd_sc_hd__or2_1
XFILLER_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11900_ _11900_/A _11900_/B vssd1 vssd1 vccd1 vccd1 _21018_/D sky130_fd_sc_hd__nor2_1
XPHY_4300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12880_ _20740_/Q _12874_/X _12879_/X _12876_/X vssd1 vssd1 vccd1 vccd1 _20740_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16796__B1 _16779_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater190 repeater233/X vssd1 vssd1 vccd1 vccd1 repeater190/X sky130_fd_sc_hd__buf_8
XPHY_4322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11831_ _11831_/A vssd1 vssd1 vccd1 vccd1 _21036_/D sky130_fd_sc_hd__inv_2
XPHY_4344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18527__S _18907_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19945__RESET_B repeater251/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14550_ _20135_/Q vssd1 vssd1 vccd1 vccd1 _15832_/A sky130_fd_sc_hd__buf_1
XANTENNA__21003__CLK _21009_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11762_ _11761_/A _19873_/Q _11761_/Y _11753_/C vssd1 vssd1 vccd1 vccd1 _11763_/B
+ sky130_fd_sc_hd__o22a_1
XPHY_3643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13501_ _20444_/Q _13499_/X _13429_/X _13500_/X vssd1 vssd1 vccd1 vccd1 _20444_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_187_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10713_ _21319_/Q _10711_/Y _10708_/B _10712_/X vssd1 vssd1 vccd1 vccd1 _21319_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14481_ _20230_/Q _14480_/Y _14472_/X _14374_/B vssd1 vssd1 vccd1 vccd1 _20230_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_3687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11693_ _21081_/Q _11689_/X _11571_/X _11690_/X vssd1 vssd1 vccd1 vccd1 _21081_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10884__A _12544_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15220__B1 _20474_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16220_ _19428_/Q _16216_/X _16113_/X _16218_/X vssd1 vssd1 vccd1 vccd1 _19428_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13432_ input39/X vssd1 vssd1 vccd1 vccd1 _13432_/X sky130_fd_sc_hd__clkbuf_2
X_10644_ _10685_/A vssd1 vssd1 vccd1 vccd1 _10677_/A sky130_fd_sc_hd__clkbuf_2
XPHY_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16151_ _16158_/A vssd1 vssd1 vccd1 vccd1 _16151_/X sky130_fd_sc_hd__buf_1
XFILLER_127_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10575_ _10575_/A _10722_/A _10575_/C vssd1 vssd1 vccd1 vccd1 _10576_/A sky130_fd_sc_hd__or3_1
X_13363_ _20511_/Q _13358_/X _13146_/X _13360_/X vssd1 vssd1 vccd1 vccd1 _20511_/D
+ sky130_fd_sc_hd__a22o_1
Xrebuffer7 _14950_/A vssd1 vssd1 vccd1 vccd1 rebuffer7/X sky130_fd_sc_hd__dlygate4sd1_1
XANTENNA__18262__S _18902_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15102_ _20460_/Q vssd1 vssd1 vccd1 vccd1 _15102_/Y sky130_fd_sc_hd__inv_2
X_12314_ _12314_/A _12372_/A vssd1 vssd1 vccd1 vccd1 _12315_/B sky130_fd_sc_hd__or2_2
XANTENNA__20432__RESET_B repeater235/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16082_ _16088_/A vssd1 vssd1 vccd1 vccd1 _16082_/X sky130_fd_sc_hd__buf_1
XFILLER_5_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13294_ _13294_/A vssd1 vssd1 vccd1 vccd1 _13294_/X sky130_fd_sc_hd__buf_1
XFILLER_181_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19910_ _21151_/CLK _19910_/D repeater223/X vssd1 vssd1 vccd1 vccd1 _19910_/Q sky130_fd_sc_hd__dfrtp_2
X_15033_ _20069_/Q vssd1 vssd1 vccd1 vccd1 _15083_/A sky130_fd_sc_hd__inv_2
X_12245_ _20939_/Q vssd1 vssd1 vccd1 vccd1 _12428_/A sky130_fd_sc_hd__inv_2
XFILLER_181_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19841_ _21193_/CLK _19841_/D repeater226/X vssd1 vssd1 vccd1 vccd1 _19841_/Q sky130_fd_sc_hd__dfrtp_1
X_12176_ _20361_/Q vssd1 vssd1 vccd1 vccd1 _12176_/Y sky130_fd_sc_hd__inv_2
XFILLER_111_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09616__C _12716_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19093__S _19870_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11127_ _11127_/A _11136_/A vssd1 vssd1 vccd1 vccd1 _11131_/B sky130_fd_sc_hd__nor2_1
X_16984_ _16984_/A vssd1 vssd1 vccd1 vccd1 _16984_/X sky130_fd_sc_hd__clkbuf_2
X_19772_ _19789_/CLK _19772_/D vssd1 vssd1 vccd1 vccd1 _19772_/Q sky130_fd_sc_hd__dfxtp_1
X_11058_ _11058_/A _11089_/A vssd1 vssd1 vccd1 vccd1 _11085_/A sky130_fd_sc_hd__or2_1
X_15935_ _15943_/A vssd1 vssd1 vccd1 vccd1 _15935_/X sky130_fd_sc_hd__buf_1
X_18723_ _18722_/X _13951_/Y _18849_/S vssd1 vssd1 vccd1 vccd1 _18723_/X sky130_fd_sc_hd__mux2_1
X_10009_ _17034_/A vssd1 vssd1 vccd1 vccd1 _10009_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18654_ _17079_/Y _12100_/Y _18908_/S vssd1 vssd1 vccd1 vccd1 _18654_/X sky130_fd_sc_hd__mux2_1
XFILLER_237_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15866_ _15875_/A vssd1 vssd1 vccd1 vccd1 _15877_/A sky130_fd_sc_hd__inv_2
XFILLER_64_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21220__RESET_B repeater235/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17605_ _11940_/A _17348_/A _11932_/X _17253_/Y _17604_/X vssd1 vssd1 vccd1 vccd1
+ _17605_/X sky130_fd_sc_hd__o221a_1
X_14817_ _20113_/Q _20114_/Q _14818_/S vssd1 vssd1 vccd1 vccd1 _20114_/D sky130_fd_sc_hd__mux2_1
X_18585_ _17079_/Y _15226_/Y _18908_/S vssd1 vssd1 vccd1 vccd1 _18585_/X sky130_fd_sc_hd__mux2_1
X_15797_ _15832_/C vssd1 vssd1 vccd1 vccd1 _16484_/B sky130_fd_sc_hd__buf_1
XANTENNA__18437__S _18841_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18528__A1 _21480_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_240_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17536_ _17536_/A vssd1 vssd1 vccd1 vccd1 _17777_/A sky130_fd_sc_hd__buf_1
XFILLER_205_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14748_ _14747_/A _14541_/A _15832_/A _14747_/Y vssd1 vssd1 vccd1 vccd1 _20135_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_189_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17736__C1 _17734_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17467_ _21189_/Q vssd1 vssd1 vccd1 vccd1 _17467_/Y sky130_fd_sc_hd__inv_2
XFILLER_220_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14679_ _14679_/A _14679_/B vssd1 vssd1 vccd1 vccd1 _14682_/A sky130_fd_sc_hd__or2_1
XFILLER_149_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16418_ _19325_/Q _16413_/X _16375_/X _16414_/X vssd1 vssd1 vccd1 vccd1 _19325_/D
+ sky130_fd_sc_hd__a22o_1
X_19206_ _19202_/X _19203_/X _19204_/X _19205_/X _21005_/Q _21006_/Q vssd1 vssd1 vccd1
+ vccd1 _19206_/X sky130_fd_sc_hd__mux4_2
X_17398_ _17575_/A vssd1 vssd1 vccd1 vccd1 _17398_/X sky130_fd_sc_hd__buf_1
XANTENNA__12576__A1 _20888_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19137_ _19680_/Q _19808_/Q _19800_/Q _19792_/Q _19285_/S0 _21017_/Q vssd1 vssd1
+ vccd1 vccd1 _19137_/X sky130_fd_sc_hd__mux4_2
X_16349_ _19364_/Q _16345_/X _16281_/X _16347_/X vssd1 vssd1 vccd1 vccd1 _19364_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_185_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18172__S _18644_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20173__RESET_B repeater248/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19068_ _16735_/X _21142_/Q _19908_/D vssd1 vssd1 vccd1 vccd1 _19068_/X sky130_fd_sc_hd__mux2_1
XFILLER_218_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20102__RESET_B repeater259/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18019_ _18019_/A vssd1 vssd1 vccd1 vccd1 _18019_/X sky130_fd_sc_hd__buf_1
XFILLER_105_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19693__CLK _19813_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18900__S _18910_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21030_ _21207_/CLK _21030_/D repeater242/X vssd1 vssd1 vccd1 vccd1 _21030_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_234_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09723_ _11112_/A _20145_/Q _21237_/Q _09719_/Y _09722_/X vssd1 vssd1 vccd1 vccd1
+ _09769_/A sky130_fd_sc_hd__o221a_1
X_09654_ input40/X vssd1 vssd1 vccd1 vccd1 _12860_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_242_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18347__S _18910_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18519__A1 _13923_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20814_ _21379_/CLK _20814_/D repeater212/X vssd1 vssd1 vccd1 vccd1 _20814_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_169_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20745_ _21319_/CLK _20745_/D repeater191/X vssd1 vssd1 vccd1 vccd1 _20745_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20676_ _21480_/CLK _20676_/D repeater208/X vssd1 vssd1 vccd1 vccd1 _20676_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10360_ _10360_/A _10360_/B _10360_/C _10360_/D vssd1 vssd1 vccd1 vccd1 _10361_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_109_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13516__B1 _13446_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10291_ _21375_/Q vssd1 vssd1 vccd1 vccd1 _10291_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18810__S _18880_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12030_ _12030_/A vssd1 vssd1 vccd1 vccd1 _12030_/X sky130_fd_sc_hd__buf_1
XFILLER_2_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21228_ _21235_/CLK _21228_/D repeater249/X vssd1 vssd1 vccd1 vccd1 _21228_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_88_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21159_ _21162_/CLK _21159_/D repeater227/X vssd1 vssd1 vccd1 vccd1 _21159_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_238_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13981_ _20318_/Q _13979_/Y _13894_/B _13979_/A _13980_/X vssd1 vssd1 vccd1 vccd1
+ _20318_/D sky130_fd_sc_hd__o221a_1
X_15720_ _19663_/Q _15716_/X _15703_/X _15717_/X vssd1 vssd1 vccd1 vccd1 _19663_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13255__A _17178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_219_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12932_ input45/X vssd1 vssd1 vccd1 vccd1 _12932_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_37_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15651_ _19695_/Q _15647_/X _15485_/X _15648_/X vssd1 vssd1 vccd1 vccd1 _19695_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_234_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12863_ _12863_/A vssd1 vssd1 vccd1 vccd1 _12863_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__18257__S _18897_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14602_ _14602_/A vssd1 vssd1 vccd1 vccd1 _14602_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15470__A _15479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11814_ _11814_/A _11824_/A vssd1 vssd1 vccd1 vccd1 _11822_/A sky130_fd_sc_hd__or2_1
X_18370_ _18369_/X _21364_/Q _18841_/S vssd1 vssd1 vccd1 vccd1 _18370_/X sky130_fd_sc_hd__mux2_1
XPHY_4174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15582_ _15785_/A vssd1 vssd1 vccd1 vccd1 _15582_/X sky130_fd_sc_hd__clkbuf_2
XPHY_4185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12794_ _20783_/Q _12791_/X _09659_/X _12792_/X vssd1 vssd1 vccd1 vccd1 _20783_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17321_ _18856_/X _17857_/A _18865_/X _17320_/X vssd1 vssd1 vccd1 vccd1 _17321_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20684__RESET_B repeater208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14533_ _14656_/A vssd1 vssd1 vccd1 vccd1 _14663_/A sky130_fd_sc_hd__buf_1
X_11745_ _19843_/Q vssd1 vssd1 vccd1 vccd1 _16502_/A sky130_fd_sc_hd__inv_2
XPHY_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18930__A1 _19276_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12007__B1 _20251_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17252_ _21214_/Q vssd1 vssd1 vccd1 vccd1 _17252_/Y sky130_fd_sc_hd__inv_2
XFILLER_230_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14464_ _20632_/Q _14464_/B vssd1 vssd1 vccd1 vccd1 _14464_/X sky130_fd_sc_hd__or2_1
XPHY_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11676_ _10894_/A _21088_/Q _11676_/S vssd1 vssd1 vccd1 vccd1 _21088_/D sky130_fd_sc_hd__mux2_1
XPHY_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16203_ _19435_/Q _16195_/X _16202_/X _16198_/X vssd1 vssd1 vccd1 vccd1 _19435_/D
+ sky130_fd_sc_hd__a22o_1
X_13415_ _20481_/Q _13410_/X _13223_/X _13411_/X vssd1 vssd1 vccd1 vccd1 _20481_/D
+ sky130_fd_sc_hd__a22o_1
X_10627_ _10540_/A _20741_/Q _10657_/A _20756_/Q vssd1 vssd1 vccd1 vccd1 _10627_/X
+ sky130_fd_sc_hd__o22a_1
X_17183_ _20738_/Q vssd1 vssd1 vccd1 vccd1 _17183_/Y sky130_fd_sc_hd__inv_2
X_14395_ _21479_/Q vssd1 vssd1 vccd1 vccd1 _14395_/Y sky130_fd_sc_hd__inv_2
XANTENNA_repeater244_A repeater245/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16134_ _19469_/Q _16130_/X _16131_/X _16133_/X vssd1 vssd1 vccd1 vccd1 _19469_/D
+ sky130_fd_sc_hd__a22o_1
X_13346_ _13352_/A vssd1 vssd1 vccd1 vccd1 _13346_/X sky130_fd_sc_hd__buf_1
XFILLER_182_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10558_ _21323_/Q vssd1 vssd1 vccd1 vccd1 _10652_/A sky130_fd_sc_hd__inv_2
XFILLER_115_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18005__B _18006_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16065_ _16071_/A vssd1 vssd1 vccd1 vccd1 _16072_/A sky130_fd_sc_hd__inv_2
XANTENNA__18720__S _18897_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13277_ input57/X vssd1 vssd1 vccd1 vccd1 _13277_/X sky130_fd_sc_hd__clkbuf_2
X_10489_ _21303_/Q _10484_/Y _10754_/A _20666_/Q _10488_/X vssd1 vssd1 vccd1 vccd1
+ _10496_/C sky130_fd_sc_hd__o221a_1
X_15016_ _20081_/Q _15015_/Y _15002_/B _14952_/X vssd1 vssd1 vccd1 vccd1 _20081_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__18446__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12228_ _12228_/A vssd1 vssd1 vccd1 vccd1 _12429_/A sky130_fd_sc_hd__buf_1
XFILLER_97_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__21472__RESET_B repeater204/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19824_ _19835_/CLK _19824_/D vssd1 vssd1 vccd1 vccd1 _19824_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12159_ _12159_/A _12159_/B _12156_/X _12158_/X vssd1 vssd1 vccd1 vccd1 _12205_/A
+ sky130_fd_sc_hd__or4bb_4
XFILLER_111_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19755_ _19765_/CLK _19755_/D vssd1 vssd1 vccd1 vccd1 _19755_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__19867__RESET_B repeater216/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16967_ _16984_/A vssd1 vssd1 vccd1 vccd1 _16967_/X sky130_fd_sc_hd__buf_1
XANTENNA__18749__A1 _20638_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18706_ _17685_/Y _19216_/X _18930_/S vssd1 vssd1 vccd1 vccd1 _18706_/X sky130_fd_sc_hd__mux2_1
X_15918_ _20127_/Q vssd1 vssd1 vccd1 vccd1 _16325_/B sky130_fd_sc_hd__buf_1
XFILLER_204_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16898_ _16915_/A vssd1 vssd1 vccd1 vccd1 _16898_/X sky130_fd_sc_hd__buf_1
X_19686_ _19811_/CLK _19686_/D vssd1 vssd1 vccd1 vccd1 _19686_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_224_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15849_ _15856_/A vssd1 vssd1 vccd1 vccd1 _15849_/X sky130_fd_sc_hd__buf_1
X_18637_ _18848_/A0 _14125_/Y _18902_/S vssd1 vssd1 vccd1 vccd1 _18637_/X sky130_fd_sc_hd__mux2_1
XANTENNA__18167__S _18891_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18568_ _18845_/A0 _10456_/Y _18896_/S vssd1 vssd1 vccd1 vccd1 _18568_/X sky130_fd_sc_hd__mux2_1
XFILLER_220_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17519_ _19618_/Q vssd1 vssd1 vccd1 vccd1 _17519_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18499_ _17079_/Y _12094_/Y _18908_/S vssd1 vssd1 vccd1 vccd1 _18499_/X sky130_fd_sc_hd__mux2_2
XFILLER_220_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20530_ _21366_/CLK _20530_/D repeater265/X vssd1 vssd1 vccd1 vccd1 _20530_/Q sky130_fd_sc_hd__dfrtp_4
X_20461_ _20495_/CLK _20461_/D repeater273/X vssd1 vssd1 vccd1 vccd1 _20461_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_192_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20392_ _20951_/CLK _20392_/D repeater272/X vssd1 vssd1 vccd1 vccd1 _20392_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_145_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18630__S _18910_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21013_ _21121_/CLK _21013_/D repeater238/X vssd1 vssd1 vccd1 vccd1 _21013_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_102_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_157_HCLK_A clkbuf_opt_1_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09706_ _21458_/Q vssd1 vssd1 vccd1 vccd1 _09783_/A sky130_fd_sc_hd__inv_2
XFILLER_244_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09637_ _21480_/Q _09632_/X _09636_/X _09634_/X vssd1 vssd1 vccd1 vccd1 _21480_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_56_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20566__CLK _20592_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12788__A1 _20787_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18805__S _18884_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19260__S1 _20131_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11530_ _21143_/Q _11527_/X _10884_/X _11529_/X vssd1 vssd1 vccd1 vccd1 _21143_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20728_ _21375_/CLK _20728_/D repeater257/X vssd1 vssd1 vccd1 vccd1 _20728_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11461_ _11480_/A vssd1 vssd1 vccd1 vccd1 _11461_/X sky130_fd_sc_hd__buf_1
XPHY_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20659_ _20661_/CLK _20659_/D repeater261/X vssd1 vssd1 vccd1 vccd1 _20659_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__18106__A hold9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13200_ _13215_/A vssd1 vssd1 vccd1 vccd1 _13200_/X sky130_fd_sc_hd__buf_1
X_10412_ _10412_/A vssd1 vssd1 vccd1 vccd1 _10412_/Y sky130_fd_sc_hd__inv_2
X_11392_ _11410_/B _11786_/A _16596_/A vssd1 vssd1 vccd1 vccd1 _11408_/A sky130_fd_sc_hd__or3_1
X_14180_ _20288_/Q _14179_/Y _14174_/X _14099_/B vssd1 vssd1 vccd1 vccd1 _20288_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_137_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13131_ _20619_/Q _13126_/X _12922_/X _13127_/X vssd1 vssd1 vccd1 vccd1 _20619_/D
+ sky130_fd_sc_hd__a22o_1
X_10343_ _20723_/Q vssd1 vssd1 vccd1 vccd1 _17982_/A sky130_fd_sc_hd__inv_2
XANTENNA__18540__S _18680_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input55_A HWDATA[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13062_ _20661_/Q _13060_/X _12996_/X _13061_/X vssd1 vssd1 vccd1 vccd1 _20661_/D
+ sky130_fd_sc_hd__a22o_1
X_10274_ _10274_/A _10394_/A vssd1 vssd1 vccd1 vccd1 _10275_/B sky130_fd_sc_hd__or2_2
XFILLER_79_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12013_ _19067_/X _12010_/X _20998_/Q _12012_/X vssd1 vssd1 vccd1 vccd1 _20998_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_3_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17870_ _18555_/X _17857_/X _18567_/X _17869_/X vssd1 vssd1 vccd1 vccd1 _17870_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_238_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16821_ _19936_/Q vssd1 vssd1 vccd1 vccd1 _16821_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19960__RESET_B repeater184/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16752_ _19918_/Q vssd1 vssd1 vccd1 vccd1 _16753_/B sky130_fd_sc_hd__inv_2
X_19540_ _21445_/CLK _19540_/D vssd1 vssd1 vccd1 vccd1 _19540_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13964_ _14070_/B vssd1 vssd1 vccd1 vccd1 _13987_/A sky130_fd_sc_hd__buf_1
XFILLER_246_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_16_HCLK_A clkbuf_4_3_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15703_ _15793_/A vssd1 vssd1 vccd1 vccd1 _15703_/X sky130_fd_sc_hd__buf_1
XANTENNA__18600__A0 _18848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20865__RESET_B repeater247/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12915_ _12924_/A vssd1 vssd1 vccd1 vccd1 _12915_/X sky130_fd_sc_hd__buf_1
X_16683_ _16683_/A vssd1 vssd1 vccd1 vccd1 _16684_/A sky130_fd_sc_hd__buf_1
XFILLER_206_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19471_ _19776_/CLK _19471_/D vssd1 vssd1 vccd1 vccd1 _19471_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_79_HCLK_A clkbuf_4_13_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13895_ _13895_/A vssd1 vssd1 vccd1 vccd1 _13896_/B sky130_fd_sc_hd__inv_2
XFILLER_206_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15634_ _19705_/Q _15632_/X _15585_/X _15633_/X vssd1 vssd1 vccd1 vccd1 _19705_/D
+ sky130_fd_sc_hd__a22o_1
X_18422_ _18421_/X _16800_/Y _18667_/S vssd1 vssd1 vccd1 vccd1 _18422_/X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_4_HCLK_A clkbuf_opt_2_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12846_ _20754_/Q _12841_/X _09638_/X _12842_/X vssd1 vssd1 vccd1 vccd1 _20754_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18353_ _18035_/Y _20797_/Q _18849_/S vssd1 vssd1 vccd1 vccd1 _18353_/X sky130_fd_sc_hd__mux2_1
X_15565_ _19740_/Q _15561_/X _15548_/X _15563_/X vssd1 vssd1 vccd1 vccd1 _19740_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12777_ _12777_/A vssd1 vssd1 vccd1 vccd1 _12777_/X sky130_fd_sc_hd__buf_1
XANTENNA__19251__S1 _20133_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18715__S _18841_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17304_ _20245_/Q vssd1 vssd1 vccd1 vccd1 _17304_/Y sky130_fd_sc_hd__inv_2
X_14516_ _20213_/Q _14520_/A _14513_/A _14453_/X vssd1 vssd1 vccd1 vccd1 _20213_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11728_ _11735_/A vssd1 vssd1 vccd1 vccd1 _11737_/A sky130_fd_sc_hd__inv_2
X_18284_ _18283_/X _10286_/A _18886_/S vssd1 vssd1 vccd1 vccd1 _18284_/X sky130_fd_sc_hd__mux2_1
X_15496_ _19772_/Q _15492_/X _15454_/X _15494_/X vssd1 vssd1 vccd1 vccd1 _19772_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_230_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13728__A0 _15766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17235_ _17235_/A _17235_/B _17235_/C _17235_/D vssd1 vssd1 vccd1 vccd1 _17235_/Y
+ sky130_fd_sc_hd__nand4_4
XPHY_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14447_ _21478_/Q _14462_/A _14384_/Y _20032_/Q vssd1 vssd1 vccd1 vccd1 _14447_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_174_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11659_ _19112_/X vssd1 vssd1 vccd1 vccd1 _11659_/Y sky130_fd_sc_hd__inv_2
XPHY_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17166_ _21186_/Q vssd1 vssd1 vccd1 vccd1 _17166_/Y sky130_fd_sc_hd__inv_2
XANTENNA__09638__A input45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14378_ _14378_/A _14378_/B vssd1 vssd1 vccd1 vccd1 _14379_/A sky130_fd_sc_hd__or2_1
X_16117_ _20328_/Q vssd1 vssd1 vccd1 vccd1 _16117_/X sky130_fd_sc_hd__clkbuf_2
X_13329_ _13329_/A _13657_/B vssd1 vssd1 vccd1 vccd1 _13357_/A sky130_fd_sc_hd__or2_2
XFILLER_115_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17097_ _19358_/Q vssd1 vssd1 vccd1 vccd1 _17097_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18450__S _18885_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16048_ _16297_/A _16107_/B _16465_/C vssd1 vssd1 vccd1 vccd1 _16056_/A sky130_fd_sc_hd__or3_4
XANTENNA__17890__B2 _17326_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12999__A input56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19807_ _20172_/CLK _19807_/D vssd1 vssd1 vccd1 vccd1 _19807_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17999_ _17925_/X _17999_/B _17999_/C vssd1 vssd1 vccd1 vccd1 _17999_/Y sky130_fd_sc_hd__nand3b_4
XFILLER_85_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19738_ _19765_/CLK _19738_/D vssd1 vssd1 vccd1 vccd1 _19738_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_226_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19669_ _19813_/CLK _19669_/D vssd1 vssd1 vccd1 vccd1 _19669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_198_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19242__S1 _21004_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18625__S _18667_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13719__A0 input73/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20513_ _20929_/CLK _20513_/D repeater267/X vssd1 vssd1 vccd1 vccd1 _20513_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_193_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20444_ _20476_/CLK _20444_/D repeater280/X vssd1 vssd1 vccd1 vccd1 _20444_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_162_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20375_ _20957_/CLK _20375_/D repeater186/X vssd1 vssd1 vccd1 vccd1 _20375_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18360__S _18666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15892__B1 _15891_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12702__A _12708_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10961_ _10956_/Y _21037_/Q _21207_/Q _11811_/A _10960_/X vssd1 vssd1 vccd1 vccd1
+ _10969_/C sky130_fd_sc_hd__o221a_1
XFILLER_43_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12700_ _20819_/Q _12693_/X _12699_/X _12694_/X vssd1 vssd1 vccd1 vccd1 _20819_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_55_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20276__RESET_B repeater262/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13680_ _13680_/A vssd1 vssd1 vccd1 vccd1 _13680_/X sky130_fd_sc_hd__buf_1
X_10892_ _10892_/A vssd1 vssd1 vccd1 vccd1 _10892_/X sky130_fd_sc_hd__buf_2
XFILLER_203_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12631_ _12637_/A vssd1 vssd1 vccd1 vccd1 _12631_/X sky130_fd_sc_hd__buf_1
XPHY_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18535__S _18666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19233__S1 _21004_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15350_ _15588_/A vssd1 vssd1 vccd1 vccd1 _15350_/X sky130_fd_sc_hd__clkbuf_2
XPHY_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12562_ _12562_/A vssd1 vssd1 vccd1 vccd1 _19984_/D sky130_fd_sc_hd__buf_1
XPHY_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14301_ _20122_/Q _14300_/Y _20122_/Q _14300_/Y vssd1 vssd1 vccd1 vccd1 _14324_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_8_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11513_ _11513_/A vssd1 vssd1 vccd1 vccd1 _21147_/D sky130_fd_sc_hd__inv_2
XPHY_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15281_ _20489_/Q vssd1 vssd1 vccd1 vccd1 _18030_/A sky130_fd_sc_hd__inv_2
XPHY_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12493_ _12493_/A vssd1 vssd1 vccd1 vccd1 _12496_/A sky130_fd_sc_hd__inv_2
XANTENNA__10892__A _10892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17020_ _17020_/A _17023_/B vssd1 vssd1 vccd1 vccd1 _20006_/D sky130_fd_sc_hd__nor2_1
XANTENNA__13186__A1 _12968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14232_ _19892_/Q _14232_/B vssd1 vssd1 vccd1 vccd1 _14233_/B sky130_fd_sc_hd__or2_1
XPHY_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11444_ _21156_/Q _11444_/B vssd1 vssd1 vccd1 vccd1 _11445_/B sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_161_HCLK clkbuf_opt_0_HCLK/A vssd1 vssd1 vccd1 vccd1 _19784_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__11197__B1 _10898_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14163_ _20536_/Q vssd1 vssd1 vccd1 vccd1 _14163_/Y sky130_fd_sc_hd__inv_2
X_11375_ _11375_/A _11375_/B vssd1 vssd1 vccd1 vccd1 _11376_/D sky130_fd_sc_hd__or2_1
XANTENNA__18270__S _18879_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17321__B1 _18865_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13114_ _13141_/A vssd1 vssd1 vccd1 vccd1 _13133_/A sky130_fd_sc_hd__buf_1
XANTENNA__19754__CLK _19765_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10326_ _20718_/Q vssd1 vssd1 vccd1 vccd1 _10326_/Y sky130_fd_sc_hd__inv_2
X_14094_ _14094_/A _14187_/A vssd1 vssd1 vccd1 vccd1 _14095_/B sky130_fd_sc_hd__or2_1
X_18971_ _16526_/Y _16491_/Y _18975_/S vssd1 vssd1 vccd1 vccd1 _18971_/X sky130_fd_sc_hd__mux2_1
XFILLER_106_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13045_ _20666_/Q _13040_/X _12884_/X _13041_/X vssd1 vssd1 vccd1 vccd1 _20666_/D
+ sky130_fd_sc_hd__a22o_1
X_17922_ _20413_/Q vssd1 vssd1 vccd1 vccd1 _17922_/Y sky130_fd_sc_hd__inv_2
X_10257_ _21346_/Q vssd1 vssd1 vccd1 vccd1 _10262_/A sky130_fd_sc_hd__inv_2
XANTENNA_repeater207_A repeater208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17853_ _17853_/A vssd1 vssd1 vccd1 vccd1 _17853_/X sky130_fd_sc_hd__buf_1
XFILLER_79_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10188_ _21395_/Q _10187_/Y _10183_/X _10157_/B vssd1 vssd1 vccd1 vccd1 _21395_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_121_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15635__B1 _15588_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16804_ _16801_/Y _16802_/X _16803_/X vssd1 vssd1 vccd1 vccd1 _16804_/X sky130_fd_sc_hd__o21a_1
X_17784_ _19840_/Q vssd1 vssd1 vccd1 vccd1 _17784_/Y sky130_fd_sc_hd__inv_2
X_14996_ _14960_/D _14866_/B _14994_/Y _14989_/X vssd1 vssd1 vccd1 vccd1 _20088_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_208_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_140_HCLK_A clkbuf_4_3_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19523_ _20327_/CLK _19523_/D vssd1 vssd1 vccd1 vccd1 _19523_/Q sky130_fd_sc_hd__dfxtp_1
X_16735_ _20997_/Q _12003_/B _12003_/X vssd1 vssd1 vccd1 vccd1 _16735_/X sky130_fd_sc_hd__a21bo_1
X_13947_ _13947_/A _13947_/B _13947_/C _13947_/D vssd1 vssd1 vccd1 vccd1 _13962_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_34_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16666_ _21154_/Q _11442_/B _11443_/B vssd1 vssd1 vccd1 vccd1 _16666_/X sky130_fd_sc_hd__a21bo_1
X_19454_ _21234_/CLK _19454_/D vssd1 vssd1 vccd1 vccd1 _19454_/Q sky130_fd_sc_hd__dfxtp_1
X_13878_ _14030_/A _13974_/A vssd1 vssd1 vccd1 vccd1 _13879_/B sky130_fd_sc_hd__or2_2
XFILLER_62_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18405_ _18404_/X _20573_/Q _18907_/S vssd1 vssd1 vccd1 vccd1 _18405_/X sky130_fd_sc_hd__mux2_1
X_15617_ _19714_/Q _15611_/X _15477_/X _15613_/X vssd1 vssd1 vccd1 vccd1 _19714_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13949__B1 _20648_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12829_ _12841_/A vssd1 vssd1 vccd1 vccd1 _12829_/X sky130_fd_sc_hd__buf_1
XFILLER_34_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16597_ _16597_/A _19875_/Q vssd1 vssd1 vccd1 vccd1 _17046_/B sky130_fd_sc_hd__or2_2
X_19385_ _21222_/CLK _19385_/D vssd1 vssd1 vccd1 vccd1 _19385_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18445__S _18875_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19224__S1 _21004_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18336_ _18845_/A0 _10484_/Y _18896_/S vssd1 vssd1 vccd1 vccd1 _18336_/X sky130_fd_sc_hd__mux2_1
X_15548_ _15661_/A vssd1 vssd1 vccd1 vccd1 _15548_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_91_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18267_ _18266_/X _14095_/A _18904_/S vssd1 vssd1 vccd1 vccd1 _18267_/X sky130_fd_sc_hd__mux2_2
X_15479_ _15479_/A vssd1 vssd1 vccd1 vccd1 _15479_/X sky130_fd_sc_hd__buf_1
X_17218_ _17581_/A vssd1 vssd1 vccd1 vccd1 _17857_/A sky130_fd_sc_hd__buf_1
X_18198_ _18848_/A0 _17958_/Y _18666_/S vssd1 vssd1 vccd1 vccd1 _18198_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20129__SET_B repeater249/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17149_ _17553_/A vssd1 vssd1 vccd1 vccd1 _17292_/A sky130_fd_sc_hd__buf_1
XANTENNA__18180__S _18903_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20160_ _21121_/CLK _20160_/D repeater237/X vssd1 vssd1 vccd1 vccd1 _20160_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_89_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09971_ _21421_/Q _09968_/X _09663_/X _09970_/X vssd1 vssd1 vccd1 vccd1 _21421_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_226_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20091_ _20496_/CLK _20091_/D repeater273/X vssd1 vssd1 vccd1 vccd1 _20091_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_58_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12152__A2 _20346_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19160__S0 _19285_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_42_HCLK clkbuf_4_11_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _21196_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_26_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20993_ _21338_/CLK _20993_/D repeater222/X vssd1 vssd1 vccd1 vccd1 _20993_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17918__A2 _17214_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11663__A1 _10892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_241_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_62_HCLK_A clkbuf_4_14_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18355__S _18902_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19215__S1 _21004_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13168__A1 _20602_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21476_ _21476_/CLK _21476_/D repeater204/X vssd1 vssd1 vccd1 vccd1 _21476_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20427_ _20428_/CLK _20427_/D repeater270/X vssd1 vssd1 vccd1 vccd1 _20427_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_119_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11160_ _13180_/A _13527_/A _13181_/C _11160_/D vssd1 vssd1 vccd1 vccd1 _16525_/C
+ sky130_fd_sc_hd__or4_4
X_20358_ _20972_/CLK _20358_/D repeater279/X vssd1 vssd1 vccd1 vccd1 _20358_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_136_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10111_ _10204_/A _20780_/Q _21383_/Q _10109_/Y _10110_/X vssd1 vssd1 vccd1 vccd1
+ _10112_/D sky130_fd_sc_hd__o221a_1
X_11091_ _11086_/B _11079_/X _11090_/Y _11082_/X _11058_/A vssd1 vssd1 vccd1 vccd1
+ _11092_/A sky130_fd_sc_hd__o32a_1
XANTENNA_clkbuf_4_2_0_HCLK_A clkbuf_4_3_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20289_ _20592_/CLK _20289_/D repeater261/X vssd1 vssd1 vccd1 vccd1 _20289_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_96_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18803__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17606__A1 _11940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10042_ _21383_/Q vssd1 vssd1 vccd1 vccd1 _10204_/A sky130_fd_sc_hd__inv_2
XFILLER_248_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17942__B _17943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20457__RESET_B repeater276/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14850_ _20079_/Q vssd1 vssd1 vccd1 vccd1 _14853_/A sky130_fd_sc_hd__inv_2
XFILLER_248_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13801_ _20624_/Q vssd1 vssd1 vccd1 vccd1 _13801_/Y sky130_fd_sc_hd__inv_2
X_14781_ _14779_/A _14779_/B _14779_/Y vssd1 vssd1 vccd1 vccd1 _20125_/D sky130_fd_sc_hd__a21oi_1
XANTENNA_input18_A HADDR[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11993_ _20987_/Q _11993_/B vssd1 vssd1 vccd1 vccd1 _11994_/B sky130_fd_sc_hd__or2_1
XFILLER_90_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16520_ _16512_/Y _16518_/Y _16519_/Y _19875_/Q vssd1 vssd1 vccd1 vccd1 _16521_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_205_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13732_ _15772_/A _15774_/A _13734_/S vssd1 vssd1 vccd1 vccd1 _20325_/D sky130_fd_sc_hd__mux2_1
XANTENNA__10457__A2 _20692_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10944_ _21210_/Q _11814_/A _10940_/Y _21025_/Q _10943_/X vssd1 vssd1 vccd1 vccd1
+ _10970_/C sky130_fd_sc_hd__o221a_1
XFILLER_17_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16451_ _16451_/A _16451_/B _16451_/C vssd1 vssd1 vccd1 vccd1 _16459_/A sky130_fd_sc_hd__or3_4
X_13663_ _20363_/Q _13659_/X _13538_/X _13662_/X vssd1 vssd1 vccd1 vccd1 _20363_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18265__S _18902_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10875_ _21261_/Q _10871_/X _09698_/X _10872_/X vssd1 vssd1 vccd1 vccd1 _21261_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19206__S1 _21006_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_231_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15402_ _19812_/Q _15398_/X _15383_/X _15400_/X vssd1 vssd1 vccd1 vccd1 _19812_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19170_ _19301_/Q _19823_/Q _19831_/Q _19415_/Q _19280_/S0 _20122_/Q vssd1 vssd1
+ vccd1 vccd1 _19170_/X sky130_fd_sc_hd__mux4_2
X_12614_ _12620_/A vssd1 vssd1 vccd1 vccd1 _12614_/X sky130_fd_sc_hd__buf_1
XPHY_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16382_ _19347_/Q _16378_/X _16200_/X _16380_/X vssd1 vssd1 vccd1 vccd1 _19347_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12603__B1 _18223_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13594_ _13594_/A vssd1 vssd1 vccd1 vccd1 _13594_/X sky130_fd_sc_hd__buf_1
XFILLER_231_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18121_ vssd1 vssd1 vccd1 vccd1 _18121_/HI _18121_/LO sky130_fd_sc_hd__conb_1
XPHY_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15333_ _20025_/Q _15329_/X _13557_/X _15330_/X vssd1 vssd1 vccd1 vccd1 _20025_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12545_ _12553_/A vssd1 vssd1 vccd1 vccd1 _12554_/A sky130_fd_sc_hd__inv_2
XANTENNA_repeater157_A _18886_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18052_ _18052_/A vssd1 vssd1 vccd1 vccd1 _18052_/Y sky130_fd_sc_hd__inv_2
X_15264_ _15260_/Y _20055_/Q _15261_/Y _20050_/Q _15263_/X vssd1 vssd1 vccd1 vccd1
+ _15285_/B sky130_fd_sc_hd__o221a_1
X_12476_ _12476_/A _12476_/B vssd1 vssd1 vccd1 vccd1 _12476_/Y sky130_fd_sc_hd__nor2_2
XFILLER_177_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17003_ _19978_/Q vssd1 vssd1 vccd1 vccd1 _17003_/Y sky130_fd_sc_hd__inv_2
XFILLER_126_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19096__S _19870_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14215_ _14215_/A _14215_/B _14215_/C vssd1 vssd1 vccd1 vccd1 _20269_/D sky130_fd_sc_hd__nor3_1
X_11427_ _11347_/B _11418_/X _11371_/B _11403_/A vssd1 vssd1 vccd1 vccd1 _21176_/D
+ sky130_fd_sc_hd__o22ai_1
X_15195_ _15195_/A vssd1 vssd1 vccd1 vccd1 _15195_/Y sky130_fd_sc_hd__inv_2
XFILLER_141_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output86_A _17936_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14146_ _20530_/Q vssd1 vssd1 vccd1 vccd1 _14146_/Y sky130_fd_sc_hd__inv_2
X_11358_ _11375_/A _21183_/Q _11374_/A _21182_/Q vssd1 vssd1 vccd1 vccd1 _11359_/A
+ sky130_fd_sc_hd__or4b_4
XFILLER_153_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17845__B2 _18064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10309_ _20716_/Q vssd1 vssd1 vccd1 vccd1 _10309_/Y sky130_fd_sc_hd__inv_2
X_18954_ _16651_/X _21082_/Q _18962_/S vssd1 vssd1 vccd1 vccd1 _18954_/X sky130_fd_sc_hd__mux2_1
X_14077_ _14077_/A _14219_/A vssd1 vssd1 vccd1 vccd1 _14078_/B sky130_fd_sc_hd__or2_2
X_11289_ _11300_/A _11299_/A vssd1 vssd1 vccd1 vccd1 _11290_/B sky130_fd_sc_hd__or2_1
XFILLER_140_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19142__S0 _19285_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_239_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13028_ _20677_/Q _13026_/X _12860_/X _13027_/X vssd1 vssd1 vccd1 vccd1 _20677_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__20880__RESET_B repeater243/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17905_ _18441_/X _17951_/A _18433_/X _17952_/A vssd1 vssd1 vccd1 vccd1 _17905_/Y
+ sky130_fd_sc_hd__a22oi_4
Xclkbuf_leaf_65_HCLK clkbuf_4_11_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _21334_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_239_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18885_ _18884_/X _10089_/Y _18885_/S vssd1 vssd1 vccd1 vccd1 _18885_/X sky130_fd_sc_hd__mux2_1
XANTENNA__16749__A _16758_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20198__RESET_B repeater193/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17836_ _21421_/Q vssd1 vssd1 vccd1 vccd1 _17836_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20127__RESET_B repeater245/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09651__A input41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17767_ _19621_/Q vssd1 vssd1 vccd1 vccd1 _17767_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13095__B1 _12954_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14979_ _20099_/Q _14977_/Y _14878_/B _14978_/X vssd1 vssd1 vccd1 vccd1 _20099_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_242_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13173__A _13714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19506_ _20327_/CLK _19506_/D vssd1 vssd1 vccd1 vccd1 _19506_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_235_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16718_ _16718_/A _18934_/X vssd1 vssd1 vccd1 vccd1 _19902_/D sky130_fd_sc_hd__and2_1
XFILLER_212_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17698_ _19331_/Q vssd1 vssd1 vccd1 vccd1 _17698_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19437_ _21453_/CLK _19437_/D vssd1 vssd1 vccd1 vccd1 _19437_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_223_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16649_ _19859_/Q _15293_/B _15294_/B vssd1 vssd1 vccd1 vccd1 _16649_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__18175__S _18875_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_4_13_0_HCLK_A clkbuf_3_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19368_ _19828_/CLK _19368_/D vssd1 vssd1 vccd1 vccd1 _19368_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18319_ _17079_/Y _12128_/Y _18908_/S vssd1 vssd1 vccd1 vccd1 _18319_/X sky130_fd_sc_hd__mux2_1
X_19299_ _20432_/CLK _19299_/D vssd1 vssd1 vccd1 vccd1 _19299_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__18903__S _18903_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21330_ _21341_/CLK _21330_/D repeater204/X vssd1 vssd1 vccd1 vccd1 _21330_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__10620__A2 _20758_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21261_ _21433_/CLK _21261_/D repeater233/X vssd1 vssd1 vccd1 vccd1 _21261_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_190_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20212_ _20220_/CLK _20212_/D repeater203/X vssd1 vssd1 vccd1 vccd1 _20212_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_190_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21192_ _21193_/CLK _21192_/D repeater224/X vssd1 vssd1 vccd1 vccd1 _21192_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__20968__RESET_B repeater186/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20143_ _21239_/CLK _20143_/D repeater249/X vssd1 vssd1 vccd1 vccd1 _20143_/Q sky130_fd_sc_hd__dfrtp_1
X_09954_ _21428_/Q _09950_/X _09676_/X _09952_/X vssd1 vssd1 vccd1 vccd1 _21428_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_143_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19133__S0 _19285_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20074_ _20075_/CLK _20074_/D repeater276/X vssd1 vssd1 vccd1 vccd1 _20074_/Q sky130_fd_sc_hd__dfrtp_4
X_09885_ _20011_/Q _09885_/B vssd1 vssd1 vccd1 vccd1 _09886_/A sky130_fd_sc_hd__nand2_1
XFILLER_100_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_opt_7_HCLK_A clkbuf_opt_7_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_245_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10439__A2 _20693_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12833__B1 _12668_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20976_ _20982_/CLK _20976_/D repeater278/X vssd1 vssd1 vccd1 vccd1 _20976_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_3825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10660_ _10660_/A _10683_/A vssd1 vssd1 vccd1 vccd1 _10661_/B sky130_fd_sc_hd__or2_1
XFILLER_213_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10591_ _10591_/A _10591_/B _10591_/C _10591_/D vssd1 vssd1 vccd1 vccd1 _10639_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__18813__S _18898_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12330_ _12330_/A _12342_/A vssd1 vssd1 vccd1 vccd1 _12331_/B sky130_fd_sc_hd__or2_2
XANTENNA__17937__B _17938_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_215_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11050__B _14309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12261_ _20937_/Q _20517_/Q _12426_/A _12260_/Y vssd1 vssd1 vccd1 vccd1 _12261_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__13010__B1 _12920_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21459_ _21459_/CLK _21459_/D repeater245/X vssd1 vssd1 vccd1 vccd1 _21459_/Q sky130_fd_sc_hd__dfrtp_4
X_14000_ _20308_/Q _13999_/Y _13885_/B _13988_/X vssd1 vssd1 vccd1 vccd1 _20308_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_5_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11212_ _21209_/Q _11206_/X _09652_/X _11208_/X vssd1 vssd1 vccd1 vccd1 _21209_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_123_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12192_ _12105_/X _20352_/Q _12089_/X _20348_/Q vssd1 vssd1 vccd1 vccd1 _12192_/X
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_88_HCLK clkbuf_4_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _21368_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_135_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11143_ _11142_/X _11128_/X _11951_/B vssd1 vssd1 vccd1 vccd1 _11143_/Y sky130_fd_sc_hd__o21ai_1
Xoutput86 _17936_/Y vssd1 vssd1 vccd1 vccd1 HRDATA[16] sky130_fd_sc_hd__clkbuf_2
XFILLER_1_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput97 _18059_/Y vssd1 vssd1 vccd1 vccd1 HRDATA[26] sky130_fd_sc_hd__clkbuf_2
XFILLER_122_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15951_ _16016_/A vssd1 vssd1 vccd1 vccd1 _15951_/X sky130_fd_sc_hd__clkbuf_2
X_11074_ _11074_/A vssd1 vssd1 vccd1 vccd1 _11075_/B sky130_fd_sc_hd__inv_2
XFILLER_95_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10127__B2 _20787_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14902_ _20578_/Q vssd1 vssd1 vccd1 vccd1 _14902_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20291__RESET_B repeater263/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10025_ _10877_/A vssd1 vssd1 vccd1 vccd1 _17060_/C sky130_fd_sc_hd__clkbuf_2
X_18670_ _18669_/X _14593_/A _18748_/S vssd1 vssd1 vccd1 vccd1 _18670_/X sky130_fd_sc_hd__mux2_1
X_15882_ _19591_/Q _15875_/X _15881_/X _15877_/X vssd1 vssd1 vccd1 vccd1 _19591_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_237_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20220__RESET_B repeater203/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17621_ _19619_/Q vssd1 vssd1 vccd1 vccd1 _17621_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14833_ _20099_/Q vssd1 vssd1 vccd1 vccd1 _14963_/C sky130_fd_sc_hd__inv_2
XANTENNA__13077__B1 _12932_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output124_A _17086_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_245_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17552_ _21068_/Q vssd1 vssd1 vccd1 vccd1 _17552_/Y sky130_fd_sc_hd__inv_2
X_14764_ _14747_/B _14548_/X _15798_/B _20130_/Q _14763_/Y vssd1 vssd1 vccd1 vccd1
+ _14769_/B sky130_fd_sc_hd__a221o_1
XFILLER_17_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11976_ _13185_/A _11961_/Y _11972_/Y _21002_/Q _11975_/X vssd1 vssd1 vccd1 vccd1
+ _21002_/D sky130_fd_sc_hd__a32o_1
XANTENNA__16015__B1 _16014_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16503_ _16503_/A _16507_/B vssd1 vssd1 vccd1 vccd1 _16503_/Y sky130_fd_sc_hd__nor2_1
X_13715_ _20332_/Q _13706_/X _13714_/X _13708_/X vssd1 vssd1 vccd1 vccd1 _20332_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_72_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10927_ _21202_/Q _21029_/Q _10925_/Y _11806_/A vssd1 vssd1 vccd1 vccd1 _10931_/C
+ sky130_fd_sc_hd__o22a_1
X_17483_ _17158_/X _17461_/X _17170_/X _17470_/X _17482_/X vssd1 vssd1 vccd1 vccd1
+ _17483_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_205_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14695_ _18247_/X _14690_/X _20164_/Q _14692_/X vssd1 vssd1 vccd1 vccd1 _20164_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_220_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19222_ _17588_/Y _17589_/Y _17590_/Y _17591_/Y _19275_/S0 _21004_/Q vssd1 vssd1
+ vccd1 vccd1 _19222_/X sky130_fd_sc_hd__mux4_2
X_13646_ _13652_/A vssd1 vssd1 vccd1 vccd1 _13646_/X sky130_fd_sc_hd__buf_1
X_16434_ _16441_/A vssd1 vssd1 vccd1 vccd1 _16434_/X sky130_fd_sc_hd__buf_1
X_10858_ _10858_/A _20887_/Q _10973_/C vssd1 vssd1 vccd1 vccd1 _13327_/C sky130_fd_sc_hd__or3_4
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16365_ _16371_/A vssd1 vssd1 vccd1 vccd1 _16365_/X sky130_fd_sc_hd__clkbuf_2
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19153_ _19763_/Q _19755_/Q _19747_/Q _19739_/Q _19285_/S0 _21017_/Q vssd1 vssd1
+ vccd1 vccd1 _19153_/X sky130_fd_sc_hd__mux4_2
XFILLER_158_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13577_ _20411_/Q _13573_/X _13422_/X _13575_/X vssd1 vssd1 vccd1 vccd1 _20411_/D
+ sky130_fd_sc_hd__a22o_1
X_10789_ _10783_/A _10783_/B _10824_/A _10784_/Y vssd1 vssd1 vccd1 vccd1 _21307_/D
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__18723__S _18849_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15316_ _21444_/Q _21443_/Q _21445_/Q _09864_/X vssd1 vssd1 vccd1 vccd1 _15316_/X
+ sky130_fd_sc_hd__a31o_1
X_18104_ _18656_/X _17219_/X _18175_/X _18064_/X _18103_/X vssd1 vssd1 vccd1 vccd1
+ _18105_/C sky130_fd_sc_hd__o221a_1
X_12528_ _12528_/A vssd1 vssd1 vccd1 vccd1 _12528_/X sky130_fd_sc_hd__buf_1
XFILLER_200_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19084_ _21049_/Q _21062_/Q _19872_/Q vssd1 vssd1 vccd1 vccd1 _19084_/X sky130_fd_sc_hd__mux2_1
X_16296_ _19390_/Q _16287_/X _16295_/X _16289_/X vssd1 vssd1 vccd1 vccd1 _19390_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_185_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15247_ _20473_/Q vssd1 vssd1 vccd1 vccd1 _17807_/A sky130_fd_sc_hd__inv_2
X_18035_ _18035_/A _18078_/B vssd1 vssd1 vccd1 vccd1 _18035_/Y sky130_fd_sc_hd__nor2_1
XFILLER_173_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12459_ _20935_/Q _12458_/Y _12448_/X _12425_/B vssd1 vssd1 vccd1 vccd1 _20935_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__14552__A _20131_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18024__A _18024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15178_ _20067_/Q _15176_/Y _15082_/B _15177_/X vssd1 vssd1 vccd1 vccd1 _20067_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_99_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20379__RESET_B repeater186/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14129_ _20549_/Q vssd1 vssd1 vccd1 vccd1 _14129_/Y sky130_fd_sc_hd__inv_2
X_19986_ _20408_/CLK _19986_/D repeater185/X vssd1 vssd1 vccd1 vccd1 _19986_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_141_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18937_ _16710_/X _21139_/Q _18946_/S vssd1 vssd1 vccd1 vccd1 _18937_/X sky130_fd_sc_hd__mux2_1
XFILLER_239_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19472__CLK _19813_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15383__A _15661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09670_ _12544_/A vssd1 vssd1 vccd1 vccd1 _09670_/X sky130_fd_sc_hd__buf_4
XFILLER_95_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18868_ _18867_/X _10940_/Y _18928_/S vssd1 vssd1 vccd1 vccd1 _18868_/X sky130_fd_sc_hd__mux2_1
XFILLER_239_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17819_ _09991_/Y _17232_/X _09890_/Y _17196_/X vssd1 vssd1 vccd1 vccd1 _17819_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_215_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13068__B1 _13006_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18799_ _18798_/X _11123_/Y _18929_/S vssd1 vssd1 vccd1 vccd1 _18799_/X sky130_fd_sc_hd__mux2_1
XFILLER_227_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20830_ _20841_/CLK _20830_/D repeater251/X vssd1 vssd1 vccd1 vccd1 _20830_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_223_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20761_ _21481_/CLK _20761_/D repeater205/X vssd1 vssd1 vccd1 vccd1 _20761_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21167__RESET_B repeater225/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20692_ _20693_/CLK _20692_/D repeater196/X vssd1 vssd1 vccd1 vccd1 _20692_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_11_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10974__B _20889_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18633__S _18748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21313_ _21321_/CLK _21313_/D repeater222/X vssd1 vssd1 vccd1 vccd1 _21313_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_191_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14740__A0 _13600_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21244_ _21433_/CLK _21244_/D repeater236/X vssd1 vssd1 vccd1 vccd1 _21244_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_117_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20731__RESET_B repeater257/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21175_ _21182_/CLK _21175_/D repeater216/X vssd1 vssd1 vccd1 vccd1 _21175_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__20049__RESET_B repeater281/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20126_ _21452_/CLK _20126_/D repeater247/X vssd1 vssd1 vccd1 vccd1 _20126_/Q sky130_fd_sc_hd__dfrtp_1
X_09937_ _10858_/A _09937_/B _10973_/C vssd1 vssd1 vccd1 vccd1 _13188_/C sky130_fd_sc_hd__or3_4
XFILLER_246_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13806__A _20603_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20057_ _20066_/CLK _20057_/D repeater281/X vssd1 vssd1 vccd1 vccd1 _20057_/Q sky130_fd_sc_hd__dfrtp_2
X_09868_ _20242_/Q _09867_/A _10843_/B _18976_/S vssd1 vssd1 vccd1 vccd1 _09869_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_219_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16245__B1 _16016_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13059__B1 _12993_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09799_ _09804_/A _09803_/A _09793_/C _21459_/Q _16620_/B vssd1 vssd1 vccd1 vccd1
+ _09800_/B sky130_fd_sc_hd__o32a_1
XFILLER_234_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18808__S _18896_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater180 _21016_/Q vssd1 vssd1 vccd1 vccd1 _19285_/S0 sky130_fd_sc_hd__clkbuf_16
XPHY_4312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater191 repeater212/X vssd1 vssd1 vccd1 vccd1 repeater191/X sky130_fd_sc_hd__buf_8
XFILLER_73_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11830_ _11825_/B _11827_/X _11829_/Y _11180_/X _11813_/A vssd1 vssd1 vccd1 vccd1
+ _11831_/A sky130_fd_sc_hd__o32a_1
XPHY_4334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10230__A _21373_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11761_ _11761_/A vssd1 vssd1 vccd1 vccd1 _11761_/Y sky130_fd_sc_hd__inv_2
XPHY_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20959_ _20981_/CLK _20959_/D repeater186/X vssd1 vssd1 vccd1 vccd1 _20959_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_42_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13500_ _13515_/A vssd1 vssd1 vccd1 vccd1 _13500_/X sky130_fd_sc_hd__buf_1
XPHY_3666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10712_ _10712_/A vssd1 vssd1 vccd1 vccd1 _10712_/X sky130_fd_sc_hd__buf_1
XPHY_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13541__A _13567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14480_ _14480_/A vssd1 vssd1 vccd1 vccd1 _14480_/Y sky130_fd_sc_hd__inv_2
XPHY_3677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11692_ _21082_/Q _11689_/X _11568_/X _11690_/X vssd1 vssd1 vccd1 vccd1 _21082_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13431_ _20476_/Q _13428_/X _13429_/X _13430_/X vssd1 vssd1 vccd1 vccd1 _20476_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_42_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10643_ _21341_/Q _10649_/A _10577_/Y _10576_/A _10642_/X vssd1 vssd1 vccd1 vccd1
+ _21341_/D sky130_fd_sc_hd__o221a_1
XFILLER_186_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17948__A _18064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13231__B1 _13146_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18543__S _18928_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16150_ _16179_/A _16150_/B _16419_/C vssd1 vssd1 vccd1 vccd1 _16158_/A sky130_fd_sc_hd__or3_4
XFILLER_127_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13362_ _20512_/Q _13358_/X _13144_/X _13360_/X vssd1 vssd1 vccd1 vccd1 _20512_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_139_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10574_ _10664_/C _10665_/A _10574_/C _10668_/A vssd1 vssd1 vccd1 vccd1 _10575_/C
+ sky130_fd_sc_hd__or4_4
X_15101_ _15096_/Y _20062_/Q _20456_/Q _15081_/A _15100_/X vssd1 vssd1 vccd1 vccd1
+ _15110_/B sky130_fd_sc_hd__a221o_1
XFILLER_10_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12313_ _12313_/A _12313_/B _12377_/A vssd1 vssd1 vccd1 vccd1 _12372_/A sky130_fd_sc_hd__or3_1
X_16081_ _16087_/A vssd1 vssd1 vccd1 vccd1 _16088_/A sky130_fd_sc_hd__inv_2
XANTENNA__15468__A _15479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13293_ _13293_/A vssd1 vssd1 vccd1 vccd1 _13293_/X sky130_fd_sc_hd__buf_1
X_15032_ _20070_/Q vssd1 vssd1 vccd1 vccd1 _15084_/A sky130_fd_sc_hd__inv_2
X_12244_ _20920_/Q vssd1 vssd1 vccd1 vccd1 _12396_/B sky130_fd_sc_hd__inv_2
X_19840_ _21151_/CLK _21055_/Q repeater223/X vssd1 vssd1 vccd1 vccd1 _19840_/Q sky130_fd_sc_hd__dfrtp_1
X_12175_ _12175_/A _12175_/B _12175_/C _12175_/D vssd1 vssd1 vccd1 vccd1 _12205_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_3_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11126_ _21003_/Q vssd1 vssd1 vccd1 vccd1 _11136_/A sky130_fd_sc_hd__inv_2
X_19771_ _19789_/CLK _19771_/D vssd1 vssd1 vccd1 vccd1 _19771_/Q sky130_fd_sc_hd__dfxtp_1
X_16983_ _19973_/Q vssd1 vssd1 vccd1 vccd1 _16983_/Y sky130_fd_sc_hd__inv_2
XFILLER_111_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18722_ _18848_/A0 _14142_/Y _18902_/S vssd1 vssd1 vccd1 vccd1 _18722_/X sky130_fd_sc_hd__mux2_1
X_15934_ _15985_/A _16325_/B _15999_/C vssd1 vssd1 vccd1 vccd1 _15943_/A sky130_fd_sc_hd__or3_4
X_11057_ _11093_/A _11093_/B vssd1 vssd1 vccd1 vccd1 _11089_/A sky130_fd_sc_hd__or2_1
XANTENNA__16236__B1 _16235_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10008_ _21417_/Q vssd1 vssd1 vccd1 vccd1 _10008_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18653_ _18652_/X _17011_/Y _18875_/S vssd1 vssd1 vccd1 vccd1 _18653_/X sky130_fd_sc_hd__mux2_1
X_15865_ _15865_/A vssd1 vssd1 vccd1 vccd1 _15865_/X sky130_fd_sc_hd__buf_1
XFILLER_36_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18718__S _18880_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17604_ _11932_/X _17253_/Y _21007_/Q _17110_/Y vssd1 vssd1 vccd1 vccd1 _17604_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_91_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14816_ _20114_/Q _20115_/Q _14818_/S vssd1 vssd1 vccd1 vccd1 _20115_/D sky130_fd_sc_hd__mux2_1
X_18584_ _18583_/X _10269_/A _18841_/S vssd1 vssd1 vccd1 vccd1 _18584_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15796_ _19630_/Q _15787_/X _15795_/X _15789_/X vssd1 vssd1 vccd1 vccd1 _19630_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_189_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17535_ _21435_/Q _17776_/B vssd1 vssd1 vccd1 vccd1 _17535_/Y sky130_fd_sc_hd__nand2_1
X_14747_ _14747_/A _14747_/B vssd1 vssd1 vccd1 vccd1 _14747_/Y sky130_fd_sc_hd__nor2_1
XFILLER_51_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11959_ _21002_/Q vssd1 vssd1 vccd1 vccd1 _13185_/A sky130_fd_sc_hd__inv_2
XANTENNA__13470__B1 _13282_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14547__A _20130_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18019__A _18019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21260__RESET_B repeater233/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13451__A _15523_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14678_ _14678_/A vssd1 vssd1 vccd1 vccd1 _20171_/D sky130_fd_sc_hd__inv_2
X_17466_ _20247_/Q vssd1 vssd1 vccd1 vccd1 _17466_/Y sky130_fd_sc_hd__inv_2
XFILLER_189_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_220_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19205_ _17750_/Y _17751_/Y _17752_/Y _17753_/Y _19275_/S0 _21004_/Q vssd1 vssd1
+ vccd1 vccd1 _19205_/X sky130_fd_sc_hd__mux4_1
X_16417_ _19326_/Q _16413_/X _16212_/X _16414_/X vssd1 vssd1 vccd1 vccd1 _19326_/D
+ sky130_fd_sc_hd__a22o_1
X_13629_ _20381_/Q _13625_/X _13487_/X _13626_/X vssd1 vssd1 vccd1 vccd1 _20381_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16762__A _16779_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17397_ _17573_/A vssd1 vssd1 vccd1 vccd1 _17397_/X sky130_fd_sc_hd__buf_1
XANTENNA__18453__S _18775_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09977__B1 _09682_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19136_ _19132_/X _19133_/X _19134_/X _19135_/X _21018_/Q _21019_/Q vssd1 vssd1 vccd1
+ vccd1 _19136_/X sky130_fd_sc_hd__mux4_2
XFILLER_192_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16348_ _19365_/Q _16345_/X _16277_/X _16347_/X vssd1 vssd1 vccd1 vccd1 _19365_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_158_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15378__A _15657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19067_ _16736_/X _21143_/Q _19908_/D vssd1 vssd1 vccd1 vccd1 _19067_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16279_ _16289_/A vssd1 vssd1 vccd1 vccd1 _16279_/X sky130_fd_sc_hd__buf_1
XFILLER_218_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18018_ _18018_/A vssd1 vssd1 vccd1 vccd1 _18018_/X sky130_fd_sc_hd__buf_1
XANTENNA__14722__B1 _13704_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11536__B1 _10894_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20142__RESET_B repeater250/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19969_ _20408_/CLK _19969_/D repeater184/X vssd1 vssd1 vccd1 vccd1 _19969_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__13289__B1 _13287_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_234_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09722_ _11060_/A _20155_/Q _21235_/Q _09721_/Y vssd1 vssd1 vccd1 vccd1 _09722_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__13626__A _13626_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_234_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09653_ _21475_/Q _09643_/X _09652_/X _09646_/X vssd1 vssd1 vccd1 vccd1 _21475_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_27_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18628__S _18908_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_216_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__21348__RESET_B repeater210/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14253__A2 _14246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_242_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20813_ _21379_/CLK _20813_/D repeater212/X vssd1 vssd1 vccd1 vccd1 _20813_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_24_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17727__B1 _16631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10985__A _10985_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20744_ _21319_/CLK _20744_/D repeater191/X vssd1 vssd1 vccd1 vccd1 _20744_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20675_ _21480_/CLK _20675_/D repeater208/X vssd1 vssd1 vccd1 vccd1 _20675_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18363__S _18680_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_117_HCLK_A clkbuf_opt_3_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20912__RESET_B repeater217/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14713__B1 _12860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10290_ _10290_/A vssd1 vssd1 vccd1 vccd1 _10290_/Y sky130_fd_sc_hd__inv_2
X_21227_ _21235_/CLK _21227_/D repeater249/X vssd1 vssd1 vccd1 vccd1 _21227_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18455__A1 _20787_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21158_ _21429_/CLK _21158_/D repeater227/X vssd1 vssd1 vccd1 vccd1 _21158_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_144_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20109_ _21433_/CLK _20109_/D repeater234/X vssd1 vssd1 vccd1 vccd1 _20109_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_144_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13980_ _13987_/A vssd1 vssd1 vccd1 vccd1 _13980_/X sky130_fd_sc_hd__buf_1
X_21089_ _21424_/CLK _21089_/D repeater230/X vssd1 vssd1 vccd1 vccd1 _21089_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_74_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_118_HCLK clkbuf_opt_3_HCLK/A vssd1 vssd1 vccd1 vccd1 _20950_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_246_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12931_ _20720_/Q _12924_/X _12930_/X _12926_/X vssd1 vssd1 vccd1 vccd1 _20720_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18538__S _18910_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12862_ _20749_/Q _12859_/X _12860_/X _12861_/X vssd1 vssd1 vccd1 vccd1 _20749_/D
+ sky130_fd_sc_hd__a22o_1
X_15650_ _19696_/Q _15647_/X _15483_/X _15648_/X vssd1 vssd1 vccd1 vccd1 _19696_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21018__RESET_B repeater238/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14601_ _14595_/A _14595_/B _14636_/A _14596_/Y vssd1 vssd1 vccd1 vccd1 _20206_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_73_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11813_ _11813_/A _11828_/A vssd1 vssd1 vccd1 vccd1 _11824_/A sky130_fd_sc_hd__or2_1
X_15581_ _19731_/Q _15576_/X _15550_/X _15578_/X vssd1 vssd1 vccd1 vccd1 _19731_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12793_ _20784_/Q _12791_/X _09655_/X _12792_/X vssd1 vssd1 vccd1 vccd1 _20784_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14532_ _16484_/A _14661_/B vssd1 vssd1 vccd1 vccd1 _14656_/A sky130_fd_sc_hd__nand2_1
X_17320_ _17320_/A vssd1 vssd1 vccd1 vccd1 _17320_/X sky130_fd_sc_hd__buf_1
XPHY_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11744_ _21056_/Q _11735_/X _11743_/X _11737_/X vssd1 vssd1 vccd1 vccd1 _21056_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_53_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14463_ _14463_/A _14463_/B _14463_/C _14463_/D vssd1 vssd1 vccd1 vccd1 _14465_/C
+ sky130_fd_sc_hd__or4_4
X_17251_ _19399_/Q vssd1 vssd1 vccd1 vccd1 _17251_/Y sky130_fd_sc_hd__inv_2
XPHY_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11675_ _11675_/A vssd1 vssd1 vccd1 vccd1 _21089_/D sky130_fd_sc_hd__inv_2
XFILLER_41_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18273__S _18906_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13204__B1 _13001_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09959__B1 _09688_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16202_ _21451_/Q vssd1 vssd1 vccd1 vccd1 _16202_/X sky130_fd_sc_hd__buf_1
X_13414_ _20482_/Q _13410_/X _13221_/X _13411_/X vssd1 vssd1 vccd1 vccd1 _20482_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10626_ _20756_/Q vssd1 vssd1 vccd1 vccd1 _10626_/Y sky130_fd_sc_hd__inv_2
XFILLER_174_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17182_ _20633_/Q _17187_/B vssd1 vssd1 vccd1 vccd1 _17182_/Y sky130_fd_sc_hd__nor2_1
X_14394_ _14394_/A _14394_/B _14391_/X _14393_/X vssd1 vssd1 vccd1 vccd1 _14401_/B
+ sky130_fd_sc_hd__or4bb_4
XFILLER_127_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16133_ _16143_/A vssd1 vssd1 vccd1 vccd1 _16133_/X sky130_fd_sc_hd__buf_1
X_13345_ _13351_/A vssd1 vssd1 vccd1 vccd1 _13345_/X sky130_fd_sc_hd__buf_1
XANTENNA__20838__CLK _20930_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10557_ _10557_/A vssd1 vssd1 vccd1 vccd1 _10659_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_repeater237_A repeater238/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_39_HCLK_A _20004_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16064_ _16071_/A vssd1 vssd1 vccd1 vccd1 _16064_/X sky130_fd_sc_hd__buf_1
XFILLER_142_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13276_ _13293_/A vssd1 vssd1 vccd1 vccd1 _13276_/X sky130_fd_sc_hd__buf_1
X_10488_ _10778_/A _20691_/Q _10764_/A _20677_/Q vssd1 vssd1 vccd1 vccd1 _10488_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_142_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15015_ _15015_/A vssd1 vssd1 vccd1 vccd1 _15015_/Y sky130_fd_sc_hd__inv_2
XFILLER_170_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12227_ _20940_/Q vssd1 vssd1 vccd1 vccd1 _12228_/A sky130_fd_sc_hd__inv_2
XANTENNA__14180__A1 _20288_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16457__B1 _11504_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19823_ _21452_/CLK _19823_/D vssd1 vssd1 vccd1 vccd1 _19823_/Q sky130_fd_sc_hd__dfxtp_1
X_12158_ _12330_/A _20359_/Q _12089_/X _20348_/Q _12157_/X vssd1 vssd1 vccd1 vccd1
+ _12158_/X sky130_fd_sc_hd__o221a_1
XFILLER_150_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13446__A _15424_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11109_ _21228_/Q _11109_/B vssd1 vssd1 vccd1 vccd1 _11109_/Y sky130_fd_sc_hd__nor2_1
X_19754_ _19765_/CLK _19754_/D vssd1 vssd1 vccd1 vccd1 _19754_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16966_ _16966_/A _16966_/B vssd1 vssd1 vccd1 vccd1 _16966_/Y sky130_fd_sc_hd__nor2_1
X_12089_ _12319_/A vssd1 vssd1 vccd1 vccd1 _12089_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_49_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18705_ _17702_/X _19339_/Q _18926_/S vssd1 vssd1 vccd1 vccd1 _18705_/X sky130_fd_sc_hd__mux2_1
X_15917_ _19574_/Q _15911_/X _15916_/X _15912_/X vssd1 vssd1 vccd1 vccd1 _19574_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_65_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19685_ _19813_/CLK _19685_/D vssd1 vssd1 vccd1 vccd1 _19685_/Q sky130_fd_sc_hd__dfxtp_1
X_16897_ _19952_/Q _16892_/A _19953_/Q vssd1 vssd1 vccd1 vccd1 _16897_/X sky130_fd_sc_hd__o21a_1
XFILLER_49_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13691__B1 _12855_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18448__S _18841_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15661__A _15661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18636_ _18635_/X _10783_/A _18898_/S vssd1 vssd1 vccd1 vccd1 _18636_/X sky130_fd_sc_hd__mux2_1
X_15848_ _15885_/A _17254_/A vssd1 vssd1 vccd1 vccd1 _15856_/A sky130_fd_sc_hd__or2_2
XFILLER_224_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18567_ _18566_/X _14934_/Y _18907_/S vssd1 vssd1 vccd1 vccd1 _18567_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13443__B1 _13442_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14277__A _20122_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15779_ _15787_/A vssd1 vssd1 vccd1 vccd1 _15779_/X sky130_fd_sc_hd__buf_1
X_17518_ _19434_/Q vssd1 vssd1 vccd1 vccd1 _17518_/Y sky130_fd_sc_hd__inv_2
XFILLER_220_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18498_ _18497_/X _12234_/Y _18910_/S vssd1 vssd1 vccd1 vccd1 _18498_/X sky130_fd_sc_hd__mux2_1
XFILLER_178_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17449_ _17449_/A _20112_/Q vssd1 vssd1 vccd1 vccd1 _17449_/X sky130_fd_sc_hd__and2_1
XANTENNA__18183__S _18748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20460_ _20495_/CLK _20460_/D repeater276/X vssd1 vssd1 vccd1 vccd1 _20460_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18134__A0 _18848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19119_ _19882_/Q _16569_/X _19908_/Q vssd1 vssd1 vccd1 vccd1 _19119_/X sky130_fd_sc_hd__mux2_1
XANTENNA__20394__RESET_B repeater270/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20391_ _20950_/CLK _20391_/D repeater278/X vssd1 vssd1 vccd1 vccd1 _20391_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_173_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21012_ _21121_/CLK _21012_/D repeater238/X vssd1 vssd1 vccd1 vccd1 _21012_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_248_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09705_ _14528_/A vssd1 vssd1 vccd1 vccd1 _09780_/A sky130_fd_sc_hd__buf_1
XANTENNA__18358__S _18909_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_243_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__21182__RESET_B repeater216/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_216_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09636_ input46/X vssd1 vssd1 vccd1 vccd1 _09636_/X sky130_fd_sc_hd__buf_4
XFILLER_16_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13434__B1 _13311_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_231_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20727_ _21375_/CLK _20727_/D repeater257/X vssd1 vssd1 vccd1 vccd1 _20727_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_211_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11460_ _11462_/A vssd1 vssd1 vccd1 vccd1 _11480_/A sky130_fd_sc_hd__clkbuf_2
XPHY_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18125__A0 _18848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20658_ _20665_/CLK _20658_/D repeater261/X vssd1 vssd1 vccd1 vccd1 _20658_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_128_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10411_ _10266_/A _10266_/B _10409_/Y _10397_/X vssd1 vssd1 vccd1 vccd1 _21350_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_137_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18676__A1 _19206_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11391_ _11412_/B _11409_/B vssd1 vssd1 vccd1 vccd1 _16596_/A sky130_fd_sc_hd__or2_1
XFILLER_192_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18821__S _18909_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20589_ _20590_/CLK _20589_/D repeater260/X vssd1 vssd1 vccd1 vccd1 _20589_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_192_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13130_ _20620_/Q _13126_/X _12920_/X _13127_/X vssd1 vssd1 vccd1 vccd1 _20620_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_99_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10342_ _20715_/Q vssd1 vssd1 vccd1 vccd1 _10342_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13061_ _13073_/A vssd1 vssd1 vccd1 vccd1 _13061_/X sky130_fd_sc_hd__buf_1
XFILLER_79_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10273_ _10273_/A _10273_/B vssd1 vssd1 vccd1 vccd1 _10394_/A sky130_fd_sc_hd__or2_1
XFILLER_79_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12012_ _12030_/A vssd1 vssd1 vccd1 vccd1 _12012_/X sky130_fd_sc_hd__buf_1
XANTENNA__16439__B1 _11504_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input48_A HWDATA[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16820_ _16820_/A _16820_/B vssd1 vssd1 vccd1 vccd1 _16820_/Y sky130_fd_sc_hd__nor2_1
XFILLER_238_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16751_ _19919_/Q vssd1 vssd1 vccd1 vccd1 _16753_/A sky130_fd_sc_hd__inv_2
XFILLER_120_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13963_ _13990_/A vssd1 vssd1 vccd1 vccd1 _14070_/B sky130_fd_sc_hd__inv_2
XFILLER_101_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18268__S _18885_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15481__A _15481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15702_ _19672_/Q _15696_/X _15701_/X _15698_/X vssd1 vssd1 vccd1 vccd1 _19672_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_246_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19470_ _19776_/CLK _19470_/D vssd1 vssd1 vccd1 vccd1 _19470_/Q sky130_fd_sc_hd__dfxtp_1
X_12914_ _20727_/Q _12909_/X _12670_/X _12910_/X vssd1 vssd1 vccd1 vccd1 _20727_/D
+ sky130_fd_sc_hd__a22o_1
X_16682_ _20001_/Q _18948_/X _16680_/B _16681_/X vssd1 vssd1 vccd1 vccd1 _16682_/X
+ sky130_fd_sc_hd__a22o_1
X_13894_ _13894_/A _13894_/B _13979_/A vssd1 vssd1 vccd1 vccd1 _13895_/A sky130_fd_sc_hd__or3_1
XFILLER_206_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18421_ _18848_/A0 _17884_/Y _18874_/S vssd1 vssd1 vccd1 vccd1 _18421_/X sky130_fd_sc_hd__mux2_1
X_12845_ _20755_/Q _12841_/X _09636_/X _12842_/X vssd1 vssd1 vccd1 vccd1 _20755_/D
+ sky130_fd_sc_hd__a22o_1
X_15633_ _15633_/A vssd1 vssd1 vccd1 vccd1 _15633_/X sky130_fd_sc_hd__buf_1
XFILLER_206_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13425__B1 _13424_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18352_ _18007_/Y _16842_/Y _18875_/S vssd1 vssd1 vccd1 vccd1 _18352_/X sky130_fd_sc_hd__mux2_1
XFILLER_187_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15564_ _19741_/Q _15561_/X _15544_/X _15563_/X vssd1 vssd1 vccd1 vccd1 _19741_/D
+ sky130_fd_sc_hd__a22o_1
X_12776_ _20793_/Q _12771_/X _09628_/X _12772_/X vssd1 vssd1 vccd1 vccd1 _20793_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17303_ _21137_/Q vssd1 vssd1 vccd1 vccd1 _17303_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14515_ _14515_/A vssd1 vssd1 vccd1 vccd1 _14520_/A sky130_fd_sc_hd__inv_2
XANTENNA__19099__S _19870_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11727_ _11735_/A vssd1 vssd1 vccd1 vccd1 _11727_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_9_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15495_ _19773_/Q _15492_/X _15450_/X _15494_/X vssd1 vssd1 vccd1 vccd1 _19773_/D
+ sky130_fd_sc_hd__a22o_1
X_18283_ _18282_/X _10080_/Y _18644_/S vssd1 vssd1 vccd1 vccd1 _18283_/X sky130_fd_sc_hd__mux2_1
XPHY_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17234_ _18875_/X _17224_/X _18925_/X _17227_/X _17233_/X vssd1 vssd1 vccd1 vccd1
+ _17235_/D sky130_fd_sc_hd__o221a_2
XANTENNA__17201__A _17201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11658_ _11658_/A vssd1 vssd1 vccd1 vccd1 _19112_/S sky130_fd_sc_hd__buf_1
X_14446_ _20028_/Q vssd1 vssd1 vccd1 vccd1 _14446_/Y sky130_fd_sc_hd__inv_2
XFILLER_174_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10609_ _20754_/Q vssd1 vssd1 vccd1 vccd1 _10609_/Y sky130_fd_sc_hd__inv_2
XPHY_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14377_ _14465_/A _14471_/A vssd1 vssd1 vccd1 vccd1 _14378_/B sky130_fd_sc_hd__or2_2
XANTENNA_clkbuf_leaf_100_HCLK_A clkbuf_4_13_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17165_ _20244_/Q vssd1 vssd1 vccd1 vccd1 _17165_/Y sky130_fd_sc_hd__inv_2
X_11589_ _21123_/Q vssd1 vssd1 vccd1 vccd1 _11589_/Y sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_163_HCLK_A clkbuf_opt_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13328_ _13328_/A _17217_/A vssd1 vssd1 vccd1 vccd1 _13657_/B sky130_fd_sc_hd__or2_2
X_16116_ _19475_/Q _16108_/X _16115_/X _16111_/X vssd1 vssd1 vccd1 vccd1 _19475_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_182_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17096_ _19470_/Q vssd1 vssd1 vccd1 vccd1 _17096_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14153__A1 _20552_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18419__A1 _20648_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16047_ _19510_/Q _16042_/X _16016_/X _16043_/X vssd1 vssd1 vccd1 vccd1 _19510_/D
+ sky130_fd_sc_hd__a22o_1
X_13259_ _17085_/A _13259_/B vssd1 vssd1 vccd1 vccd1 _13260_/S sky130_fd_sc_hd__or2_1
XFILLER_143_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17890__A2 _18020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09654__A input40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19092__A1 _21086_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19806_ _19820_/CLK _19806_/D vssd1 vssd1 vccd1 vccd1 _19806_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17998_ _18347_/X _17931_/X _18151_/X _17995_/X _17997_/X vssd1 vssd1 vccd1 vccd1
+ _17999_/C sky130_fd_sc_hd__o221a_1
XFILLER_245_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_238_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19737_ _21011_/CLK _19737_/D vssd1 vssd1 vccd1 vccd1 _19737_/Q sky130_fd_sc_hd__dfxtp_1
X_16949_ _19966_/Q _16949_/B vssd1 vssd1 vccd1 vccd1 _16958_/C sky130_fd_sc_hd__or2_2
XFILLER_49_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18178__S _18898_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13664__B1 _13543_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_238_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19668_ _19812_/CLK _19668_/D vssd1 vssd1 vccd1 vccd1 _19668_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18619_ _18618_/X _20288_/Q _18904_/S vssd1 vssd1 vccd1 vccd1 _18619_/X sky130_fd_sc_hd__mux2_1
XFILLER_198_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12219__B2 _20504_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_241_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19599_ _19821_/CLK _19599_/D vssd1 vssd1 vccd1 vccd1 _19599_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18906__S _18906_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18355__A0 _18848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20512_ _20947_/CLK _20512_/D repeater267/X vssd1 vssd1 vccd1 vccd1 _20512_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__20504__RESET_B repeater267/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19406__CLK _19813_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20443_ _20476_/CLK _20443_/D repeater280/X vssd1 vssd1 vccd1 vccd1 _20443_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18641__S _18906_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_opt_0_HCLK clkbuf_opt_0_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_opt_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_16
X_20374_ _20957_/CLK _20374_/D repeater186/X vssd1 vssd1 vccd1 vccd1 _20374_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_107_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15341__B1 _14262_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_22_HCLK_A clkbuf_4_3_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17881__A2 _17839_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_85_HCLK_A clkbuf_4_12_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21363__RESET_B repeater254/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13655__B1 _13452_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10960_ _10958_/Y _21032_/Q _21205_/Q _11845_/A vssd1 vssd1 vccd1 vccd1 _10960_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__18594__A0 _17079_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09619_ _09672_/A vssd1 vssd1 vccd1 vccd1 _09657_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_43_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13407__B1 _13209_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10891_ _21255_/Q _10888_/X _10889_/X _10890_/X vssd1 vssd1 vccd1 vccd1 _21255_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18816__S _18850_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12630_ input32/X _12625_/X _20852_/Q _12626_/X vssd1 vssd1 vccd1 vccd1 _20852_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_43_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12561_ _19983_/Q _12561_/B vssd1 vssd1 vccd1 vccd1 _12562_/A sky130_fd_sc_hd__and2_1
XPHY_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11512_ _16711_/A _11497_/A _11508_/Y _11509_/Y _11523_/S vssd1 vssd1 vccd1 vccd1
+ _11513_/A sky130_fd_sc_hd__o32a_1
X_14300_ _15574_/A _15335_/B _14315_/A vssd1 vssd1 vccd1 vccd1 _14300_/Y sky130_fd_sc_hd__o21ai_1
XPHY_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15280_ _20469_/Q _15128_/X _17540_/A _20048_/Q _15279_/X vssd1 vssd1 vccd1 vccd1
+ _15284_/C sky130_fd_sc_hd__o221a_1
XPHY_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12492_ _12492_/A _12492_/B _12496_/C vssd1 vssd1 vccd1 vccd1 _20921_/D sky130_fd_sc_hd__nor3_1
XPHY_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14231_ _19890_/Q _19891_/Q vssd1 vssd1 vccd1 vccd1 _14232_/B sky130_fd_sc_hd__or2_1
XPHY_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11443_ _21155_/Q _11443_/B vssd1 vssd1 vccd1 vccd1 _11444_/B sky130_fd_sc_hd__or2_1
XPHY_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15580__B1 _15548_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18551__S _18885_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14162_ _14159_/Y _20280_/Q _14160_/Y _20268_/Q _14161_/X vssd1 vssd1 vccd1 vccd1
+ _14170_/B sky130_fd_sc_hd__o221a_1
X_11374_ _11374_/A _11783_/C vssd1 vssd1 vccd1 vccd1 _11375_/B sky130_fd_sc_hd__or2_1
XFILLER_4_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13113_ _13138_/A vssd1 vssd1 vccd1 vccd1 _13141_/A sky130_fd_sc_hd__inv_2
X_10325_ _20720_/Q vssd1 vssd1 vccd1 vccd1 _17943_/A sky130_fd_sc_hd__inv_2
X_18970_ _11542_/A _12506_/B _20917_/Q vssd1 vssd1 vccd1 vccd1 _18970_/X sky130_fd_sc_hd__mux2_1
X_14093_ _14093_/A _14093_/B vssd1 vssd1 vccd1 vccd1 _14187_/A sky130_fd_sc_hd__or2_1
XANTENNA__17872__A2 _17839_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15332__B1 _13555_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13044_ _20667_/Q _13040_/X _12881_/X _13041_/X vssd1 vssd1 vccd1 vccd1 _20667_/D
+ sky130_fd_sc_hd__a22o_1
X_17921_ _20827_/Q vssd1 vssd1 vccd1 vccd1 _17921_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19074__A1 _21136_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10256_ _21347_/Q vssd1 vssd1 vccd1 vccd1 _10263_/A sky130_fd_sc_hd__inv_2
XFILLER_239_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11509__A _16338_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17852_ _17852_/A vssd1 vssd1 vccd1 vccd1 _17852_/X sky130_fd_sc_hd__clkbuf_4
X_10187_ _10187_/A vssd1 vssd1 vccd1 vccd1 _10187_/Y sky130_fd_sc_hd__inv_2
XFILLER_227_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__21033__RESET_B repeater242/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16803_ _16848_/A vssd1 vssd1 vccd1 vccd1 _16803_/X sky130_fd_sc_hd__buf_1
XFILLER_120_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17783_ _21087_/Q vssd1 vssd1 vccd1 vccd1 _17783_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14995_ _20089_/Q _14994_/Y _14973_/X _14868_/B vssd1 vssd1 vccd1 vccd1 _20089_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_82_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19522_ _20327_/CLK _19522_/D vssd1 vssd1 vccd1 vccd1 _19522_/Q sky130_fd_sc_hd__dfxtp_1
X_16734_ _20996_/Q _12002_/B _12003_/B vssd1 vssd1 vccd1 vccd1 _16734_/X sky130_fd_sc_hd__a21bo_1
XFILLER_35_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13946_ _13942_/Y _20292_/Q _13943_/Y _20294_/Q _13945_/X vssd1 vssd1 vccd1 vccd1
+ _13947_/D sky130_fd_sc_hd__o221a_1
XANTENNA__18585__A0 _17079_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19453_ _21453_/CLK _19453_/D vssd1 vssd1 vccd1 vccd1 _19453_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16665_ _21153_/Q _21152_/Q _11442_/B vssd1 vssd1 vccd1 vccd1 _16665_/X sky130_fd_sc_hd__a21bo_1
XFILLER_61_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18726__S _18784_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13877_ _14011_/A _14010_/C _13877_/C _13877_/D vssd1 vssd1 vccd1 vccd1 _13974_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_62_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18404_ _17807_/Y _20441_/Q _18906_/S vssd1 vssd1 vccd1 vccd1 _18404_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15616_ _19715_/Q _15611_/X _15475_/X _15613_/X vssd1 vssd1 vccd1 vccd1 _19715_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_201_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12828_ _20766_/Q _12821_/X _12660_/X _12824_/X vssd1 vssd1 vccd1 vccd1 _20766_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_50_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19384_ _19521_/CLK _19384_/D vssd1 vssd1 vccd1 vccd1 _19384_/Q sky130_fd_sc_hd__dfxtp_1
X_16596_ _16596_/A _16596_/B _16596_/C _16596_/D vssd1 vssd1 vccd1 vccd1 _16596_/X
+ sky130_fd_sc_hd__or4_4
XFILLER_15_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18335_ _18334_/X _20283_/Q _18904_/S vssd1 vssd1 vccd1 vccd1 _18335_/X sky130_fd_sc_hd__mux2_1
X_15547_ _19749_/Q _15543_/X _15544_/X _15546_/X vssd1 vssd1 vccd1 vccd1 _19749_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12759_ _12785_/A vssd1 vssd1 vccd1 vccd1 _12778_/A sky130_fd_sc_hd__buf_1
XFILLER_188_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09649__A _12855_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18266_ _18265_/X _13931_/Y _18903_/S vssd1 vssd1 vccd1 vccd1 _18266_/X sky130_fd_sc_hd__mux2_1
X_15478_ _19778_/Q _15468_/X _15477_/X _15471_/X vssd1 vssd1 vccd1 vccd1 _19778_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_30_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17217_ _17217_/A vssd1 vssd1 vccd1 vccd1 _17581_/A sky130_fd_sc_hd__buf_1
X_14429_ _14427_/Y _20216_/Q _21470_/Q _14501_/A _14428_/X vssd1 vssd1 vccd1 vccd1
+ _14434_/C sky130_fd_sc_hd__o221a_1
X_18197_ _18196_/X _10772_/A _18617_/S vssd1 vssd1 vccd1 vccd1 _18197_/X sky130_fd_sc_hd__mux2_1
XANTENNA__18461__S _18884_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17148_ _21064_/Q vssd1 vssd1 vccd1 vccd1 _17148_/Y sky130_fd_sc_hd__inv_2
XFILLER_144_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17312__B2 _17232_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15386__A _15663_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09970_ _09976_/A vssd1 vssd1 vccd1 vccd1 _09970_/X sky130_fd_sc_hd__buf_1
X_17079_ _17174_/B vssd1 vssd1 vccd1 vccd1 _17079_/Y sky130_fd_sc_hd__clkinv_16
XFILLER_104_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17863__A2 _17839_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20556__CLK _20592_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20090_ _20495_/CLK _20090_/D repeater273/X vssd1 vssd1 vccd1 vccd1 _20090_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_124_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19160__S1 _21017_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13637__B1 _13424_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20992_ _21338_/CLK _20992_/D repeater222/X vssd1 vssd1 vccd1 vccd1 _20992_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_225_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20756__RESET_B repeater205/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18636__S _18898_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11154__A _20891_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_3_0_HCLK clkbuf_2_3_0_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__17000__B1 _16984_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15011__C1 _14970_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21475_ _21477_/CLK _21475_/D repeater201/X vssd1 vssd1 vccd1 vccd1 _21475_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__18371__S _18909_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20426_ _20951_/CLK _20426_/D repeater269/X vssd1 vssd1 vccd1 vccd1 _20426_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_146_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18500__A0 _18499_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20357_ _20980_/CLK _20357_/D repeater279/X vssd1 vssd1 vccd1 vccd1 _20357_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_134_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10110_ _21400_/Q _20797_/Q _21400_/Q _20797_/Q vssd1 vssd1 vccd1 vccd1 _10110_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_136_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11090_ _21233_/Q _11090_/B vssd1 vssd1 vccd1 vccd1 _11090_/Y sky130_fd_sc_hd__nor2_1
X_20288_ _20665_/CLK _20288_/D repeater261/X vssd1 vssd1 vccd1 vccd1 _20288_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_121_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10041_ _10041_/A _10041_/B _10221_/C vssd1 vssd1 vccd1 vccd1 _10200_/C sky130_fd_sc_hd__or3_1
XFILLER_195_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13800_ _20599_/Q vssd1 vssd1 vccd1 vccd1 _13800_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11992_ _20986_/Q _11992_/B vssd1 vssd1 vccd1 vccd1 _11993_/B sky130_fd_sc_hd__or2_1
X_14780_ _14779_/A _14315_/A _15574_/A _14779_/Y vssd1 vssd1 vccd1 vccd1 _20126_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_17_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13731_ _20325_/Q vssd1 vssd1 vccd1 vccd1 _15774_/A sky130_fd_sc_hd__buf_1
XFILLER_72_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10943_ _10941_/Y _21036_/Q _21209_/Q _11813_/A vssd1 vssd1 vccd1 vccd1 _10943_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_90_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18546__S _18617_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16450_ _17054_/B _11457_/C _19851_/D _19308_/Q _16449_/X vssd1 vssd1 vccd1 vccd1
+ _19308_/D sky130_fd_sc_hd__a32o_1
XANTENNA__18319__A0 _17079_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13662_ _13680_/A vssd1 vssd1 vccd1 vccd1 _13662_/X sky130_fd_sc_hd__buf_1
X_10874_ _21262_/Q _10871_/X _09693_/X _10872_/X vssd1 vssd1 vccd1 vccd1 _21262_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_25_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15401_ _19813_/Q _15398_/X _15378_/X _15400_/X vssd1 vssd1 vccd1 vccd1 _19813_/D
+ sky130_fd_sc_hd__a22o_1
X_12613_ _12619_/A vssd1 vssd1 vccd1 vccd1 _12613_/X sky130_fd_sc_hd__buf_1
XFILLER_43_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13593_ _20401_/Q _13588_/X _13442_/X _13589_/X vssd1 vssd1 vccd1 vccd1 _20401_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_31_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16381_ _19348_/Q _16378_/X _16196_/X _16380_/X vssd1 vssd1 vccd1 vccd1 _19348_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12603__B2 _12601_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18120_ vssd1 vssd1 vccd1 vccd1 _18120_/HI _18120_/LO sky130_fd_sc_hd__conb_1
XPHY_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12544_ _12544_/A vssd1 vssd1 vccd1 vccd1 _12544_/X sky130_fd_sc_hd__clkbuf_2
X_15332_ _20026_/Q _15329_/X _13555_/X _15330_/X vssd1 vssd1 vccd1 vccd1 _20026_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18051_ _18018_/X _18051_/B _18051_/C vssd1 vssd1 vccd1 vccd1 _18051_/Y sky130_fd_sc_hd__nand3b_4
X_15263_ _20486_/Q _15079_/A _15262_/Y _15098_/X vssd1 vssd1 vccd1 vccd1 _15263_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_8_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12475_ _12475_/A _12479_/A vssd1 vssd1 vccd1 vccd1 _12476_/B sky130_fd_sc_hd__or2_2
X_17002_ _17001_/Y _16998_/A _19977_/Q _16998_/Y _16915_/A vssd1 vssd1 vccd1 vccd1
+ _17002_/X sky130_fd_sc_hd__o221a_1
X_11426_ _11426_/A vssd1 vssd1 vccd1 vccd1 _21177_/D sky130_fd_sc_hd__inv_2
X_14214_ _14103_/X _14216_/A _14079_/A vssd1 vssd1 vccd1 vccd1 _14215_/C sky130_fd_sc_hd__o21a_1
XFILLER_126_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15194_ _15099_/X _15072_/B _15191_/Y _15193_/X vssd1 vssd1 vccd1 vccd1 _20058_/D
+ sky130_fd_sc_hd__a211oi_4
XANTENNA__21285__RESET_B repeater207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14145_ _14142_/Y _20264_/Q _20533_/Q _14073_/A _14144_/X vssd1 vssd1 vccd1 vccd1
+ _14155_/B sky130_fd_sc_hd__o221a_1
X_11357_ _11357_/A _11783_/C _11357_/C _11357_/D vssd1 vssd1 vccd1 vccd1 _11409_/A
+ sky130_fd_sc_hd__nor4_2
XFILLER_153_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17845__A2 _17324_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10308_ _20705_/Q vssd1 vssd1 vccd1 vccd1 _10308_/Y sky130_fd_sc_hd__inv_2
X_18953_ _16653_/X _21083_/Q _18962_/S vssd1 vssd1 vccd1 vccd1 _18953_/X sky130_fd_sc_hd__mux2_1
XANTENNA_output79_A _17235_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14076_ _14076_/A _14076_/B vssd1 vssd1 vccd1 vccd1 _14219_/A sky130_fd_sc_hd__or2_1
X_11288_ _20905_/Q vssd1 vssd1 vccd1 vccd1 _11290_/A sky130_fd_sc_hd__inv_2
XFILLER_193_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13027_ _13041_/A vssd1 vssd1 vccd1 vccd1 _13027_/X sky130_fd_sc_hd__buf_1
X_17904_ _18457_/X _17227_/X _18466_/X _17817_/X vssd1 vssd1 vccd1 vccd1 _17904_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_79_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19142__S1 _21017_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10239_ _21364_/Q vssd1 vssd1 vccd1 vccd1 _10279_/A sky130_fd_sc_hd__inv_2
X_18884_ _18883_/X _10316_/Y _18884_/S vssd1 vssd1 vccd1 vccd1 _18884_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17835_ _21259_/Q vssd1 vssd1 vccd1 vccd1 _17835_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13454__A _13714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17766_ _19437_/Q vssd1 vssd1 vccd1 vccd1 _17766_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18558__A0 _17281_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14978_ _14978_/A vssd1 vssd1 vccd1 vccd1 _14978_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_19_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19505_ _19521_/CLK _19505_/D vssd1 vssd1 vccd1 vccd1 _19505_/Q sky130_fd_sc_hd__dfxtp_1
X_16717_ _19902_/Q _14242_/B _14243_/B vssd1 vssd1 vccd1 vccd1 _16717_/X sky130_fd_sc_hd__a21bo_1
XFILLER_19_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13929_ _13928_/Y _13865_/B _20636_/Q _20293_/Q vssd1 vssd1 vccd1 vccd1 _13930_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_35_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17697_ _19355_/Q vssd1 vssd1 vccd1 vccd1 _17697_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18456__S _18850_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19436_ _21453_/CLK _19436_/D vssd1 vssd1 vccd1 vccd1 _19436_/Q sky130_fd_sc_hd__dfxtp_1
X_16648_ _16652_/A _18956_/X vssd1 vssd1 vccd1 vccd1 _19858_/D sky130_fd_sc_hd__and2_1
XFILLER_23_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19367_ _19828_/CLK _19367_/D vssd1 vssd1 vccd1 vccd1 _19367_/Q sky130_fd_sc_hd__dfxtp_1
X_16579_ _16495_/Y _16632_/B _16686_/A _11437_/Y _16575_/Y vssd1 vssd1 vccd1 vccd1
+ _16580_/A sky130_fd_sc_hd__o32a_1
XANTENNA__15792__B1 _15791_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18318_ _18317_/X _16847_/Y _18667_/S vssd1 vssd1 vccd1 vccd1 _18318_/X sky130_fd_sc_hd__mux2_1
XANTENNA__18730__A0 _18729_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19298_ _20432_/CLK _19298_/D vssd1 vssd1 vccd1 vccd1 _19298_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18249_ _19161_/X _20167_/Q _18249_/S vssd1 vssd1 vccd1 vccd1 _18249_/X sky130_fd_sc_hd__mux2_1
XANTENNA__18191__S _18748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21260_ _21433_/CLK _21260_/D repeater233/X vssd1 vssd1 vccd1 vccd1 _21260_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_190_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20211_ _21476_/CLK _20211_/D repeater203/X vssd1 vssd1 vccd1 vccd1 _20211_/Q sky130_fd_sc_hd__dfrtp_1
X_21191_ _21191_/CLK _21191_/D repeater224/X vssd1 vssd1 vccd1 vccd1 _21191_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_171_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20142_ _20142_/CLK _20142_/D repeater250/X vssd1 vssd1 vccd1 vccd1 _20142_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_103_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09953_ _21429_/Q _09950_/X _09670_/X _09952_/X vssd1 vssd1 vccd1 vccd1 _21429_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19133__S1 _21017_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20073_ _20075_/CLK _20073_/D repeater276/X vssd1 vssd1 vccd1 vccd1 _20073_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_58_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09884_ _09884_/A vssd1 vssd1 vccd1 vccd1 _09885_/B sky130_fd_sc_hd__inv_2
XFILLER_112_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_151_HCLK clkbuf_4_4_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19961_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_26_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20590__RESET_B repeater259/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12833__A1 _20763_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20975_ _20980_/CLK _20975_/D repeater278/X vssd1 vssd1 vccd1 vccd1 _20975_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_4549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18366__S _18875_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17221__B1 _18892_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19744__CLK _19765_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12708__A _12708_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10590_ _10656_/A _20755_/Q _10651_/A _20750_/Q _10589_/X vssd1 vssd1 vccd1 vccd1
+ _10591_/D sky130_fd_sc_hd__o221a_1
XFILLER_178_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12260_ _20517_/Q vssd1 vssd1 vccd1 vccd1 _12260_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21458_ _21459_/CLK _21458_/D repeater245/X vssd1 vssd1 vccd1 vccd1 _21458_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_119_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11211_ _21210_/Q _11206_/X _09649_/X _11208_/X vssd1 vssd1 vccd1 vccd1 _21210_/D
+ sky130_fd_sc_hd__a22o_1
X_20409_ _20413_/CLK _20409_/D repeater185/X vssd1 vssd1 vccd1 vccd1 _20409_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_135_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12191_ _20358_/Q vssd1 vssd1 vccd1 vccd1 _12191_/Y sky130_fd_sc_hd__inv_2
XFILLER_162_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21389_ _21390_/CLK _21389_/D repeater239/X vssd1 vssd1 vccd1 vccd1 _21389_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_123_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11142_ _21005_/Q vssd1 vssd1 vccd1 vccd1 _11142_/X sky130_fd_sc_hd__buf_1
Xoutput87 _17957_/X vssd1 vssd1 vccd1 vccd1 HRDATA[17] sky130_fd_sc_hd__clkbuf_2
X_15950_ _19559_/Q _15943_/X _15949_/X _15945_/X vssd1 vssd1 vccd1 vccd1 _19559_/D
+ sky130_fd_sc_hd__a22o_1
X_11073_ _11063_/B _11066_/B _11072_/X _11050_/A _21237_/Q vssd1 vssd1 vccd1 vccd1
+ _21237_/D sky130_fd_sc_hd__a32o_1
XFILLER_95_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput98 _18068_/Y vssd1 vssd1 vccd1 vccd1 HRDATA[27] sky130_fd_sc_hd__clkbuf_2
XANTENNA__18788__A0 _18787_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10024_ _18984_/X _14813_/D _21410_/Q _17038_/B vssd1 vssd1 vccd1 vccd1 _21410_/D
+ sky130_fd_sc_hd__o22a_1
XANTENNA_input30_A HADDR[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14901_ _14901_/A _14901_/B _14901_/C _14900_/X vssd1 vssd1 vccd1 vccd1 _14901_/X
+ sky130_fd_sc_hd__or4b_1
X_15881_ _15881_/A vssd1 vssd1 vccd1 vccd1 _15881_/X sky130_fd_sc_hd__buf_1
XFILLER_48_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17620_ _19435_/Q vssd1 vssd1 vccd1 vccd1 _17620_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13274__A input58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14832_ _20100_/Q vssd1 vssd1 vccd1 vccd1 _14965_/B sky130_fd_sc_hd__inv_2
XANTENNA__14274__A0 _13600_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17551_ _21084_/Q vssd1 vssd1 vccd1 vccd1 _17551_/Y sky130_fd_sc_hd__inv_2
XFILLER_91_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14763_ _19124_/X vssd1 vssd1 vccd1 vccd1 _14763_/Y sky130_fd_sc_hd__inv_2
XFILLER_245_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11975_ _13175_/A _11974_/X _13185_/B _11978_/B vssd1 vssd1 vccd1 vccd1 _11975_/X
+ sky130_fd_sc_hd__a31o_1
X_16502_ _16502_/A vssd1 vssd1 vccd1 vccd1 _16507_/B sky130_fd_sc_hd__buf_1
X_13714_ _13714_/A vssd1 vssd1 vccd1 vccd1 _13714_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__20260__RESET_B repeater262/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10926_ _21029_/Q vssd1 vssd1 vccd1 vccd1 _11806_/A sky130_fd_sc_hd__inv_2
X_17482_ _17060_/B _17475_/X _17477_/X _17479_/X _17481_/X vssd1 vssd1 vccd1 vccd1
+ _17482_/X sky130_fd_sc_hd__o2111a_1
X_14694_ _18248_/X _14690_/X _20165_/Q _14692_/X vssd1 vssd1 vccd1 vccd1 _20165_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_205_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19221_ _19217_/X _19218_/X _19219_/X _19220_/X _20132_/Q _20133_/Q vssd1 vssd1 vccd1
+ vccd1 _19221_/X sky130_fd_sc_hd__mux4_2
XFILLER_71_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16433_ _16433_/A _17254_/A vssd1 vssd1 vccd1 vccd1 _16441_/A sky130_fd_sc_hd__or2_2
XFILLER_220_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13645_ _13651_/A vssd1 vssd1 vccd1 vccd1 _13645_/X sky130_fd_sc_hd__buf_1
X_10857_ _21269_/Q _10853_/X _18275_/X _10846_/X vssd1 vssd1 vccd1 vccd1 _21269_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_71_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19152_ _19683_/Q _19811_/Q _19803_/Q _19795_/Q _19285_/S0 _21017_/Q vssd1 vssd1
+ vccd1 vccd1 _19152_/X sky130_fd_sc_hd__mux4_1
X_16364_ _16370_/A vssd1 vssd1 vccd1 vccd1 _16371_/A sky130_fd_sc_hd__inv_2
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10788_ _21308_/Q _10784_/Y _10422_/Y _10784_/A _10787_/X vssd1 vssd1 vccd1 vccd1
+ _21308_/D sky130_fd_sc_hd__o221a_1
X_13576_ _20412_/Q _13573_/X _13418_/X _13575_/X vssd1 vssd1 vccd1 vccd1 _20412_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18103_ _18171_/X _17862_/A _18173_/X _18065_/X vssd1 vssd1 vccd1 vccd1 _18103_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__21466__RESET_B repeater204/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15315_ _18976_/X vssd1 vssd1 vccd1 vccd1 _15315_/Y sky130_fd_sc_hd__inv_2
X_12527_ _12527_/A vssd1 vssd1 vccd1 vccd1 _12527_/X sky130_fd_sc_hd__clkbuf_2
X_19083_ _21050_/Q _21063_/Q _19872_/Q vssd1 vssd1 vccd1 vccd1 _19083_/X sky130_fd_sc_hd__mux2_1
X_16295_ _20324_/Q vssd1 vssd1 vccd1 vccd1 _16295_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_185_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18034_ _18034_/A _18078_/B vssd1 vssd1 vccd1 vccd1 _18034_/Y sky130_fd_sc_hd__nor2_1
X_15246_ _20490_/Q vssd1 vssd1 vccd1 vccd1 _15246_/Y sky130_fd_sc_hd__inv_2
X_12458_ _12458_/A vssd1 vssd1 vccd1 vccd1 _12458_/Y sky130_fd_sc_hd__inv_2
XFILLER_126_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_32_HCLK clkbuf_opt_4_HCLK/A vssd1 vssd1 vccd1 vccd1 _21125_/CLK sky130_fd_sc_hd__clkbuf_16
X_11409_ _11409_/A _11409_/B _11409_/C _11376_/C vssd1 vssd1 vccd1 vccd1 _11776_/B
+ sky130_fd_sc_hd__or4b_4
XANTENNA__13449__A _13710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15177_ _15177_/A vssd1 vssd1 vccd1 vccd1 _15177_/X sky130_fd_sc_hd__clkbuf_2
X_12389_ _12389_/A vssd1 vssd1 vccd1 vccd1 _12389_/Y sky130_fd_sc_hd__inv_2
XFILLER_181_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14128_ _14125_/Y _20289_/Q _20560_/Q _14099_/A _14127_/X vssd1 vssd1 vccd1 vccd1
+ _14138_/B sky130_fd_sc_hd__o221a_1
X_19985_ _19985_/CLK _19985_/D repeater281/X vssd1 vssd1 vccd1 vccd1 _19985_/Q sky130_fd_sc_hd__dfstp_1
X_18936_ _16713_/X _21140_/Q _18946_/S vssd1 vssd1 vccd1 vccd1 _18936_/X sky130_fd_sc_hd__mux2_1
X_14059_ _20269_/Q vssd1 vssd1 vccd1 vccd1 _14079_/A sky130_fd_sc_hd__inv_2
XFILLER_141_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09662__A input69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_239_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18867_ _18866_/X _17252_/Y _18927_/S vssd1 vssd1 vccd1 vccd1 _18867_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17818_ _09762_/Y _17853_/A _10958_/Y _17817_/X vssd1 vssd1 vccd1 vccd1 _17818_/X
+ sky130_fd_sc_hd__o22a_1
X_18798_ _18797_/X _10948_/Y _18928_/S vssd1 vssd1 vccd1 vccd1 _18798_/X sky130_fd_sc_hd__mux2_1
XANTENNA__14265__B1 _14264_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17749_ _19725_/Q vssd1 vssd1 vccd1 vccd1 _17749_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18186__S _18896_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20760_ _21481_/CLK _20760_/D repeater201/X vssd1 vssd1 vccd1 vccd1 _20760_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_50_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19419_ _19828_/CLK _19419_/D vssd1 vssd1 vccd1 vccd1 _19419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20691_ _20693_/CLK _20691_/D repeater194/X vssd1 vssd1 vccd1 vccd1 _20691_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_195_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21312_ _21338_/CLK _21312_/D repeater222/X vssd1 vssd1 vccd1 vccd1 _21312_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_175_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21243_ _21433_/CLK _21243_/D repeater190/X vssd1 vssd1 vccd1 vccd1 _21243_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_105_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21174_ _21182_/CLK _21174_/D repeater216/X vssd1 vssd1 vccd1 vccd1 _21174_/Q sky130_fd_sc_hd__dfrtp_1
X_20125_ _21452_/CLK _20125_/D repeater247/X vssd1 vssd1 vccd1 vccd1 _20125_/Q sky130_fd_sc_hd__dfrtp_1
X_09936_ _20888_/Q vssd1 vssd1 vccd1 vccd1 _10858_/A sky130_fd_sc_hd__inv_2
XFILLER_246_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20056_ _20480_/CLK _20056_/D repeater183/X vssd1 vssd1 vccd1 vccd1 _20056_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__20771__RESET_B repeater255/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09867_ _09867_/A vssd1 vssd1 vccd1 vccd1 _09870_/A sky130_fd_sc_hd__buf_1
XFILLER_85_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09798_ _21458_/Q vssd1 vssd1 vccd1 vccd1 _16620_/B sky130_fd_sc_hd__buf_1
XFILLER_133_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater170 _18897_/S vssd1 vssd1 vccd1 vccd1 _18669_/S sky130_fd_sc_hd__buf_6
Xrepeater181 _21003_/Q vssd1 vssd1 vccd1 vccd1 _19275_/S0 sky130_fd_sc_hd__clkbuf_16
XPHY_4313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater192 repeater212/X vssd1 vssd1 vccd1 vccd1 repeater192/X sky130_fd_sc_hd__buf_8
XPHY_4324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11760_ _21053_/Q _11759_/X _19872_/Q _11755_/Y vssd1 vssd1 vccd1 vccd1 _21053_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_26_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20958_ _20981_/CLK _20958_/D repeater186/X vssd1 vssd1 vccd1 vccd1 _20958_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_4379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09683__B1 _09682_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_199_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10711_ _10711_/A vssd1 vssd1 vccd1 vccd1 _10711_/Y sky130_fd_sc_hd__inv_2
XPHY_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11691_ _21083_/Q _11689_/X _11565_/X _11690_/X vssd1 vssd1 vccd1 vccd1 _21083_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_241_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20889_ _20890_/CLK _20889_/D repeater185/X vssd1 vssd1 vccd1 vccd1 _20889_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_3689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10642_ _10694_/A vssd1 vssd1 vccd1 vccd1 _10642_/X sky130_fd_sc_hd__buf_1
XPHY_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13430_ _13447_/A vssd1 vssd1 vccd1 vccd1 _13430_/X sky130_fd_sc_hd__buf_1
XPHY_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_55_HCLK clkbuf_4_12_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _21406_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13361_ _20513_/Q _13358_/X _13140_/X _13360_/X vssd1 vssd1 vccd1 vccd1 _20513_/D
+ sky130_fd_sc_hd__a22o_1
X_10573_ _10650_/B _10573_/B _10573_/C vssd1 vssd1 vccd1 vccd1 _10668_/A sky130_fd_sc_hd__or3_1
XFILLER_167_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18170__A1 _10086_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15100_ _15097_/Y _15098_/X _20447_/Q _15099_/X vssd1 vssd1 vccd1 vccd1 _15100_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_139_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12990__B1 _12989_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12312_ _12312_/A _12312_/B vssd1 vssd1 vccd1 vccd1 _12377_/A sky130_fd_sc_hd__or2_2
XFILLER_139_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16080_ _16087_/A vssd1 vssd1 vccd1 vccd1 _16080_/X sky130_fd_sc_hd__buf_1
XFILLER_10_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13292_ _20550_/Q _13286_/X _13213_/X _13288_/X vssd1 vssd1 vccd1 vccd1 _20550_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_input78_A sda_i_S5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15031_ _20071_/Q vssd1 vssd1 vccd1 vccd1 _15085_/A sky130_fd_sc_hd__inv_2
X_12243_ _20945_/Q vssd1 vssd1 vccd1 vccd1 _12395_/B sky130_fd_sc_hd__inv_2
XFILLER_170_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12174_ _12333_/A _20362_/Q _20975_/Q _12172_/Y _12173_/X vssd1 vssd1 vccd1 vccd1
+ _12175_/D sky130_fd_sc_hd__a221o_1
XANTENNA__20859__RESET_B repeater243/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11125_ _21004_/Q vssd1 vssd1 vccd1 vccd1 _11127_/A sky130_fd_sc_hd__inv_2
X_19770_ _19789_/CLK _19770_/D vssd1 vssd1 vccd1 vccd1 _19770_/Q sky130_fd_sc_hd__dfxtp_1
X_16982_ _16980_/Y _16981_/X _16967_/X vssd1 vssd1 vccd1 vccd1 _16982_/X sky130_fd_sc_hd__o21a_1
XFILLER_123_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18721_ _18720_/X _14571_/A _18898_/S vssd1 vssd1 vccd1 vccd1 _18721_/X sky130_fd_sc_hd__mux2_2
X_15933_ _20128_/Q vssd1 vssd1 vccd1 vccd1 _15985_/A sky130_fd_sc_hd__buf_1
X_11056_ _11096_/A _11096_/B vssd1 vssd1 vccd1 vccd1 _11093_/B sky130_fd_sc_hd__nand2_1
XFILLER_77_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10007_ _20016_/Q vssd1 vssd1 vccd1 vccd1 _17032_/A sky130_fd_sc_hd__buf_1
X_18652_ _17281_/X _18092_/Y _18874_/S vssd1 vssd1 vccd1 vccd1 _18652_/X sky130_fd_sc_hd__mux2_1
X_15864_ _15875_/A vssd1 vssd1 vccd1 vccd1 _15864_/X sky130_fd_sc_hd__buf_1
XFILLER_236_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20767__CLK _21342_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16787__A2 _16777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_224_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17603_ _19403_/Q vssd1 vssd1 vccd1 vccd1 _17603_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14815_ _20115_/Q _20116_/Q _14818_/S vssd1 vssd1 vccd1 vccd1 _20116_/D sky130_fd_sc_hd__mux2_1
X_18583_ _18582_/X _10094_/Y _18885_/S vssd1 vssd1 vccd1 vccd1 _18583_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15795_ _16016_/A vssd1 vssd1 vccd1 vccd1 _15795_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_217_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17204__A _17204_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17534_ _17536_/A vssd1 vssd1 vccd1 vccd1 _17776_/B sky130_fd_sc_hd__buf_1
X_14746_ _19122_/X _14561_/Y _14745_/X vssd1 vssd1 vccd1 vccd1 _20136_/D sky130_fd_sc_hd__a21oi_1
XANTENNA__19281__S0 _20123_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11958_ _11951_/A _11136_/X _19109_/X _21003_/Q vssd1 vssd1 vccd1 vccd1 _21003_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_44_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_232_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17465_ _21144_/Q vssd1 vssd1 vccd1 vccd1 _17465_/Y sky130_fd_sc_hd__inv_2
X_10909_ _10898_/A _21247_/Q _10910_/S vssd1 vssd1 vccd1 vccd1 _21247_/D sky130_fd_sc_hd__mux2_1
XANTENNA__18734__S _18929_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14677_ _20171_/Q _10918_/B _14673_/Y _10918_/A _14676_/Y vssd1 vssd1 vccd1 vccd1
+ _14678_/A sky130_fd_sc_hd__o32a_1
XFILLER_32_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11889_ _19115_/S _11889_/B vssd1 vssd1 vccd1 vccd1 _11889_/X sky130_fd_sc_hd__or2_2
XFILLER_60_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19204_ _17746_/Y _17747_/Y _17748_/Y _17749_/Y _19275_/S0 _21004_/Q vssd1 vssd1
+ vccd1 vccd1 _19204_/X sky130_fd_sc_hd__mux4_2
X_16416_ _19327_/Q _16413_/X _16210_/X _16414_/X vssd1 vssd1 vccd1 vccd1 _19327_/D
+ sky130_fd_sc_hd__a22o_1
X_13628_ _20382_/Q _13625_/X _13485_/X _13626_/X vssd1 vssd1 vccd1 vccd1 _20382_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__20254__SET_B repeater217/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17396_ _17394_/Y _17196_/X _17395_/Y _17232_/X vssd1 vssd1 vccd1 vccd1 _17396_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_186_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19135_ _19655_/Q _19647_/Q _19631_/Q _19815_/Q _19285_/S0 _21017_/Q vssd1 vssd1
+ vccd1 vccd1 _19135_/X sky130_fd_sc_hd__mux4_2
X_16347_ _16353_/A vssd1 vssd1 vccd1 vccd1 _16347_/X sky130_fd_sc_hd__buf_1
XFILLER_158_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13559_ _13566_/A vssd1 vssd1 vccd1 vccd1 _13559_/X sky130_fd_sc_hd__buf_1
XANTENNA__18161__A1 _21485_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19066_ _19357_/Q _21127_/Q _19910_/Q vssd1 vssd1 vccd1 vccd1 _19066_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16278_ _16287_/A vssd1 vssd1 vccd1 vccd1 _16289_/A sky130_fd_sc_hd__inv_2
XFILLER_173_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18017_ _20420_/Q vssd1 vssd1 vccd1 vccd1 _18017_/Y sky130_fd_sc_hd__inv_2
X_15229_ _20487_/Q vssd1 vssd1 vccd1 vccd1 _18001_/A sky130_fd_sc_hd__inv_2
XFILLER_218_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11536__A1 _21139_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19968_ _20413_/CLK _19968_/D repeater185/X vssd1 vssd1 vccd1 vccd1 _19968_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_234_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09721_ _20155_/Q vssd1 vssd1 vccd1 vccd1 _09721_/Y sky130_fd_sc_hd__inv_2
XFILLER_228_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18919_ _18918_/X _21246_/Q _20869_/Q vssd1 vssd1 vccd1 vccd1 _18919_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19899_ _21185_/CLK _19899_/D repeater224/X vssd1 vssd1 vccd1 vccd1 _19899_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18909__S _18909_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20182__RESET_B repeater193/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09652_ _12857_/A vssd1 vssd1 vccd1 vccd1 _09652_/X sky130_fd_sc_hd__buf_4
XFILLER_216_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20812_ _21379_/CLK _20812_/D repeater213/X vssd1 vssd1 vccd1 vccd1 _20812_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_82_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19272__S0 _19275_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_78_HCLK clkbuf_4_13_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20622_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20743_ _21319_/CLK _20743_/D repeater191/X vssd1 vssd1 vccd1 vccd1 _20743_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18644__S _18644_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20674_ _21480_/CLK _20674_/D repeater208/X vssd1 vssd1 vccd1 vccd1 _20674_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11224__B1 _10892_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20039__SET_B repeater216/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12724__A0 _11179_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21226_ _21235_/CLK _21226_/D repeater249/X vssd1 vssd1 vccd1 vccd1 _21226_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_88_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17663__B1 _18721_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21157_ _21429_/CLK _21157_/D repeater229/X vssd1 vssd1 vccd1 vccd1 _21157_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_160_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20108_ _20724_/CLK _20108_/D repeater264/X vssd1 vssd1 vccd1 vccd1 _20108_/Q sky130_fd_sc_hd__dfrtp_1
X_09919_ _21244_/Q _09919_/B _21249_/Q _11591_/A vssd1 vssd1 vccd1 vccd1 _09925_/A
+ sky130_fd_sc_hd__or4_4
X_21088_ _21419_/CLK _21088_/D repeater230/X vssd1 vssd1 vccd1 vccd1 _21088_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_120_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18819__S _18907_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20039_ _21183_/CLK _20039_/D repeater216/X vssd1 vssd1 vccd1 vccd1 _20039_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_74_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12930_ input46/X vssd1 vssd1 vccd1 vccd1 _12930_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_246_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12861_ _12876_/A vssd1 vssd1 vccd1 vccd1 _12861_/X sky130_fd_sc_hd__buf_1
XFILLER_234_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14600_ _20207_/Q _14596_/Y _13832_/Y _14596_/A _14599_/X vssd1 vssd1 vccd1 vccd1
+ _20207_/D sky130_fd_sc_hd__o221a_1
XPHY_4143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11812_ _11812_/A _11832_/A vssd1 vssd1 vccd1 vccd1 _11828_/A sky130_fd_sc_hd__or2_1
XPHY_4154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15580_ _19732_/Q _15576_/X _15548_/X _15578_/X vssd1 vssd1 vccd1 vccd1 _19732_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09656__B1 _09655_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19263__S0 _19275_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12792_ _12804_/A vssd1 vssd1 vccd1 vccd1 _12792_/X sky130_fd_sc_hd__buf_1
XPHY_4176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14531_ _15832_/C vssd1 vssd1 vccd1 vccd1 _14661_/B sky130_fd_sc_hd__inv_2
XFILLER_242_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11743_ _11743_/A vssd1 vssd1 vccd1 vccd1 _11743_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_42_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18554__S _18909_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21058__RESET_B repeater212/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17250_ _19293_/Q vssd1 vssd1 vccd1 vccd1 _17250_/Y sky130_fd_sc_hd__inv_2
XPHY_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14462_ _14462_/A _14462_/B _14462_/C _14462_/D vssd1 vssd1 vccd1 vccd1 _14463_/B
+ sky130_fd_sc_hd__or4_4
XPHY_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11674_ _16654_/A _11657_/A _17046_/A _11520_/Y _11676_/S vssd1 vssd1 vccd1 vccd1
+ _11675_/A sky130_fd_sc_hd__o32a_1
XPHY_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16201_ _19436_/Q _16195_/X _16200_/X _16198_/X vssd1 vssd1 vccd1 vccd1 _19436_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13413_ _20483_/Q _13410_/X _13219_/X _13411_/X vssd1 vssd1 vccd1 vccd1 _20483_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11215__B1 _09655_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10625_ _10700_/A _20738_/Q _21324_/Q _10619_/Y _10624_/X vssd1 vssd1 vccd1 vccd1
+ _10625_/X sky130_fd_sc_hd__a221o_1
X_17181_ _20323_/Q vssd1 vssd1 vccd1 vccd1 _17181_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15479__A _15479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14393_ _20234_/Q _14392_/Y _21477_/Q _14343_/A vssd1 vssd1 vccd1 vccd1 _14393_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_139_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16132_ _16141_/A vssd1 vssd1 vccd1 vccd1 _16143_/A sky130_fd_sc_hd__inv_2
XANTENNA__11800__A _11800_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12963__B1 _12879_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10556_ _21330_/Q vssd1 vssd1 vccd1 vccd1 _10557_/A sky130_fd_sc_hd__inv_2
X_13344_ _20522_/Q _13339_/X _13284_/X _13340_/X vssd1 vssd1 vccd1 vccd1 _20522_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_185_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16063_ _16247_/A _16107_/B _16344_/C vssd1 vssd1 vccd1 vccd1 _16071_/A sky130_fd_sc_hd__or3_4
X_10487_ _21288_/Q vssd1 vssd1 vccd1 vccd1 _10764_/A sky130_fd_sc_hd__inv_2
XANTENNA__15901__B1 _15795_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13275_ _20558_/Q _13264_/X _13274_/X _13268_/X vssd1 vssd1 vccd1 vccd1 _20558_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_170_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15014_ _15002_/A _15002_/B _15012_/Y _14970_/X vssd1 vssd1 vccd1 vccd1 _20082_/D
+ sky130_fd_sc_hd__a211oi_2
X_12226_ _20930_/Q vssd1 vssd1 vccd1 vccd1 _12419_/A sky130_fd_sc_hd__inv_2
XFILLER_97_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12157_ _12036_/X _20346_/Q _12324_/A _20353_/Q vssd1 vssd1 vccd1 vccd1 _12157_/X
+ sky130_fd_sc_hd__o22a_1
X_19822_ _19835_/CLK _19822_/D vssd1 vssd1 vccd1 vccd1 _19822_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13727__A _13727_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11108_ _11108_/A vssd1 vssd1 vccd1 vccd1 _11109_/B sky130_fd_sc_hd__inv_2
XFILLER_238_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16965_ _16965_/A vssd1 vssd1 vccd1 vccd1 _16965_/Y sky130_fd_sc_hd__inv_2
X_12088_ _20966_/Q vssd1 vssd1 vccd1 vccd1 _12319_/A sky130_fd_sc_hd__inv_2
X_19753_ _21011_/CLK _19753_/D vssd1 vssd1 vccd1 vccd1 _19753_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18729__S _18787_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15916_ _16163_/A vssd1 vssd1 vccd1 vccd1 _15916_/X sky130_fd_sc_hd__clkbuf_2
X_11039_ _19967_/Q _19968_/Q _11039_/C _16979_/A vssd1 vssd1 vccd1 vccd1 _11040_/B
+ sky130_fd_sc_hd__or4_1
X_18704_ _17703_/X _20150_/Q _18928_/S vssd1 vssd1 vccd1 vccd1 _18704_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19684_ _19812_/CLK _19684_/D vssd1 vssd1 vccd1 vccd1 _19684_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16896_ _16896_/A vssd1 vssd1 vccd1 vccd1 _16902_/B sky130_fd_sc_hd__inv_2
XANTENNA__13691__A1 _20345_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18635_ _18634_/X _10615_/Y _18891_/S vssd1 vssd1 vccd1 vccd1 _18635_/X sky130_fd_sc_hd__mux2_1
XFILLER_237_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15847_ _15847_/A _15847_/B vssd1 vssd1 vccd1 vccd1 _17254_/A sky130_fd_sc_hd__or2_2
XFILLER_92_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_123_HCLK_A clkbuf_4_4_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18566_ _18565_/X _15138_/Y _18906_/S vssd1 vssd1 vccd1 vccd1 _18566_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09647__B1 _09645_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19254__S0 _19275_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15778_ _16311_/A _15778_/B _15778_/C vssd1 vssd1 vccd1 vccd1 _15787_/A sky130_fd_sc_hd__or3_4
XFILLER_17_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__21481__RESET_B repeater200/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17517_ _19490_/Q vssd1 vssd1 vccd1 vccd1 _17517_/Y sky130_fd_sc_hd__inv_2
X_14729_ _16487_/A vssd1 vssd1 vccd1 vccd1 _17774_/B sky130_fd_sc_hd__buf_1
XFILLER_21_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18497_ _18496_/X _12179_/Y _18787_/S vssd1 vssd1 vccd1 vccd1 _18497_/X sky130_fd_sc_hd__mux2_2
XANTENNA__18464__S _18775_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_232_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17448_ _21434_/Q _17536_/A vssd1 vssd1 vccd1 vccd1 _17448_/X sky130_fd_sc_hd__and2_1
XFILLER_178_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_7_HCLK clkbuf_opt_2_HCLK/A vssd1 vssd1 vccd1 vccd1 _19521_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__15389__A _15389_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17379_ _21066_/Q vssd1 vssd1 vccd1 vccd1 _17379_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14293__A _20123_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11710__A _21071_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19118_ _19115_/S _10985_/Y _19118_/S vssd1 vssd1 vccd1 vccd1 _19118_/X sky130_fd_sc_hd__mux2_1
XFILLER_192_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20390_ _20980_/CLK _20390_/D repeater278/X vssd1 vssd1 vccd1 vccd1 _20390_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_173_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11011__A1_N _21017_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19049_ _16788_/X _20820_/Q _19058_/S vssd1 vssd1 vccd1 vccd1 _19927_/D sky130_fd_sc_hd__mux2_1
XFILLER_146_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12706__B1 _11733_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10717__C1 _10677_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21011_ _21011_/CLK _21011_/D repeater235/X vssd1 vssd1 vccd1 vccd1 _21011_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12182__B2 _20345_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18639__S _18904_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13131__B1 _12922_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09704_ _21459_/Q vssd1 vssd1 vccd1 vccd1 _14528_/A sky130_fd_sc_hd__inv_2
XFILLER_74_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09635_ _21481_/Q _09632_/X _09633_/X _09634_/X vssd1 vssd1 vccd1 vccd1 _21481_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_28_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15959__B1 _15893_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_216_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13434__A1 _20474_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19245__S0 _19275_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_45_HCLK_A clkbuf_4_11_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18374__S _18910_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20726_ _21366_/CLK _20726_/D repeater254/X vssd1 vssd1 vccd1 vccd1 _20726_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_212_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13198__B1 _12991_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20657_ _20657_/CLK _20657_/D repeater197/X vssd1 vssd1 vccd1 vccd1 _20657_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12716__A _17639_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12945__B1 _12863_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10410_ _21351_/Q _10409_/Y _10395_/X _10268_/B vssd1 vssd1 vccd1 vccd1 _21351_/D
+ sky130_fd_sc_hd__o211a_1
X_11390_ _11390_/A _11390_/B _11390_/C _11390_/D vssd1 vssd1 vccd1 vccd1 _11409_/B
+ sky130_fd_sc_hd__nor4_2
X_20588_ _20946_/CLK _20588_/D repeater258/X vssd1 vssd1 vccd1 vccd1 _20588_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_109_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10341_ _20707_/Q vssd1 vssd1 vccd1 vccd1 _17545_/A sky130_fd_sc_hd__inv_2
XFILLER_192_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13060_ _13072_/A vssd1 vssd1 vccd1 vccd1 _13060_/X sky130_fd_sc_hd__buf_1
XFILLER_124_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10272_ _10272_/A _10399_/A vssd1 vssd1 vccd1 vccd1 _10273_/B sky130_fd_sc_hd__or2_2
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12011_ _12011_/A vssd1 vssd1 vccd1 vccd1 _12030_/A sky130_fd_sc_hd__inv_2
XFILLER_3_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13370__B1 _13313_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13547__A input58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21209_ _21401_/CLK _21209_/D repeater242/X vssd1 vssd1 vccd1 vccd1 _21209_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_79_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18549__S _18904_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13122__B1 _12996_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16750_ _16750_/A vssd1 vssd1 vccd1 vccd1 _16756_/A sky130_fd_sc_hd__buf_1
X_13962_ _13962_/A _13962_/B _13962_/C _13962_/D vssd1 vssd1 vccd1 vccd1 _13990_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_235_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15701_ _16012_/A vssd1 vssd1 vccd1 vccd1 _15701_/X sky130_fd_sc_hd__buf_1
X_12913_ _20728_/Q _12909_/X _12668_/X _12910_/X vssd1 vssd1 vccd1 vccd1 _20728_/D
+ sky130_fd_sc_hd__a22o_1
X_16681_ _21088_/Q _16681_/B vssd1 vssd1 vccd1 vccd1 _16681_/X sky130_fd_sc_hd__or2_1
XFILLER_74_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13893_ _13893_/A _13983_/A _13893_/C vssd1 vssd1 vccd1 vccd1 _13979_/A sky130_fd_sc_hd__or3_4
XFILLER_246_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13282__A input55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18420_ _18419_/X _20273_/Q _18904_/S vssd1 vssd1 vccd1 vccd1 _18420_/X sky130_fd_sc_hd__mux2_1
X_15632_ _15632_/A vssd1 vssd1 vccd1 vccd1 _15632_/X sky130_fd_sc_hd__buf_1
XANTENNA__21239__RESET_B repeater251/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12844_ _20756_/Q _12841_/X _09633_/X _12842_/X vssd1 vssd1 vccd1 vccd1 _20756_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09629__B1 _09628_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19236__S0 _21005_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_221_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18351_ _18036_/Y _16850_/Y _18667_/S vssd1 vssd1 vccd1 vccd1 _18351_/X sky130_fd_sc_hd__mux2_1
X_15563_ _15569_/A vssd1 vssd1 vccd1 vccd1 _15563_/X sky130_fd_sc_hd__buf_1
XPHY_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18284__S _18886_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12775_ _20794_/Q _12771_/X _09626_/X _12772_/X vssd1 vssd1 vccd1 vccd1 _20794_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_221_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18364__A1 _20762_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16593__A _16616_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_214_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17302_ _11514_/Y _17151_/X _17300_/Y _17301_/X vssd1 vssd1 vccd1 vccd1 _17302_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_70_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14514_ _20214_/Q _14513_/Y _14500_/B _14453_/X vssd1 vssd1 vccd1 vccd1 _20214_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11726_ _17387_/A _11726_/B vssd1 vssd1 vccd1 vccd1 _11735_/A sky130_fd_sc_hd__or2_2
X_18282_ _18848_/A0 _10348_/Y _18884_/S vssd1 vssd1 vccd1 vccd1 _18282_/X sky130_fd_sc_hd__mux2_1
XPHY_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15494_ _15500_/A vssd1 vssd1 vccd1 vccd1 _15494_/X sky130_fd_sc_hd__buf_1
XPHY_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17233_ _18907_/X _18019_/A _17230_/Y _17232_/X vssd1 vssd1 vccd1 vccd1 _17233_/X
+ sky130_fd_sc_hd__o22a_1
X_14445_ _21465_/Q _14351_/B _20238_/Q _14387_/Y _14444_/X vssd1 vssd1 vccd1 vccd1
+ _14449_/C sky130_fd_sc_hd__o221a_1
XPHY_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11657_ _11657_/A vssd1 vssd1 vccd1 vccd1 _11658_/A sky130_fd_sc_hd__inv_2
XPHY_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10608_ _10704_/A _20744_/Q _10659_/A _20758_/Q _10607_/X vssd1 vssd1 vccd1 vccd1
+ _10608_/X sky130_fd_sc_hd__a221o_1
XFILLER_174_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17164_ _21136_/Q vssd1 vssd1 vccd1 vccd1 _17164_/Y sky130_fd_sc_hd__inv_2
XPHY_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14376_ _14465_/B _14376_/B vssd1 vssd1 vccd1 vccd1 _14471_/A sky130_fd_sc_hd__or2_1
X_11588_ _21124_/Q _11587_/X _11583_/B vssd1 vssd1 vccd1 vccd1 _21124_/D sky130_fd_sc_hd__o21a_1
XFILLER_116_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16115_ _20329_/Q vssd1 vssd1 vccd1 vccd1 _16115_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13327_ _13327_/A _13327_/B _13327_/C vssd1 vssd1 vccd1 vccd1 _17217_/A sky130_fd_sc_hd__or3_4
XFILLER_116_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10539_ _21311_/Q vssd1 vssd1 vccd1 vccd1 _10723_/C sky130_fd_sc_hd__inv_2
X_17095_ _19694_/Q vssd1 vssd1 vccd1 vccd1 _17095_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16046_ _19511_/Q _16042_/X _16014_/X _16043_/X vssd1 vssd1 vccd1 vccd1 _19511_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_143_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13258_ _13254_/X _20563_/Q _13258_/S vssd1 vssd1 vccd1 vccd1 _20563_/D sky130_fd_sc_hd__mux2_1
XFILLER_124_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18032__B _18032_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13361__B1 _13140_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12209_ _20501_/Q vssd1 vssd1 vccd1 vccd1 _12209_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13189_ _13328_/A _17228_/A vssd1 vssd1 vccd1 vccd1 _13456_/B sky130_fd_sc_hd__or2_2
XFILLER_151_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19805_ _19820_/CLK _19805_/D vssd1 vssd1 vccd1 vccd1 _19805_/Q sky130_fd_sc_hd__dfxtp_1
X_17997_ _18147_/X _17963_/X _18160_/X _17996_/X vssd1 vssd1 vccd1 vccd1 _17997_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_111_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18459__S _18897_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16948_ _19966_/Q vssd1 vssd1 vccd1 vccd1 _16951_/A sky130_fd_sc_hd__inv_2
X_19736_ _19765_/CLK _19736_/D vssd1 vssd1 vccd1 vccd1 _19736_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09670__A _12544_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_238_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19667_ _19813_/CLK _19667_/D vssd1 vssd1 vccd1 vccd1 _19667_/Q sky130_fd_sc_hd__dfxtp_1
X_16879_ _19948_/Q _16872_/A _19949_/Q vssd1 vssd1 vccd1 vccd1 _16879_/X sky130_fd_sc_hd__o21a_1
XFILLER_92_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18618_ _18080_/Y _20663_/Q _18903_/S vssd1 vssd1 vccd1 vccd1 _18618_/X sky130_fd_sc_hd__mux2_1
XFILLER_213_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19227__S0 _20130_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19598_ _21021_/CLK _19598_/D vssd1 vssd1 vccd1 vccd1 _19598_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_240_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18194__S _18886_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18549_ _18548_/X _14080_/A _18904_/S vssd1 vssd1 vccd1 vccd1 _18549_/X sky130_fd_sc_hd__mux2_1
XFILLER_221_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20511_ _20947_/CLK _20511_/D repeater267/X vssd1 vssd1 vccd1 vccd1 _20511_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_193_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18922__S _18927_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12927__B1 _12925_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20442_ _20476_/CLK _20442_/D repeater280/X vssd1 vssd1 vccd1 vccd1 _20442_/Q sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_108_HCLK clkbuf_4_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20496_/CLK sky130_fd_sc_hd__clkbuf_16
X_20373_ _20957_/CLK _20373_/D repeater186/X vssd1 vssd1 vccd1 vccd1 _20373_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__20544__RESET_B repeater264/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18369__S _18885_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18594__A1 _12083_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21332__RESET_B repeater203/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09618_ _13108_/A _13046_/A vssd1 vssd1 vccd1 vccd1 _09672_/A sky130_fd_sc_hd__or2_2
XFILLER_18_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19218__S0 _20130_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10890_ _10890_/A vssd1 vssd1 vccd1 vccd1 _10890_/X sky130_fd_sc_hd__buf_1
XFILLER_203_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12560_ _19984_/Q vssd1 vssd1 vccd1 vccd1 _12561_/B sky130_fd_sc_hd__inv_2
XFILLER_11_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11511_ _16691_/A _11511_/B vssd1 vssd1 vccd1 vccd1 _11523_/S sky130_fd_sc_hd__or2_2
XPHY_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20709_ _21357_/CLK _20709_/D repeater210/X vssd1 vssd1 vccd1 vccd1 _20709_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12491_ _12396_/B _12493_/A _12396_/A vssd1 vssd1 vccd1 vccd1 _12492_/B sky130_fd_sc_hd__o21a_1
XANTENNA__18832__S _18928_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14230_ _20259_/Q _14004_/A _14228_/A _14174_/X vssd1 vssd1 vccd1 vccd1 _20259_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_138_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11442_ _21154_/Q _11442_/B vssd1 vssd1 vccd1 vccd1 _11443_/B sky130_fd_sc_hd__or2_1
XPHY_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13591__B1 _13509_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11373_ _11373_/A _21176_/Q _11373_/C vssd1 vssd1 vccd1 vccd1 _11376_/C sky130_fd_sc_hd__or3_4
XFILLER_166_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14161_ _20531_/Q _14071_/A _20557_/Q _14096_/A vssd1 vssd1 vccd1 vccd1 _14161_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__20285__RESET_B repeater262/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13112_ _13132_/A vssd1 vssd1 vccd1 vccd1 _13112_/X sky130_fd_sc_hd__buf_1
XANTENNA_input60_A HWDATA[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10324_ _20724_/Q vssd1 vssd1 vccd1 vccd1 _10324_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20214__RESET_B repeater202/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15332__A1 _20026_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14092_ _14092_/A _14190_/A vssd1 vssd1 vccd1 vccd1 _14093_/B sky130_fd_sc_hd__or2_2
XFILLER_79_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13343__B1 _13282_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13277__A input57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13043_ _20668_/Q _13040_/X _12879_/X _13041_/X vssd1 vssd1 vccd1 vccd1 _20668_/D
+ sky130_fd_sc_hd__a22o_1
X_17920_ _20348_/Q vssd1 vssd1 vccd1 vccd1 _17920_/Y sky130_fd_sc_hd__inv_2
X_10255_ _21348_/Q vssd1 vssd1 vccd1 vccd1 _10264_/A sky130_fd_sc_hd__inv_2
XFILLER_140_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18282__A0 _18848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_239_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17851_ _20407_/Q vssd1 vssd1 vccd1 vccd1 _17851_/Y sky130_fd_sc_hd__inv_2
X_10186_ _10157_/A _10157_/B _10185_/X _10182_/Y vssd1 vssd1 vccd1 vccd1 _21396_/D
+ sky130_fd_sc_hd__a211oi_2
X_16802_ _19930_/Q _16794_/A _19931_/Q vssd1 vssd1 vccd1 vccd1 _16802_/X sky130_fd_sc_hd__o21a_1
X_17782_ _17780_/Y _17139_/A _17781_/Y _17136_/A vssd1 vssd1 vccd1 vccd1 _17782_/X
+ sky130_fd_sc_hd__o22a_1
X_14994_ _14994_/A vssd1 vssd1 vccd1 vccd1 _14994_/Y sky130_fd_sc_hd__inv_2
XFILLER_94_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16733_ _20995_/Q _12001_/B _12002_/B vssd1 vssd1 vccd1 vccd1 _16733_/X sky130_fd_sc_hd__a21bo_1
X_19521_ _19521_/CLK _19521_/D vssd1 vssd1 vccd1 vccd1 _19521_/Q sky130_fd_sc_hd__dfxtp_1
X_13945_ _13944_/Y _13897_/A _20664_/Q _20321_/Q vssd1 vssd1 vccd1 vccd1 _13945_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_235_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19452_ _19834_/CLK _19452_/D vssd1 vssd1 vccd1 vccd1 _19452_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16664_ _21152_/Q vssd1 vssd1 vccd1 vccd1 _16664_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19209__S0 _20130_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13876_ _14016_/A _14015_/A _13876_/C _14017_/A vssd1 vssd1 vccd1 vccd1 _13877_/D
+ sky130_fd_sc_hd__or4_4
XFILLER_201_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18403_ _18402_/X _20506_/Q _18910_/S vssd1 vssd1 vccd1 vccd1 _18403_/X sky130_fd_sc_hd__mux2_1
X_15615_ _19716_/Q _15611_/X _15473_/X _15613_/X vssd1 vssd1 vccd1 vccd1 _19716_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__21002__RESET_B repeater190/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12827_ _20767_/Q _12821_/X _12658_/X _12824_/X vssd1 vssd1 vccd1 vccd1 _20767_/D
+ sky130_fd_sc_hd__a22o_1
X_19383_ _19521_/CLK _19383_/D vssd1 vssd1 vccd1 vccd1 _19383_/Q sky130_fd_sc_hd__dfxtp_1
X_16595_ _16595_/A _16595_/B vssd1 vssd1 vccd1 vccd1 _16596_/B sky130_fd_sc_hd__or2_1
XANTENNA__18337__A1 _10614_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18334_ _18031_/Y _20658_/Q _18903_/S vssd1 vssd1 vccd1 vccd1 _18334_/X sky130_fd_sc_hd__mux2_1
XANTENNA__17212__A _17212_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15546_ _15554_/A vssd1 vssd1 vccd1 vccd1 _15546_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_188_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12758_ _12783_/A vssd1 vssd1 vccd1 vccd1 _12785_/A sky130_fd_sc_hd__inv_2
XPHY_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18027__B _18027_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11709_ _21072_/Q _11704_/X _11573_/X _11705_/X vssd1 vssd1 vccd1 vccd1 _21072_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_91_HCLK_A clkbuf_4_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18265_ _18848_/A0 _14126_/Y _18902_/S vssd1 vssd1 vccd1 vccd1 _18265_/X sky130_fd_sc_hd__mux2_1
X_15477_ _15766_/A vssd1 vssd1 vccd1 vccd1 _15477_/X sky130_fd_sc_hd__buf_1
XFILLER_175_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18742__S _18880_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12689_ _20826_/Q _12686_/X _09641_/X _12688_/X vssd1 vssd1 vccd1 vccd1 _20826_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17216_ _17216_/A vssd1 vssd1 vccd1 vccd1 _17854_/A sky130_fd_sc_hd__clkbuf_2
X_14428_ _21475_/Q _14460_/D _21468_/Q _14499_/A vssd1 vssd1 vccd1 vccd1 _14428_/X
+ sky130_fd_sc_hd__o22a_1
X_18196_ _18195_/X _10606_/Y _18891_/S vssd1 vssd1 vccd1 vccd1 _18196_/X sky130_fd_sc_hd__mux2_1
X_17147_ _17376_/A vssd1 vssd1 vccd1 vccd1 _17147_/X sky130_fd_sc_hd__buf_1
XFILLER_156_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13582__B1 _13429_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14359_ _20220_/Q vssd1 vssd1 vccd1 vccd1 _14361_/C sky130_fd_sc_hd__inv_2
XFILLER_171_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09665__A input68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17078_ _20243_/Q _19876_/Q vssd1 vssd1 vccd1 vccd1 _17078_/X sky130_fd_sc_hd__and2_2
XFILLER_170_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16029_ _16029_/A vssd1 vssd1 vccd1 vccd1 _16029_/X sky130_fd_sc_hd__buf_1
XFILLER_226_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__21283__CLK _21342_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18189__S _18896_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19719_ _20326_/CLK _19719_/D vssd1 vssd1 vccd1 vccd1 _19719_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20991_ _21319_/CLK _20991_/D repeater222/X vssd1 vssd1 vccd1 vccd1 _20991_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_225_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_225_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11154__B _17169_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20796__RESET_B repeater252/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20725__RESET_B repeater264/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18652__S _18874_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21474_ _21477_/CLK _21474_/D repeater204/X vssd1 vssd1 vccd1 vccd1 _21474_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_153_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20425_ _20951_/CLK _20425_/D repeater270/X vssd1 vssd1 vccd1 vccd1 _20425_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_106_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20356_ _20980_/CLK _20356_/D repeater279/X vssd1 vssd1 vccd1 vccd1 _20356_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__13325__B1 _13171_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17792__A _21143_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20287_ _20592_/CLK _20287_/D repeater260/X vssd1 vssd1 vccd1 vccd1 _20287_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_96_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10040_ _10040_/A vssd1 vssd1 vccd1 vccd1 _10221_/C sky130_fd_sc_hd__buf_1
XFILLER_248_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19979__RESET_B repeater270/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_217_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11991_ _20985_/Q _11991_/B vssd1 vssd1 vccd1 vccd1 _11992_/B sky130_fd_sc_hd__or2_1
XFILLER_152_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18827__S _18928_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_217_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13730_ _15769_/A _15772_/A _13734_/S vssd1 vssd1 vccd1 vccd1 _20326_/D sky130_fd_sc_hd__mux2_1
XFILLER_84_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10942_ _21036_/Q vssd1 vssd1 vccd1 vccd1 _11813_/A sky130_fd_sc_hd__inv_2
XANTENNA__21006__CLK _21009_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19869__D _19869_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13661_ _13687_/A vssd1 vssd1 vccd1 vccd1 _13680_/A sky130_fd_sc_hd__clkbuf_2
X_10873_ _21263_/Q _10871_/X _09688_/X _10872_/X vssd1 vssd1 vccd1 vccd1 _21263_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_43_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13560__A input53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15400_ _15406_/A vssd1 vssd1 vccd1 vccd1 _15400_/X sky130_fd_sc_hd__buf_1
XPHY_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12612_ input14/X _11793_/X _20864_/Q _11797_/X vssd1 vssd1 vccd1 vccd1 _20864_/D
+ sky130_fd_sc_hd__o22a_1
XPHY_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16380_ _16386_/A vssd1 vssd1 vccd1 vccd1 _16380_/X sky130_fd_sc_hd__buf_1
XFILLER_25_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13592_ _20402_/Q _13588_/X _13511_/X _13589_/X vssd1 vssd1 vccd1 vccd1 _20402_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12603__A2 _12600_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15331_ _15331_/A1 _15329_/X _13553_/X _15330_/X vssd1 vssd1 vccd1 vccd1 _20027_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12543_ _12553_/A vssd1 vssd1 vccd1 vccd1 _12543_/X sky130_fd_sc_hd__buf_1
XFILLER_212_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18562__S _18748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12176__A _20361_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18050_ _18383_/X _18024_/X _18363_/X _17995_/X _18049_/X vssd1 vssd1 vccd1 vccd1
+ _18051_/C sky130_fd_sc_hd__o221a_1
X_15262_ _20484_/Q vssd1 vssd1 vccd1 vccd1 _15262_/Y sky130_fd_sc_hd__inv_2
XFILLER_157_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12474_ _12474_/A _12474_/B vssd1 vssd1 vccd1 vccd1 _12479_/A sky130_fd_sc_hd__or2_1
XFILLER_8_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17001_ _19977_/Q vssd1 vssd1 vccd1 vccd1 _17001_/Y sky130_fd_sc_hd__inv_2
X_14213_ _20270_/Q _14215_/A _14205_/X _14081_/B vssd1 vssd1 vccd1 vccd1 _20270_/D
+ sky130_fd_sc_hd__o211a_1
X_11425_ _11424_/Y _11408_/X _11413_/X _11373_/A _11414_/X vssd1 vssd1 vccd1 vccd1
+ _11426_/A sky130_fd_sc_hd__o32a_1
XFILLER_172_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15193_ _15193_/A vssd1 vssd1 vccd1 vccd1 _15193_/X sky130_fd_sc_hd__buf_2
X_14144_ _20553_/Q _14092_/A _14143_/Y _20271_/Q vssd1 vssd1 vccd1 vccd1 _14144_/X
+ sky130_fd_sc_hd__o22a_1
X_11356_ _21181_/Q vssd1 vssd1 vccd1 vccd1 _11357_/C sky130_fd_sc_hd__inv_2
XFILLER_141_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10307_ _10307_/A _10307_/B _10307_/C _10307_/D vssd1 vssd1 vccd1 vccd1 _10361_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_113_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18952_ _16656_/X _21084_/Q _18962_/S vssd1 vssd1 vccd1 vccd1 _18952_/X sky130_fd_sc_hd__mux2_1
XFILLER_180_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14075_ _14075_/A _14222_/A vssd1 vssd1 vccd1 vccd1 _14076_/B sky130_fd_sc_hd__or2_2
X_11287_ _11313_/C _11313_/B _11287_/C vssd1 vssd1 vccd1 vccd1 _11545_/A sky130_fd_sc_hd__nor3_4
X_13026_ _13040_/A vssd1 vssd1 vccd1 vccd1 _13026_/X sky130_fd_sc_hd__buf_1
X_17903_ _20411_/Q _17944_/B vssd1 vssd1 vccd1 vccd1 _17903_/Y sky130_fd_sc_hd__nand2_1
X_10238_ _21365_/Q vssd1 vssd1 vccd1 vccd1 _10280_/A sky130_fd_sc_hd__inv_2
X_18883_ _18882_/X _17186_/Y _18901_/S vssd1 vssd1 vccd1 vccd1 _18883_/X sky130_fd_sc_hd__mux2_1
X_17834_ _18930_/S _18929_/S vssd1 vssd1 vccd1 vccd1 _17852_/A sky130_fd_sc_hd__or2_4
X_10169_ _21403_/Q _21402_/Q _10169_/C vssd1 vssd1 vccd1 vccd1 _10169_/X sky130_fd_sc_hd__and3_1
XFILLER_66_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_239_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17765_ _19493_/Q vssd1 vssd1 vccd1 vccd1 _17765_/Y sky130_fd_sc_hd__inv_2
X_14977_ _14977_/A vssd1 vssd1 vccd1 vccd1 _14977_/Y sky130_fd_sc_hd__inv_2
XFILLER_207_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18737__S _18928_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19504_ _19521_/CLK _19504_/D vssd1 vssd1 vccd1 vccd1 _19504_/Q sky130_fd_sc_hd__dfxtp_1
X_16716_ _16718_/A _18935_/X vssd1 vssd1 vccd1 vccd1 _19901_/D sky130_fd_sc_hd__and2_1
X_13928_ _20636_/Q vssd1 vssd1 vccd1 vccd1 _13928_/Y sky130_fd_sc_hd__inv_2
XFILLER_235_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17696_ _19620_/Q vssd1 vssd1 vccd1 vccd1 _17696_/Y sky130_fd_sc_hd__inv_2
XFILLER_222_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16647_ _19858_/Q _15292_/B _15293_/B vssd1 vssd1 vccd1 vccd1 _16647_/X sky130_fd_sc_hd__a21bo_1
X_19435_ _21453_/CLK _19435_/D vssd1 vssd1 vccd1 vccd1 _19435_/Q sky130_fd_sc_hd__dfxtp_1
X_13859_ _20303_/Q vssd1 vssd1 vccd1 vccd1 _13972_/C sky130_fd_sc_hd__inv_2
XANTENNA__14566__A _14566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16578_ _11430_/Y _16575_/Y _16624_/A vssd1 vssd1 vccd1 vccd1 _19916_/D sky130_fd_sc_hd__o21ai_1
X_19366_ _19828_/CLK _19366_/D vssd1 vssd1 vccd1 vccd1 _19366_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18317_ _18848_/A0 _18016_/Y _18666_/S vssd1 vssd1 vccd1 vccd1 _18317_/X sky130_fd_sc_hd__mux2_1
X_15529_ _15536_/A vssd1 vssd1 vccd1 vccd1 _15529_/X sky130_fd_sc_hd__buf_1
X_19297_ _20432_/CLK _19297_/D vssd1 vssd1 vccd1 vccd1 _19297_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__18472__S _18896_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18248_ _19156_/X _20166_/Q _18249_/S vssd1 vssd1 vccd1 vccd1 _18248_/X sky130_fd_sc_hd__mux2_1
XANTENNA__20136__RESET_B repeater248/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18179_ _18848_/A0 _14129_/Y _18902_/S vssd1 vssd1 vccd1 vccd1 _18179_/X sky130_fd_sc_hd__mux2_1
X_20210_ _21477_/CLK _20210_/D repeater203/X vssd1 vssd1 vccd1 vccd1 _20210_/Q sky130_fd_sc_hd__dfrtp_1
X_21190_ _21191_/CLK _21190_/D repeater224/X vssd1 vssd1 vccd1 vccd1 _21190_/Q sky130_fd_sc_hd__dfrtp_1
X_20141_ _20142_/CLK _20141_/D repeater250/X vssd1 vssd1 vccd1 vccd1 _20141_/Q sky130_fd_sc_hd__dfrtp_1
X_09952_ _09958_/A vssd1 vssd1 vccd1 vccd1 _09952_/X sky130_fd_sc_hd__buf_1
XFILLER_89_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20072_ _20495_/CLK _20072_/D repeater276/X vssd1 vssd1 vccd1 vccd1 _20072_/Q sky130_fd_sc_hd__dfrtp_1
X_09883_ _20010_/Q _09912_/A vssd1 vssd1 vccd1 vccd1 _09884_/A sky130_fd_sc_hd__nand2_1
XFILLER_218_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18647__S _18908_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20974_ _20980_/CLK _20974_/D repeater278/X vssd1 vssd1 vccd1 vccd1 _20974_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__20977__RESET_B repeater278/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17221__B2 _17214_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20906__RESET_B repeater217/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12597__A1 _20875_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18382__S _18909_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13546__B1 _13545_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21457_ _21457_/CLK _21457_/D repeater245/X vssd1 vssd1 vccd1 vccd1 _21457_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_193_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11210_ _21211_/Q _11206_/X _09645_/X _11208_/X vssd1 vssd1 vccd1 vccd1 _21211_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_119_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12190_ _12190_/A _12190_/B _12190_/C _12190_/D vssd1 vssd1 vccd1 vccd1 _12190_/X
+ sky130_fd_sc_hd__and4_1
X_20408_ _20408_/CLK _20408_/D repeater184/X vssd1 vssd1 vccd1 vccd1 _20408_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_135_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21388_ _21390_/CLK _21388_/D repeater239/X vssd1 vssd1 vccd1 vccd1 _21388_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_107_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11141_ _15756_/B vssd1 vssd1 vccd1 vccd1 _11141_/X sky130_fd_sc_hd__buf_1
XFILLER_162_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20339_ _20422_/CLK _20339_/D repeater271/X vssd1 vssd1 vccd1 vccd1 _20339_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_89_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11072_ _21237_/Q _11072_/B vssd1 vssd1 vccd1 vccd1 _11072_/X sky130_fd_sc_hd__or2_1
Xoutput88 _17966_/Y vssd1 vssd1 vccd1 vccd1 HRDATA[18] sky130_fd_sc_hd__clkbuf_2
Xoutput99 _18076_/Y vssd1 vssd1 vccd1 vccd1 HRDATA[28] sky130_fd_sc_hd__clkbuf_2
X_10023_ _17031_/A vssd1 vssd1 vccd1 vccd1 _17038_/B sky130_fd_sc_hd__clkbuf_2
X_14900_ _20571_/Q _15002_/A _20585_/Q _14960_/B vssd1 vssd1 vccd1 vccd1 _14900_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__13555__A input55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15880_ _19592_/Q _15875_/X _15879_/X _15877_/X vssd1 vssd1 vccd1 vccd1 _19592_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_130_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input23_A HADDR[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14831_ _20101_/Q vssd1 vssd1 vccd1 vccd1 _14965_/A sky130_fd_sc_hd__inv_2
XANTENNA__18557__S _18928_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17550_ _17550_/A vssd1 vssd1 vccd1 vccd1 _17550_/X sky130_fd_sc_hd__buf_1
X_14762_ _14753_/A _14548_/X _19123_/X _20130_/Q vssd1 vssd1 vccd1 vccd1 _20130_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_16_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11974_ _13182_/B vssd1 vssd1 vccd1 vccd1 _11974_/X sky130_fd_sc_hd__buf_1
XFILLER_44_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16501_ _16509_/C vssd1 vssd1 vccd1 vccd1 _16501_/X sky130_fd_sc_hd__buf_1
XFILLER_217_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13713_ _20333_/Q _13706_/X _13712_/X _13708_/X vssd1 vssd1 vccd1 vccd1 _20333_/D
+ sky130_fd_sc_hd__a22o_1
X_17481_ _18770_/X _17324_/X _18779_/X _17480_/X vssd1 vssd1 vccd1 vccd1 _17481_/X
+ sky130_fd_sc_hd__o22a_1
X_10925_ _21202_/Q vssd1 vssd1 vccd1 vccd1 _10925_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14693_ _18249_/X _14690_/X _20166_/Q _14692_/X vssd1 vssd1 vccd1 vccd1 _20166_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_232_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19220_ _17623_/Y _17624_/Y _17625_/Y _17626_/Y _20130_/Q _20131_/Q vssd1 vssd1 vccd1
+ vccd1 _19220_/X sky130_fd_sc_hd__mux4_2
X_16432_ _19317_/Q _16427_/X _16375_/X _16428_/X vssd1 vssd1 vccd1 vccd1 _19317_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_177_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13644_ _20372_/Q _13639_/X _13586_/X _13640_/X vssd1 vssd1 vccd1 vccd1 _20372_/D
+ sky130_fd_sc_hd__a22o_1
X_10856_ _18276_/X _10853_/X _21270_/Q _10846_/X vssd1 vssd1 vccd1 vccd1 _21270_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_220_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19151_ _19147_/X _19148_/X _19149_/X _19150_/X _21018_/Q _21019_/Q vssd1 vssd1 vccd1
+ vccd1 _19151_/X sky130_fd_sc_hd__mux4_2
X_16363_ _16370_/A vssd1 vssd1 vccd1 vccd1 _16363_/X sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_repeater162_A _18880_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13575_ _13595_/A vssd1 vssd1 vccd1 vccd1 _13575_/X sky130_fd_sc_hd__buf_1
XANTENNA__18292__S _18910_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10787_ _10812_/A vssd1 vssd1 vccd1 vccd1 _10787_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_8_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18102_ _18649_/X _17858_/X _18165_/X _17211_/X _18101_/X vssd1 vssd1 vccd1 vccd1
+ _18105_/B sky130_fd_sc_hd__o221a_2
XFILLER_12_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15314_ _15314_/A vssd1 vssd1 vccd1 vccd1 _18281_/S sky130_fd_sc_hd__clkinv_4
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12526_ _12524_/X _12525_/Y _19988_/Q _11541_/A _12518_/X vssd1 vssd1 vccd1 vccd1
+ _20914_/D sky130_fd_sc_hd__a32o_1
X_19082_ _16721_/Y _20893_/Q _19908_/D vssd1 vssd1 vccd1 vccd1 _19082_/X sky130_fd_sc_hd__mux2_1
XFILLER_158_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16294_ _19391_/Q _16287_/X _16293_/X _16289_/X vssd1 vssd1 vccd1 vccd1 _19391_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_200_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18033_ _18033_/A vssd1 vssd1 vccd1 vccd1 _18078_/B sky130_fd_sc_hd__buf_4
X_15245_ _20481_/Q _15074_/A _17976_/A _20064_/Q _15244_/X vssd1 vssd1 vccd1 vccd1
+ _15250_/C sky130_fd_sc_hd__o221a_1
XFILLER_172_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12457_ _12425_/A _12425_/B _12453_/X _12455_/Y vssd1 vssd1 vccd1 vccd1 _20936_/D
+ sky130_fd_sc_hd__a211oi_2
XANTENNA_output91_A _17989_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11408_ _11408_/A vssd1 vssd1 vccd1 vccd1 _11408_/X sky130_fd_sc_hd__buf_1
X_15176_ _15176_/A vssd1 vssd1 vccd1 vccd1 _15176_/Y sky130_fd_sc_hd__inv_2
X_12388_ _12306_/A _12306_/B _12350_/A _12386_/Y vssd1 vssd1 vccd1 vccd1 _20952_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_181_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14127_ _14126_/Y _20285_/Q _20541_/Q _14080_/A vssd1 vssd1 vccd1 vccd1 _14127_/X
+ sky130_fd_sc_hd__o22a_1
X_11339_ _11374_/A _21182_/Q _21183_/Q vssd1 vssd1 vccd1 vccd1 _11340_/A sky130_fd_sc_hd__or3b_2
XFILLER_207_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19984_ _20890_/CLK _19984_/D repeater185/X vssd1 vssd1 vccd1 vccd1 _19984_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__10154__A _10154_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18935_ _16715_/X _21141_/Q _18946_/S vssd1 vssd1 vccd1 vccd1 _18935_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14058_ _20270_/Q vssd1 vssd1 vccd1 vccd1 _14080_/A sky130_fd_sc_hd__inv_2
XFILLER_67_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13009_ _20688_/Q _13005_/X _12918_/X _13007_/X vssd1 vssd1 vccd1 vccd1 _20688_/D
+ sky130_fd_sc_hd__a22o_1
X_18866_ _17256_/Y _17253_/Y _18926_/S vssd1 vssd1 vccd1 vccd1 _18866_/X sky130_fd_sc_hd__mux2_1
XFILLER_227_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17817_ _17854_/A vssd1 vssd1 vccd1 vccd1 _17817_/X sky130_fd_sc_hd__buf_1
XANTENNA__18467__S _18896_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18797_ _18796_/X _17423_/Y _18927_/S vssd1 vssd1 vccd1 vccd1 _18797_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17748_ _19509_/Q vssd1 vssd1 vccd1 vccd1 _17748_/Y sky130_fd_sc_hd__inv_2
XFILLER_223_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20388__RESET_B repeater278/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17679_ _19780_/Q vssd1 vssd1 vccd1 vccd1 _17679_/Y sky130_fd_sc_hd__inv_2
XFILLER_223_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18951__A1 _21085_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12809__A _16342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19418_ _19835_/CLK _19418_/D vssd1 vssd1 vccd1 vccd1 _19418_/Q sky130_fd_sc_hd__dfxtp_1
X_20690_ _20693_/CLK _20690_/D repeater194/X vssd1 vssd1 vccd1 vccd1 _20690_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__20317__RESET_B repeater262/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19349_ _20137_/CLK _19349_/D vssd1 vssd1 vccd1 vccd1 _19349_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18703__A1 _19211_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17911__C1 _17910_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21311_ _21341_/CLK _21311_/D repeater201/X vssd1 vssd1 vccd1 vccd1 _21311_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_163_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12544__A _12544_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18930__S _18930_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16016__A _16016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18467__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21242_ _21242_/CLK _21242_/D repeater189/X vssd1 vssd1 vccd1 vccd1 _21242_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_105_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21176__RESET_B repeater216/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21173_ _21184_/CLK _21173_/D repeater220/X vssd1 vssd1 vccd1 vccd1 _21173_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_117_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20124_ _21273_/CLK _20124_/D repeater246/X vssd1 vssd1 vccd1 vccd1 _20124_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_77_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09935_ _13327_/A vssd1 vssd1 vccd1 vccd1 _13188_/A sky130_fd_sc_hd__buf_2
XFILLER_104_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20055_ _20066_/CLK _20055_/D repeater281/X vssd1 vssd1 vccd1 vccd1 _20055_/Q sky130_fd_sc_hd__dfrtp_2
X_09866_ _20034_/Q _10843_/B vssd1 vssd1 vccd1 vccd1 _09867_/A sky130_fd_sc_hd__nor2_1
XFILLER_85_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18377__S _18879_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09797_ _09804_/C vssd1 vssd1 vccd1 vccd1 _09806_/B sky130_fd_sc_hd__buf_1
XFILLER_218_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15453__B1 _15450_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater160 _18841_/S vssd1 vssd1 vccd1 vccd1 _18850_/S sky130_fd_sc_hd__buf_8
XFILLER_234_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater171 _18891_/S vssd1 vssd1 vccd1 vccd1 _18897_/S sky130_fd_sc_hd__buf_8
XPHY_4303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater182 _20121_/Q vssd1 vssd1 vccd1 vccd1 _19280_/S0 sky130_fd_sc_hd__clkbuf_16
XPHY_4314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater193 repeater194/X vssd1 vssd1 vccd1 vccd1 repeater193/X sky130_fd_sc_hd__clkbuf_8
XPHY_4336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20740__RESET_B repeater207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20957_ _20957_/CLK _20957_/D repeater187/X vssd1 vssd1 vccd1 vccd1 _20957_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_3635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10710_ _10708_/A _10708_/B _10677_/A _10708_/Y vssd1 vssd1 vccd1 vccd1 _21320_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_242_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20058__RESET_B repeater281/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11690_ _11690_/A vssd1 vssd1 vccd1 vccd1 _11690_/X sky130_fd_sc_hd__buf_1
XPHY_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20888_ _21444_/CLK _20888_/D repeater247/X vssd1 vssd1 vccd1 vccd1 _20888_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10641_ _10754_/B vssd1 vssd1 vccd1 vccd1 _10694_/A sky130_fd_sc_hd__buf_1
XPHY_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19001__S _19019_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13360_ _13378_/A vssd1 vssd1 vccd1 vccd1 _13360_/X sky130_fd_sc_hd__buf_1
XFILLER_220_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10572_ _10662_/A _10661_/A _10664_/A _10663_/A vssd1 vssd1 vccd1 vccd1 _10573_/C
+ sky130_fd_sc_hd__or4_4
XFILLER_158_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12990__A1 _20696_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12311_ _12311_/A _12380_/A vssd1 vssd1 vccd1 vccd1 _12312_/B sky130_fd_sc_hd__or2_2
XFILLER_10_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13519__B1 _13454_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13291_ _20551_/Q _13286_/X _13211_/X _13288_/X vssd1 vssd1 vccd1 vccd1 _20551_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18840__S _18885_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18458__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15030_ _20072_/Q vssd1 vssd1 vccd1 vccd1 _15086_/A sky130_fd_sc_hd__inv_2
X_12242_ _20926_/Q _12239_/Y _12474_/A _20506_/Q _12241_/X vssd1 vssd1 vccd1 vccd1
+ _12255_/B sky130_fd_sc_hd__o221a_1
XFILLER_174_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12173_ _12081_/X _20342_/Q _12097_/X _20340_/Q vssd1 vssd1 vccd1 vccd1 _12173_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19994__RESET_B repeater220/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11124_ _21006_/Q vssd1 vssd1 vccd1 vccd1 _11124_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16981_ _19971_/Q _16970_/A _16965_/A _19972_/Q vssd1 vssd1 vccd1 vccd1 _16981_/X
+ sky130_fd_sc_hd__o31a_1
X_18720_ _18719_/X _14443_/Y _18897_/S vssd1 vssd1 vccd1 vccd1 _18720_/X sky130_fd_sc_hd__mux2_1
X_11055_ _11055_/A _11098_/A vssd1 vssd1 vccd1 vccd1 _11096_/B sky130_fd_sc_hd__nor2_1
X_15932_ _19566_/Q _15927_/X _15795_/X _15928_/X vssd1 vssd1 vccd1 vccd1 _19566_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_190_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10006_ _10003_/Y _17033_/A _21416_/Q _10005_/A vssd1 vssd1 vccd1 vccd1 _10006_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_236_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15863_ _16093_/A _16150_/B _16419_/C vssd1 vssd1 vccd1 vccd1 _15875_/A sky130_fd_sc_hd__or3_4
X_18651_ _18650_/X _16875_/Y _18886_/S vssd1 vssd1 vccd1 vccd1 _18651_/X sky130_fd_sc_hd__mux2_1
XANTENNA__18287__S _18617_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20828__RESET_B repeater251/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14247__B2 _18946_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17602_ _19297_/Q vssd1 vssd1 vccd1 vccd1 _17602_/Y sky130_fd_sc_hd__inv_2
X_14814_ _14819_/A vssd1 vssd1 vccd1 vccd1 _14818_/S sky130_fd_sc_hd__clkbuf_2
X_15794_ _19631_/Q _15787_/X _15793_/X _15789_/X vssd1 vssd1 vccd1 vccd1 _19631_/D
+ sky130_fd_sc_hd__a22o_1
X_18582_ _18845_/A0 _10336_/Y _18884_/S vssd1 vssd1 vccd1 vccd1 _18582_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14745_ _14747_/A _14541_/A _15833_/B vssd1 vssd1 vccd1 vccd1 _14745_/X sky130_fd_sc_hd__o21a_1
X_17533_ _19313_/Q _17533_/B vssd1 vssd1 vccd1 vccd1 _17533_/Y sky130_fd_sc_hd__nand2_1
XFILLER_33_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11957_ _19109_/X _11128_/X _11956_/X vssd1 vssd1 vccd1 vccd1 _21004_/D sky130_fd_sc_hd__a21oi_1
XANTENNA__18933__A1 _21143_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19281__S1 _20124_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17464_ _21130_/Q vssd1 vssd1 vccd1 vccd1 _17464_/Y sky130_fd_sc_hd__inv_2
X_10908_ _10908_/A _10908_/B _17060_/C vssd1 vssd1 vccd1 vccd1 _10910_/S sky130_fd_sc_hd__or3_4
XANTENNA__20410__RESET_B repeater185/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14676_ _10918_/B _14674_/X _14679_/B vssd1 vssd1 vccd1 vccd1 _14676_/Y sky130_fd_sc_hd__a21oi_2
X_11888_ _21023_/Q _11887_/X _21023_/Q _11887_/X vssd1 vssd1 vccd1 vccd1 _21023_/D
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_199_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16415_ _19328_/Q _16413_/X _16207_/X _16414_/X vssd1 vssd1 vccd1 vccd1 _19328_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_20_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19203_ _17742_/Y _17743_/Y _17744_/Y _17745_/Y _19275_/S0 _21004_/Q vssd1 vssd1
+ vccd1 vccd1 _19203_/X sky130_fd_sc_hd__mux4_2
X_13627_ _20383_/Q _13625_/X _13482_/X _13626_/X vssd1 vssd1 vccd1 vccd1 _20383_/D
+ sky130_fd_sc_hd__a22o_1
X_10839_ _10839_/A vssd1 vssd1 vccd1 vccd1 _10839_/Y sky130_fd_sc_hd__inv_2
X_17395_ _18823_/X vssd1 vssd1 vccd1 vccd1 _17395_/Y sky130_fd_sc_hd__inv_2
XFILLER_220_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18697__A0 _18696_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09938__A _13188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19134_ _19687_/Q _19375_/Q _19671_/Q _19663_/Q _19285_/S0 _21017_/Q vssd1 vssd1
+ vccd1 vccd1 _19134_/X sky130_fd_sc_hd__mux4_1
X_16346_ _16352_/A vssd1 vssd1 vccd1 vccd1 _16353_/A sky130_fd_sc_hd__inv_2
X_13558_ _20421_/Q _13549_/X _13557_/X _13551_/X vssd1 vssd1 vccd1 vccd1 _20421_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_200_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18035__B _18078_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12509_ _12498_/Y _16609_/A _11316_/X _11280_/A _12512_/A vssd1 vssd1 vccd1 vccd1
+ _12510_/A sky130_fd_sc_hd__o32a_1
X_19065_ _21186_/Q _21128_/Q _19910_/Q vssd1 vssd1 vccd1 vccd1 _19065_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16277_ _20331_/Q vssd1 vssd1 vccd1 vccd1 _16277_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_157_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13489_ input45/X vssd1 vssd1 vccd1 vccd1 _13489_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__18750__S _18850_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18449__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15228_ _20479_/Q _15099_/X _17896_/A _20058_/Q _15227_/X vssd1 vssd1 vccd1 vccd1
+ _15232_/C sky130_fd_sc_hd__o221a_1
X_18016_ _20834_/Q vssd1 vssd1 vccd1 vccd1 _18016_/Y sky130_fd_sc_hd__inv_2
XFILLER_173_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_141_HCLK clkbuf_4_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _21238_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_clkbuf_leaf_146_HCLK_A clkbuf_opt_1_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19110__A1 _11916_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15159_ _15185_/A vssd1 vssd1 vccd1 vccd1 _15177_/A sky130_fd_sc_hd__buf_1
XFILLER_5_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09673__A _15329_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19967_ _20413_/CLK _19967_/D repeater184/X vssd1 vssd1 vccd1 vccd1 _19967_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__15683__B1 _15585_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09720_ _21235_/Q vssd1 vssd1 vccd1 vccd1 _11060_/A sky130_fd_sc_hd__inv_2
XANTENNA__13195__A _13217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18918_ _18917_/X _21250_/Q _20870_/Q vssd1 vssd1 vccd1 vccd1 _18918_/X sky130_fd_sc_hd__mux2_1
XFILLER_234_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19898_ _21193_/CLK _19898_/D repeater224/X vssd1 vssd1 vccd1 vccd1 _19898_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_228_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09651_ input41/X vssd1 vssd1 vccd1 vccd1 _12857_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_228_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18849_ _18848_/X _13942_/Y _18849_/S vssd1 vssd1 vccd1 vccd1 _18849_/X sky130_fd_sc_hd__mux2_1
XANTENNA__18197__S _18617_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_216_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20811_ _21379_/CLK _20811_/D repeater213/X vssd1 vssd1 vccd1 vccd1 _20811_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_36_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18924__A1 _14313_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18925__S _18930_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19272__S1 _21004_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20742_ _21319_/CLK _20742_/D repeater191/X vssd1 vssd1 vccd1 vccd1 _20742_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20151__RESET_B repeater250/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20673_ _21294_/CLK _20673_/D repeater209/X vssd1 vssd1 vccd1 vccd1 _20673_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18660__S _18875_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21225_ _21235_/CLK _21225_/D repeater249/X vssd1 vssd1 vccd1 vccd1 _21225_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_104_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21156_ _21429_/CLK _21156_/D repeater229/X vssd1 vssd1 vccd1 vccd1 _21156_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_104_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20107_ _20107_/CLK _20107_/D repeater259/X vssd1 vssd1 vccd1 vccd1 _20107_/Q sky130_fd_sc_hd__dfrtp_4
X_09918_ _21121_/Q vssd1 vssd1 vccd1 vccd1 _11591_/A sky130_fd_sc_hd__buf_1
X_21087_ _21087_/CLK _21087_/D repeater228/X vssd1 vssd1 vccd1 vccd1 _21087_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_144_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20038_ _21183_/CLK _20038_/D repeater216/X vssd1 vssd1 vccd1 vccd1 _20038_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_218_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09849_ _09861_/B _09864_/A vssd1 vssd1 vccd1 vccd1 _09849_/X sky130_fd_sc_hd__or2_1
XFILLER_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15426__B1 _15424_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12860_ _12860_/A vssd1 vssd1 vccd1 vccd1 _12860_/X sky130_fd_sc_hd__clkbuf_4
XPHY_4100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11811_ _11811_/A _11837_/A vssd1 vssd1 vccd1 vccd1 _11832_/A sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_22_HCLK clkbuf_4_3_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _21255_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_4144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12791_ _12803_/A vssd1 vssd1 vccd1 vccd1 _12791_/X sky130_fd_sc_hd__buf_1
XPHY_4155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18835__S _18835_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19263__S1 _21004_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14530_ _20208_/Q _16618_/A _14530_/C vssd1 vssd1 vccd1 vccd1 _15832_/C sky130_fd_sc_hd__or3_4
XFILLER_14_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11742_ _21057_/Q _11735_/X _11741_/X _11737_/X vssd1 vssd1 vccd1 vccd1 _21057_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14461_ _14461_/A _14461_/B _14461_/C _14461_/D vssd1 vssd1 vccd1 vccd1 _14462_/D
+ sky130_fd_sc_hd__or4_4
XPHY_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11673_ _21089_/Q vssd1 vssd1 vccd1 vccd1 _17046_/A sky130_fd_sc_hd__inv_2
XPHY_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16200_ _21452_/Q vssd1 vssd1 vccd1 vccd1 _16200_/X sky130_fd_sc_hd__buf_1
XPHY_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18679__A0 _17281_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13412_ _20484_/Q _13410_/X _13216_/X _13411_/X vssd1 vssd1 vccd1 vccd1 _20484_/D
+ sky130_fd_sc_hd__a22o_1
X_10624_ _21321_/Q _20749_/Q _10551_/C _10623_/Y vssd1 vssd1 vccd1 vccd1 _10624_/X
+ sky130_fd_sc_hd__o22a_1
X_17180_ _20564_/Q _17187_/B vssd1 vssd1 vccd1 vccd1 _17180_/Y sky130_fd_sc_hd__nor2_1
XPHY_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14392_ _20026_/Q vssd1 vssd1 vccd1 vccd1 _14392_/Y sky130_fd_sc_hd__inv_2
XPHY_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_164_HCLK clkbuf_opt_0_HCLK/A vssd1 vssd1 vccd1 vccd1 _21444_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_139_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16131_ _21453_/Q vssd1 vssd1 vccd1 vccd1 _16131_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13343_ _20523_/Q _13339_/X _13282_/X _13340_/X vssd1 vssd1 vccd1 vccd1 _20523_/D
+ sky130_fd_sc_hd__a22o_1
X_10555_ _21331_/Q vssd1 vssd1 vccd1 vccd1 _10660_/A sky130_fd_sc_hd__inv_2
XFILLER_154_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18570__S _18617_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19757__CLK _19765_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21027__RESET_B repeater242/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16062_ _21222_/Q vssd1 vssd1 vccd1 vccd1 _16247_/A sky130_fd_sc_hd__buf_1
X_13274_ input58/X vssd1 vssd1 vccd1 vccd1 _13274_/X sky130_fd_sc_hd__buf_2
X_10486_ _21302_/Q vssd1 vssd1 vccd1 vccd1 _10778_/A sky130_fd_sc_hd__inv_2
X_15013_ _20083_/Q _15012_/Y _15004_/B _14952_/X vssd1 vssd1 vccd1 vccd1 _20083_/D
+ sky130_fd_sc_hd__o211a_1
X_12225_ _12473_/A _20505_/Q _20925_/Q _12221_/Y _12224_/X vssd1 vssd1 vccd1 vccd1
+ _12232_/C sky130_fd_sc_hd__o221a_1
XANTENNA__13912__B1 _13911_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18851__A0 _17079_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19821_ _19821_/CLK _19821_/D vssd1 vssd1 vccd1 vccd1 _19821_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12156_ _12309_/A _20337_/Q _12093_/X _20344_/Q _12155_/X vssd1 vssd1 vccd1 vccd1
+ _12156_/X sky130_fd_sc_hd__o221a_1
XFILLER_123_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11107_ _11107_/A vssd1 vssd1 vccd1 vccd1 _21229_/D sky130_fd_sc_hd__inv_2
X_19752_ _19765_/CLK _19752_/D vssd1 vssd1 vccd1 vccd1 _19752_/Q sky130_fd_sc_hd__dfxtp_1
X_16964_ _16979_/B vssd1 vssd1 vccd1 vccd1 _16965_/A sky130_fd_sc_hd__clkbuf_2
X_12087_ _12087_/A _12087_/B _12087_/C _12087_/D vssd1 vssd1 vccd1 vccd1 _12087_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_238_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18703_ _17704_/Y _19211_/X _18930_/S vssd1 vssd1 vccd1 vccd1 _18703_/X sky130_fd_sc_hd__mux2_2
X_11038_ _19971_/Q _19970_/Q _19972_/Q vssd1 vssd1 vccd1 vccd1 _16979_/A sky130_fd_sc_hd__or3_1
X_15915_ _19575_/Q _15911_/X _15881_/X _15912_/X vssd1 vssd1 vccd1 vccd1 _19575_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_110_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19683_ _19811_/CLK _19683_/D vssd1 vssd1 vccd1 vccd1 _19683_/Q sky130_fd_sc_hd__dfxtp_1
X_16895_ _19953_/Q vssd1 vssd1 vccd1 vccd1 _16895_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18634_ _18845_/A0 _10454_/Y _18896_/S vssd1 vssd1 vccd1 vccd1 _18634_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15846_ _19606_/Q _15841_/X _15812_/X _15842_/X vssd1 vssd1 vccd1 vccd1 _19606_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_237_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09647__A1 _21477_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18565_ _17079_/Y _15260_/Y _18908_/S vssd1 vssd1 vccd1 vccd1 _18565_/X sky130_fd_sc_hd__mux2_1
XANTENNA__18745__S _18775_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12359__A _12359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15777_ _19638_/Q _15768_/X _15776_/X _15770_/X vssd1 vssd1 vccd1 vccd1 _19638_/D
+ sky130_fd_sc_hd__a22o_1
X_12989_ input61/X vssd1 vssd1 vccd1 vccd1 _12989_/X sky130_fd_sc_hd__buf_2
XFILLER_18_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19254__S1 _21004_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_1_0_HCLK clkbuf_4_1_0_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_opt_1_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_221_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17516_ _19578_/Q vssd1 vssd1 vccd1 vccd1 _17516_/Y sky130_fd_sc_hd__inv_2
XFILLER_178_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14728_ _20144_/Q _14723_/X _13714_/X _14724_/X vssd1 vssd1 vccd1 vccd1 _20144_/D
+ sky130_fd_sc_hd__a22o_1
X_18496_ _17079_/Y _12062_/Y _18908_/S vssd1 vssd1 vccd1 vccd1 _18496_/X sky130_fd_sc_hd__mux2_1
XFILLER_205_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_232_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14659_ _14659_/A _14659_/B vssd1 vssd1 vccd1 vccd1 _14660_/A sky130_fd_sc_hd__nand2_1
X_17447_ _19312_/Q _17631_/B vssd1 vssd1 vccd1 vccd1 _17447_/Y sky130_fd_sc_hd__nor2_1
XFILLER_21_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09668__A input67/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17378_ _17378_/A vssd1 vssd1 vccd1 vccd1 _17378_/X sky130_fd_sc_hd__buf_1
XFILLER_174_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19117_ _19116_/S _11123_/Y _19117_/S vssd1 vssd1 vccd1 vccd1 _19117_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10414__C1 _10375_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21450__RESET_B repeater247/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16329_ _19373_/Q _16326_/X _16231_/X _16328_/X vssd1 vssd1 vccd1 vccd1 _19373_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_119_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18480__S _18904_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19048_ _16792_/X _20821_/Q _19058_/S vssd1 vssd1 vccd1 vccd1 _19928_/D sky130_fd_sc_hd__mux2_1
XFILLER_161_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18842__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19190__S0 _19280_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21010_ _21431_/CLK _21010_/D repeater238/X vssd1 vssd1 vccd1 vccd1 _21010_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_59_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09703_ _21463_/Q _09690_/X _09702_/X _09694_/X vssd1 vssd1 vccd1 vccd1 _21463_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_68_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_45_HCLK clkbuf_4_11_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _21193_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_67_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09634_ _09660_/A vssd1 vssd1 vccd1 vccd1 _09634_/X sky130_fd_sc_hd__buf_1
XANTENNA__11693__A1 _21081_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_215_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18655__S _18787_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19245__S1 _21004_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_231_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20725_ _21366_/CLK _20725_/D repeater264/X vssd1 vssd1 vccd1 vccd1 _20725_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_211_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13198__A1 _20594_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20656_ _20657_/CLK _20656_/D repeater197/X vssd1 vssd1 vccd1 vccd1 _20656_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_137_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18390__S _18908_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20587_ _20947_/CLK _20587_/D repeater258/X vssd1 vssd1 vccd1 vccd1 _20587_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_99_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10340_ _10340_/A _10340_/B _10340_/C _10340_/D vssd1 vssd1 vccd1 vccd1 _10361_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_137_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15895__B1 _15785_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10271_ _10271_/A _10271_/B vssd1 vssd1 vccd1 vccd1 _10399_/A sky130_fd_sc_hd__or2_1
XFILLER_2_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12010_ _12029_/A vssd1 vssd1 vccd1 vccd1 _12010_/X sky130_fd_sc_hd__buf_1
XANTENNA__19181__S0 _20123_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21208_ _21401_/CLK _21208_/D repeater256/X vssd1 vssd1 vccd1 vccd1 _21208_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_79_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21139_ _21147_/CLK _21139_/D repeater215/X vssd1 vssd1 vccd1 vccd1 _21139_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_48_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13961_ _13950_/X _13961_/B _13961_/C _13961_/D vssd1 vssd1 vccd1 vccd1 _13962_/D
+ sky130_fd_sc_hd__and4b_1
XFILLER_59_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15700_ input60/X vssd1 vssd1 vccd1 vccd1 _16012_/A sky130_fd_sc_hd__clkbuf_2
X_12912_ _20729_/Q _12909_/X _12666_/X _12910_/X vssd1 vssd1 vccd1 vccd1 _20729_/D
+ sky130_fd_sc_hd__a22o_1
X_16680_ _20001_/Q _16680_/B vssd1 vssd1 vccd1 vccd1 _18947_/S sky130_fd_sc_hd__nor2_1
XANTENNA__20073__RESET_B repeater276/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13892_ _20317_/Q vssd1 vssd1 vccd1 vccd1 _13893_/C sky130_fd_sc_hd__inv_2
XFILLER_219_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20002__RESET_B repeater220/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12843_ _20757_/Q _12841_/X _09630_/X _12842_/X vssd1 vssd1 vccd1 vccd1 _20757_/D
+ sky130_fd_sc_hd__a22o_1
X_15631_ _19706_/Q _15625_/X _15582_/X _15627_/X vssd1 vssd1 vccd1 vccd1 _19706_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12179__A _20345_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18565__S _18908_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19236__S1 _21006_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_234_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15562_ _15568_/A vssd1 vssd1 vccd1 vccd1 _15569_/A sky130_fd_sc_hd__inv_2
X_18350_ _18349_/X _10282_/A _18886_/S vssd1 vssd1 vccd1 vccd1 _18350_/X sky130_fd_sc_hd__mux2_1
X_12774_ _20795_/Q _12771_/X _09621_/X _12772_/X vssd1 vssd1 vccd1 vccd1 _20795_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14513_ _14513_/A vssd1 vssd1 vccd1 vccd1 _14513_/Y sky130_fd_sc_hd__inv_2
XPHY_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17301_ _17301_/A vssd1 vssd1 vccd1 vccd1 _17301_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__20287__CLK _20592_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_214_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21279__RESET_B repeater207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11725_ _21064_/Q _11720_/X _11573_/X _11721_/X vssd1 vssd1 vccd1 vccd1 _21064_/D
+ sky130_fd_sc_hd__a22o_1
X_18281_ _19196_/X _21276_/Q _18281_/S vssd1 vssd1 vccd1 vccd1 _18281_/X sky130_fd_sc_hd__mux2_1
X_15493_ _15499_/A vssd1 vssd1 vccd1 vccd1 _15500_/A sky130_fd_sc_hd__inv_2
XFILLER_70_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14444_ _20237_/Q _14442_/Y _14443_/Y _20214_/Q vssd1 vssd1 vccd1 vccd1 _14444_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_147_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17232_ _17474_/A vssd1 vssd1 vccd1 vccd1 _17232_/X sky130_fd_sc_hd__buf_2
XPHY_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11656_ _11667_/B vssd1 vssd1 vccd1 vccd1 _11657_/A sky130_fd_sc_hd__clkbuf_2
XPHY_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10607_ _21329_/Q _20757_/Q _10658_/A _10606_/Y vssd1 vssd1 vccd1 vccd1 _10607_/X
+ sky130_fd_sc_hd__o22a_1
X_17163_ _17160_/Y _17175_/B _17161_/Y _17177_/B _17162_/X vssd1 vssd1 vccd1 vccd1
+ _17163_/X sky130_fd_sc_hd__o221a_1
XPHY_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14375_ _14463_/C _14476_/A vssd1 vssd1 vccd1 vccd1 _14376_/B sky130_fd_sc_hd__or2_2
XPHY_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_repeater242_A repeater250/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11587_ _21123_/Q _21122_/Q _11596_/B vssd1 vssd1 vccd1 vccd1 _11587_/X sky130_fd_sc_hd__and3_1
XFILLER_10_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16114_ _19476_/Q _16108_/X _16113_/X _16111_/X vssd1 vssd1 vccd1 vccd1 _19476_/D
+ sky130_fd_sc_hd__a22o_1
X_13326_ _20530_/Q _13321_/X _13173_/X _13322_/X vssd1 vssd1 vccd1 vccd1 _20530_/D
+ sky130_fd_sc_hd__a22o_1
X_10538_ _21312_/Q vssd1 vssd1 vccd1 vccd1 _10540_/B sky130_fd_sc_hd__inv_2
XFILLER_171_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17094_ _19638_/Q vssd1 vssd1 vccd1 vccd1 _17094_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16045_ _19512_/Q _16042_/X _16012_/X _16043_/X vssd1 vssd1 vccd1 vccd1 _19512_/D
+ sky130_fd_sc_hd__a22o_1
X_13257_ _17087_/A _13259_/B vssd1 vssd1 vccd1 vccd1 _13258_/S sky130_fd_sc_hd__or2_1
X_10469_ _10763_/A _20676_/Q _10773_/A _20686_/Q vssd1 vssd1 vccd1 vccd1 _10469_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__19172__S0 _19280_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12208_ _20946_/Q vssd1 vssd1 vccd1 vccd1 _12395_/A sky130_fd_sc_hd__inv_2
XFILLER_124_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13188_ _13188_/A _13327_/B _13188_/C vssd1 vssd1 vccd1 vccd1 _17228_/A sky130_fd_sc_hd__or3_4
XFILLER_69_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19804_ _19820_/CLK _19804_/D vssd1 vssd1 vccd1 vccd1 _19804_/Q sky130_fd_sc_hd__dfxtp_1
X_12139_ _12313_/B vssd1 vssd1 vccd1 vccd1 _12139_/X sky130_fd_sc_hd__buf_1
XFILLER_215_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17996_ _18065_/A vssd1 vssd1 vccd1 vccd1 _17996_/X sky130_fd_sc_hd__buf_1
XANTENNA_clkbuf_leaf_51_HCLK_A clkbuf_4_11_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09951__A _09957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19735_ _19765_/CLK _19735_/D vssd1 vssd1 vccd1 vccd1 _19735_/Q sky130_fd_sc_hd__dfxtp_1
X_16947_ _16951_/B _16946_/X _16939_/X vssd1 vssd1 vccd1 vccd1 _16947_/X sky130_fd_sc_hd__o21a_1
XFILLER_96_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13473__A _13483_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21062__CLK _21134_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19666_ _19812_/CLK _19666_/D vssd1 vssd1 vccd1 vccd1 _19666_/Q sky130_fd_sc_hd__dfxtp_1
X_16878_ _19949_/Q vssd1 vssd1 vccd1 vccd1 _16878_/Y sky130_fd_sc_hd__inv_2
XFILLER_225_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18617_ _18616_/X _21306_/Q _18617_/S vssd1 vssd1 vccd1 vccd1 _18617_/X sky130_fd_sc_hd__mux2_2
X_15829_ _19614_/Q _15824_/X _15812_/X _15825_/X vssd1 vssd1 vccd1 vccd1 _19614_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_64_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19227__S1 _20131_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19597_ _21040_/CLK _19597_/D vssd1 vssd1 vccd1 vccd1 _19597_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18475__S _18884_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_213_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18548_ _18547_/X _13903_/Y _18903_/S vssd1 vssd1 vccd1 vccd1 _18548_/X sky130_fd_sc_hd__mux2_1
XFILLER_178_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18479_ _18478_/X _13957_/Y _18903_/S vssd1 vssd1 vccd1 vccd1 _18479_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_221_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20510_ _20929_/CLK _20510_/D repeater267/X vssd1 vssd1 vccd1 vccd1 _20510_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_20_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20441_ _20476_/CLK _20441_/D repeater280/X vssd1 vssd1 vccd1 vccd1 _20441_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_118_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20372_ _20957_/CLK _20372_/D repeater186/X vssd1 vssd1 vccd1 vccd1 _20372_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__15847__B _15847_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19163__S0 _19280_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15629__B1 _15548_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20513__RESET_B repeater267/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14301__B1 _20122_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13383__A _13383_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09617_ _11182_/A _12898_/A vssd1 vssd1 vccd1 vccd1 _13046_/A sky130_fd_sc_hd__or2_4
XANTENNA__18385__S _18909_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19218__S1 _20131_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_243_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21372__RESET_B repeater257/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12727__A _13329_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11510_ _20251_/Q vssd1 vssd1 vccd1 vccd1 _16691_/A sky130_fd_sc_hd__inv_2
XPHY_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21301__RESET_B repeater208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20708_ _21357_/CLK _20708_/D repeater210/X vssd1 vssd1 vccd1 vccd1 _20708_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_12_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12490_ _12490_/A _12490_/B _12490_/C vssd1 vssd1 vccd1 vccd1 _12493_/A sky130_fd_sc_hd__or3_4
XFILLER_211_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11441_ _21153_/Q _21152_/Q vssd1 vssd1 vccd1 vccd1 _11442_/B sky130_fd_sc_hd__or2_1
XPHY_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20639_ _20657_/CLK _20639_/D repeater198/X vssd1 vssd1 vccd1 vccd1 _20639_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_7_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14160_ _20539_/Q vssd1 vssd1 vccd1 vccd1 _14160_/Y sky130_fd_sc_hd__inv_2
X_11372_ _21177_/Q vssd1 vssd1 vccd1 vccd1 _11373_/A sky130_fd_sc_hd__inv_2
XFILLER_50_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13111_ _13138_/A vssd1 vssd1 vccd1 vccd1 _13132_/A sky130_fd_sc_hd__buf_1
XFILLER_125_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10323_ _10311_/X _10323_/B _10323_/C _10323_/D vssd1 vssd1 vccd1 vccd1 _10361_/B
+ sky130_fd_sc_hd__and4b_1
XFILLER_166_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14091_ _14091_/A _14091_/B vssd1 vssd1 vccd1 vccd1 _14190_/A sky130_fd_sc_hd__or2_1
XFILLER_180_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19154__S0 _19285_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13042_ _20669_/Q _13040_/X _12875_/X _13041_/X vssd1 vssd1 vccd1 vccd1 _20669_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_input53_A HWDATA[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10254_ _21349_/Q vssd1 vssd1 vccd1 vccd1 _10265_/A sky130_fd_sc_hd__inv_2
XFILLER_78_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17850_ _20821_/Q vssd1 vssd1 vccd1 vccd1 _17850_/Y sky130_fd_sc_hd__inv_2
X_10185_ _10185_/A vssd1 vssd1 vccd1 vccd1 _10185_/X sky130_fd_sc_hd__buf_2
XFILLER_120_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_239_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16801_ _16801_/A vssd1 vssd1 vccd1 vccd1 _16801_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17781_ _21079_/Q vssd1 vssd1 vccd1 vccd1 _17781_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14993_ _14962_/B _14868_/B _14991_/Y _14989_/X vssd1 vssd1 vccd1 vccd1 _20090_/D
+ sky130_fd_sc_hd__a211oi_2
X_19520_ _19521_/CLK _19520_/D vssd1 vssd1 vccd1 vccd1 _19520_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_247_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16732_ _20994_/Q _12000_/B _12001_/B vssd1 vssd1 vccd1 vccd1 _16732_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__12854__B1 _12853_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13944_ _20664_/Q vssd1 vssd1 vccd1 vccd1 _13944_/Y sky130_fd_sc_hd__inv_2
XFILLER_235_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16045__B1 _16012_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19451_ _19834_/CLK _19451_/D vssd1 vssd1 vccd1 vccd1 _19451_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_235_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16663_ _16663_/A _18949_/X vssd1 vssd1 vccd1 vccd1 _19865_/D sky130_fd_sc_hd__and2_1
X_13875_ _13875_/A vssd1 vssd1 vccd1 vccd1 _14017_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_repeater192_A repeater212/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18295__S _18680_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19209__S1 _20131_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18402_ _17806_/Y _20340_/Q _18874_/S vssd1 vssd1 vccd1 vccd1 _18402_/X sky130_fd_sc_hd__mux2_1
XFILLER_201_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12826_ _20768_/Q _12821_/X _12656_/X _12824_/X vssd1 vssd1 vccd1 vccd1 _20768_/D
+ sky130_fd_sc_hd__a22o_1
X_15614_ _19717_/Q _15611_/X _15469_/X _15613_/X vssd1 vssd1 vccd1 vccd1 _19717_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_222_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19382_ _19521_/CLK _19382_/D vssd1 vssd1 vccd1 vccd1 _19382_/Q sky130_fd_sc_hd__dfxtp_1
X_16594_ _16594_/A _16594_/B vssd1 vssd1 vccd1 vccd1 _16594_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__20922__CLK _20930_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18333_ _18332_/X _16858_/A _18667_/S vssd1 vssd1 vccd1 vccd1 _18333_/X sky130_fd_sc_hd__mux2_1
XFILLER_203_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15545_ _15553_/A vssd1 vssd1 vccd1 vccd1 _15554_/A sky130_fd_sc_hd__inv_2
X_12757_ _12777_/A vssd1 vssd1 vccd1 vccd1 _12757_/X sky130_fd_sc_hd__buf_1
XPHY_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11708_ _21073_/Q _11704_/X _11571_/X _11705_/X vssd1 vssd1 vccd1 vccd1 _21073_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10632__A2 _10631_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15476_ _19779_/Q _15468_/X _15475_/X _15471_/X vssd1 vssd1 vccd1 vccd1 _19779_/D
+ sky130_fd_sc_hd__a22o_1
X_18264_ _18263_/X _14094_/A _18904_/S vssd1 vssd1 vccd1 vccd1 _18264_/X sky130_fd_sc_hd__mux2_2
X_12688_ _12708_/A vssd1 vssd1 vccd1 vccd1 _12688_/X sky130_fd_sc_hd__buf_1
XPHY_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14427_ _21470_/Q vssd1 vssd1 vccd1 vccd1 _14427_/Y sky130_fd_sc_hd__inv_2
X_17215_ _17315_/A vssd1 vssd1 vccd1 vccd1 _17216_/A sky130_fd_sc_hd__buf_1
XANTENNA__13031__B1 _13030_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11639_ _11641_/A vssd1 vssd1 vccd1 vccd1 _11640_/A sky130_fd_sc_hd__buf_1
X_18195_ _18845_/A0 _10430_/Y _18896_/S vssd1 vssd1 vccd1 vccd1 _18195_/X sky130_fd_sc_hd__mux2_1
XPHY_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14358_ _20217_/Q vssd1 vssd1 vccd1 vccd1 _14502_/A sky130_fd_sc_hd__inv_2
X_17146_ _17290_/A vssd1 vssd1 vccd1 vccd1 _17376_/A sky130_fd_sc_hd__buf_1
XFILLER_128_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15859__B1 _15791_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13309_ _20541_/Q _13307_/X _13151_/X _13308_/X vssd1 vssd1 vccd1 vccd1 _20541_/D
+ sky130_fd_sc_hd__a22o_1
X_17077_ _17075_/Y _19885_/Q _12506_/X _17076_/X vssd1 vssd1 vccd1 vccd1 _19882_/D
+ sky130_fd_sc_hd__a31o_1
X_14289_ _20125_/Q vssd1 vssd1 vccd1 vccd1 _15335_/B sky130_fd_sc_hd__buf_1
XANTENNA__19145__S0 _19285_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16028_ _16028_/A vssd1 vssd1 vccd1 vccd1 _16028_/X sky130_fd_sc_hd__buf_1
XFILLER_112_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16779__A _16779_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17979_ _18079_/A vssd1 vssd1 vccd1 vccd1 _18033_/A sky130_fd_sc_hd__buf_1
XANTENNA__18025__A1 _18350_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19718_ _19774_/CLK _19718_/D vssd1 vssd1 vccd1 vccd1 _19718_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_242_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12845__B1 _09636_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20990_ _21319_/CLK _20990_/D repeater222/X vssd1 vssd1 vccd1 vccd1 _20990_/Q sky130_fd_sc_hd__dfrtp_1
X_19649_ _21021_/CLK _19649_/D vssd1 vssd1 vccd1 vccd1 _19649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18933__S _18946_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_221_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19860__RESET_B repeater226/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21473_ _21477_/CLK _21473_/D repeater204/X vssd1 vssd1 vccd1 vccd1 _21473_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__13022__B1 _12849_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20424_ _20951_/CLK _20424_/D repeater271/X vssd1 vssd1 vccd1 vccd1 _20424_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_135_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20765__RESET_B repeater211/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20355_ _20972_/CLK _20355_/D repeater280/X vssd1 vssd1 vccd1 vccd1 _20355_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20286_ _20286_/CLK _20286_/D repeater262/X vssd1 vssd1 vccd1 vccd1 _20286_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_48_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13089__B1 _12863_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10530__A _20699_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11990_ _20984_/Q _20983_/Q vssd1 vssd1 vccd1 vccd1 _11991_/B sky130_fd_sc_hd__or2_1
XFILLER_152_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10941_ _21209_/Q vssd1 vssd1 vccd1 vccd1 _10941_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19004__S _19019_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13660_ _13685_/A vssd1 vssd1 vccd1 vccd1 _13687_/A sky130_fd_sc_hd__inv_2
XFILLER_44_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10872_ _10872_/A vssd1 vssd1 vccd1 vccd1 _10872_/X sky130_fd_sc_hd__buf_1
XFILLER_220_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12611_ input15/X _11793_/X _20865_/Q _11797_/X vssd1 vssd1 vccd1 vccd1 _20865_/D
+ sky130_fd_sc_hd__o22a_1
XPHY_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13591_ _20403_/Q _13588_/X _13509_/X _13589_/X vssd1 vssd1 vccd1 vccd1 _20403_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_197_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18843__S _18891_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17527__B1 _20119_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15330_ _15330_/A vssd1 vssd1 vccd1 vccd1 _15330_/X sky130_fd_sc_hd__buf_1
XPHY_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12542_ _17286_/A _14273_/D vssd1 vssd1 vccd1 vccd1 _12553_/A sky130_fd_sc_hd__or2_2
XFILLER_12_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15261_ _20471_/Q vssd1 vssd1 vccd1 vccd1 _15261_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12473_ _12473_/A _12483_/A vssd1 vssd1 vccd1 vccd1 _12474_/B sky130_fd_sc_hd__or2_1
X_17000_ _16998_/Y _16999_/Y _16984_/X vssd1 vssd1 vccd1 vccd1 _17000_/X sky130_fd_sc_hd__o21a_1
X_14212_ _14212_/A vssd1 vssd1 vccd1 vccd1 _14215_/A sky130_fd_sc_hd__inv_2
X_11424_ _19914_/Q vssd1 vssd1 vccd1 vccd1 _11424_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15192_ _20059_/Q _15191_/Y _15185_/X _15074_/B vssd1 vssd1 vccd1 vccd1 _20059_/D
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_3_5_0_HCLK clkbuf_3_5_0_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_137_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14143_ _20542_/Q vssd1 vssd1 vccd1 vccd1 _14143_/Y sky130_fd_sc_hd__inv_2
X_11355_ _11410_/C _11409_/C vssd1 vssd1 vccd1 vccd1 _16632_/C sky130_fd_sc_hd__nor2_2
XFILLER_153_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20435__RESET_B repeater278/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19127__S0 _19285_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10306_ _10267_/A _20710_/Q _21349_/Q _10303_/Y _10305_/X vssd1 vssd1 vccd1 vccd1
+ _10307_/D sky130_fd_sc_hd__o221a_1
X_18951_ _16658_/X _21085_/Q _18962_/S vssd1 vssd1 vccd1 vccd1 _18951_/X sky130_fd_sc_hd__mux2_1
X_14074_ _14074_/A _14074_/B vssd1 vssd1 vccd1 vccd1 _14222_/A sky130_fd_sc_hd__or2_1
X_11286_ _11300_/A _20912_/Q _11286_/C _12505_/A vssd1 vssd1 vccd1 vccd1 _11287_/C
+ sky130_fd_sc_hd__or4_4
XFILLER_141_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17902_ _20825_/Q _17944_/B vssd1 vssd1 vccd1 vccd1 _17902_/Y sky130_fd_sc_hd__nand2_1
X_13025_ _20678_/Q _13019_/X _12857_/X _13021_/X vssd1 vssd1 vccd1 vccd1 _20678_/D
+ sky130_fd_sc_hd__a22o_1
X_10237_ _21366_/Q vssd1 vssd1 vccd1 vccd1 _10281_/A sky130_fd_sc_hd__inv_2
XANTENNA__12920__A input51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18882_ _18881_/X _10527_/Y _18910_/S vssd1 vssd1 vccd1 vccd1 _18882_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17833_ _18615_/X _17227_/X _18290_/X _17817_/X vssd1 vssd1 vccd1 vccd1 _17833_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_239_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10168_ _10168_/A _10168_/B vssd1 vssd1 vccd1 vccd1 _10169_/C sky130_fd_sc_hd__nor2_1
XFILLER_120_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12827__B1 _12658_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17764_ _19581_/Q vssd1 vssd1 vccd1 vccd1 _17764_/Y sky130_fd_sc_hd__inv_2
X_14976_ _14965_/B _14878_/B _14972_/Y _14975_/X vssd1 vssd1 vccd1 vccd1 _20100_/D
+ sky130_fd_sc_hd__a211oi_2
X_10099_ _20791_/Q vssd1 vssd1 vccd1 vccd1 _10099_/Y sky130_fd_sc_hd__inv_2
XFILLER_212_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19503_ _19521_/CLK _19503_/D vssd1 vssd1 vccd1 vccd1 _19503_/Q sky130_fd_sc_hd__dfxtp_1
X_16715_ _19901_/Q _14241_/B _14242_/B vssd1 vssd1 vccd1 vccd1 _16715_/X sky130_fd_sc_hd__a21bo_1
XFILLER_81_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13927_ _13925_/Y _20300_/Q _20643_/Q _14016_/A _13926_/X vssd1 vssd1 vccd1 vccd1
+ _13930_/C sky130_fd_sc_hd__o221a_1
X_17695_ _19436_/Q vssd1 vssd1 vccd1 vccd1 _17695_/Y sky130_fd_sc_hd__inv_2
XFILLER_207_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19434_ _19626_/CLK _19434_/D vssd1 vssd1 vccd1 vccd1 _19434_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16646_ _16652_/A _18957_/X vssd1 vssd1 vccd1 vccd1 _19857_/D sky130_fd_sc_hd__and2_1
XFILLER_179_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13858_ _20304_/Q vssd1 vssd1 vccd1 vccd1 _13971_/D sky130_fd_sc_hd__inv_2
XFILLER_204_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12809_ _16342_/A vssd1 vssd1 vccd1 vccd1 _12809_/X sky130_fd_sc_hd__clkbuf_2
X_19365_ _21001_/CLK _19365_/D vssd1 vssd1 vccd1 vccd1 _19365_/Q sky130_fd_sc_hd__dfxtp_1
X_16577_ _11749_/A _16576_/X _16519_/Y _16516_/A vssd1 vssd1 vccd1 vccd1 _16624_/A
+ sky130_fd_sc_hd__a211o_1
XANTENNA__18753__S _18909_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13252__B1 _13171_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13789_ _20614_/Q vssd1 vssd1 vccd1 vccd1 _13789_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18316_ _18315_/X _20589_/Q _18907_/S vssd1 vssd1 vccd1 vccd1 _18316_/X sky130_fd_sc_hd__mux2_1
X_15528_ _15528_/A _15542_/B _16311_/C vssd1 vssd1 vccd1 vccd1 _15536_/A sky130_fd_sc_hd__or3_4
X_19296_ _20432_/CLK _19296_/D vssd1 vssd1 vccd1 vccd1 _19296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13004__B1 _13003_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18247_ _19151_/X _20165_/Q _18249_/S vssd1 vssd1 vccd1 vccd1 _18247_/X sky130_fd_sc_hd__mux2_1
X_15459_ _15459_/A vssd1 vssd1 vccd1 vccd1 _15459_/X sky130_fd_sc_hd__buf_1
XFILLER_117_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09676__A _12548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18178_ _18177_/X _14583_/A _18898_/S vssd1 vssd1 vccd1 vccd1 _18178_/X sky130_fd_sc_hd__mux2_1
XFILLER_143_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17129_ _19462_/Q vssd1 vssd1 vccd1 vccd1 _17129_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20176__RESET_B repeater200/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09951_ _09957_/A vssd1 vssd1 vccd1 vccd1 _09958_/A sky130_fd_sc_hd__inv_2
X_20140_ _20142_/CLK _20140_/D repeater250/X vssd1 vssd1 vccd1 vccd1 _20140_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__20105__RESET_B repeater259/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20071_ _20075_/CLK _20071_/D repeater276/X vssd1 vssd1 vccd1 vccd1 _20071_/Q sky130_fd_sc_hd__dfrtp_2
X_09882_ _20006_/Q _20007_/Q _20008_/Q _20009_/Q vssd1 vssd1 vccd1 vccd1 _09912_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_131_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12830__A _12842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18928__S _18928_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_239_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20973_ _20982_/CLK _20973_/D repeater187/X vssd1 vssd1 vccd1 vccd1 _20973_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_54_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18663__S _18906_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15588__A _15588_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21456_ _21461_/CLK _21456_/D repeater245/X vssd1 vssd1 vccd1 vccd1 _21456_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__11557__B1 _10889_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20407_ _20408_/CLK _20407_/D repeater184/X vssd1 vssd1 vccd1 vccd1 _20407_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_162_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21387_ _21390_/CLK _21387_/D repeater252/X vssd1 vssd1 vccd1 vccd1 _21387_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_162_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11140_ _21221_/Q vssd1 vssd1 vccd1 vccd1 _15756_/B sky130_fd_sc_hd__buf_1
X_20338_ _20951_/CLK _20338_/D repeater271/X vssd1 vssd1 vccd1 vccd1 _20338_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_123_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11071_ _11071_/A vssd1 vssd1 vccd1 vccd1 _11072_/B sky130_fd_sc_hd__inv_2
X_20269_ _20293_/CLK _20269_/D repeater263/X vssd1 vssd1 vccd1 vccd1 _20269_/Q sky130_fd_sc_hd__dfrtp_1
Xoutput89 _17973_/Y vssd1 vssd1 vccd1 vccd1 HRDATA[19] sky130_fd_sc_hd__clkbuf_2
X_10022_ _21411_/Q _14813_/D _11614_/B vssd1 vssd1 vccd1 vccd1 _21411_/D sky130_fd_sc_hd__a21o_1
XFILLER_248_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18838__S _18880_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_236_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14830_ _20102_/Q vssd1 vssd1 vccd1 vccd1 _14880_/A sky130_fd_sc_hd__inv_2
XFILLER_56_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input16_A HADDR[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14761_ _19123_/X _14758_/B _14760_/X vssd1 vssd1 vccd1 vccd1 _20131_/D sky130_fd_sc_hd__a21oi_1
XFILLER_63_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11973_ _11973_/A vssd1 vssd1 vccd1 vccd1 _13175_/A sky130_fd_sc_hd__buf_1
X_16500_ _21053_/Q _21052_/Q _21054_/Q vssd1 vssd1 vccd1 vccd1 _16509_/C sky130_fd_sc_hd__or3_1
XFILLER_17_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13712_ _15429_/A vssd1 vssd1 vccd1 vccd1 _13712_/X sky130_fd_sc_hd__clkbuf_4
X_10924_ _21201_/Q _21028_/Q _10922_/Y _11805_/A vssd1 vssd1 vccd1 vccd1 _10931_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_232_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17480_ _17928_/A vssd1 vssd1 vccd1 vccd1 _17480_/X sky130_fd_sc_hd__buf_1
X_14692_ _14692_/A vssd1 vssd1 vccd1 vccd1 _14692_/X sky130_fd_sc_hd__buf_1
XFILLER_232_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16431_ _19318_/Q _16427_/X _15881_/A _16428_/X vssd1 vssd1 vccd1 vccd1 _19318_/D
+ sky130_fd_sc_hd__a22o_1
X_10855_ _18277_/X _10853_/X _21271_/Q _10846_/X vssd1 vssd1 vccd1 vccd1 _21271_/D
+ sky130_fd_sc_hd__o22a_1
X_13643_ _20373_/Q _13639_/X _13584_/X _13640_/X vssd1 vssd1 vccd1 vccd1 _20373_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18573__S _18928_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19150_ _19658_/Q _19650_/Q _19634_/Q _19818_/Q _19285_/S0 _21017_/Q vssd1 vssd1
+ vccd1 vccd1 _19150_/X sky130_fd_sc_hd__mux4_2
X_16362_ _16405_/A _16419_/B _16377_/C vssd1 vssd1 vccd1 vccd1 _16370_/A sky130_fd_sc_hd__or3_4
X_13574_ _13574_/A vssd1 vssd1 vccd1 vccd1 _13595_/A sky130_fd_sc_hd__clkbuf_2
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10786_ _10830_/A vssd1 vssd1 vccd1 vccd1 _10812_/A sky130_fd_sc_hd__clkbuf_2
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18101_ _18144_/X _17205_/X _18168_/X _17861_/A vssd1 vssd1 vccd1 vccd1 _18101_/X
+ sky130_fd_sc_hd__o22a_2
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12525_ _16564_/A _12525_/B _12525_/C vssd1 vssd1 vccd1 vccd1 _12525_/Y sky130_fd_sc_hd__nor3_4
X_15313_ _13600_/X _20035_/Q _15313_/S vssd1 vssd1 vccd1 vccd1 _20035_/D sky130_fd_sc_hd__mux2_1
X_19081_ _16722_/X _20894_/Q _19908_/D vssd1 vssd1 vccd1 vccd1 _19081_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16293_ _20325_/Q vssd1 vssd1 vccd1 vccd1 _16293_/X sky130_fd_sc_hd__clkbuf_2
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_repeater155_A _18875_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18032_ _18032_/A _18032_/B vssd1 vssd1 vccd1 vccd1 _18032_/Y sky130_fd_sc_hd__nor2_1
XFILLER_172_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15244_ _20478_/Q _15071_/A _15243_/Y _20047_/Q vssd1 vssd1 vccd1 vccd1 _15244_/X
+ sky130_fd_sc_hd__o22a_1
X_12456_ _20937_/Q _12455_/Y _12448_/X _12427_/B vssd1 vssd1 vccd1 vccd1 _20937_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__14734__B1 _13704_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11548__A0 _21135_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11407_ _19915_/Q vssd1 vssd1 vccd1 vccd1 _11407_/Y sky130_fd_sc_hd__inv_2
X_15175_ _15104_/X _15082_/B _15173_/Y _15201_/B vssd1 vssd1 vccd1 vccd1 _20068_/D
+ sky130_fd_sc_hd__a211oi_2
X_12387_ _20953_/Q _12386_/Y _12373_/X _12308_/B vssd1 vssd1 vccd1 vccd1 _20953_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_207_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output84_A _17911_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14126_ _20556_/Q vssd1 vssd1 vccd1 vccd1 _14126_/Y sky130_fd_sc_hd__inv_2
X_11338_ _21181_/Q _11357_/D vssd1 vssd1 vccd1 vccd1 _11374_/A sky130_fd_sc_hd__or2_1
XFILLER_140_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19983_ _20890_/CLK _19983_/D repeater185/X vssd1 vssd1 vccd1 vccd1 _19983_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_4_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18934_ _16717_/X _21142_/Q _18946_/S vssd1 vssd1 vccd1 vccd1 _18934_/X sky130_fd_sc_hd__mux2_1
X_14057_ _20271_/Q vssd1 vssd1 vccd1 vccd1 _14081_/A sky130_fd_sc_hd__inv_2
X_11269_ _20910_/Q _11313_/B _12505_/A vssd1 vssd1 vccd1 vccd1 _11271_/C sky130_fd_sc_hd__or3_1
XANTENNA__16239__B1 _16006_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13008_ _20689_/Q _13005_/X _13006_/X _13007_/X vssd1 vssd1 vccd1 vccd1 _20689_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_140_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18865_ _18864_/X _19261_/X _18930_/S vssd1 vssd1 vccd1 vccd1 _18865_/X sky130_fd_sc_hd__mux2_2
XFILLER_228_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18748__S _18748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17816_ _20405_/Q _17944_/B vssd1 vssd1 vccd1 vccd1 _17816_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__15961__A _15961_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__21404__RESET_B repeater252/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18796_ _17427_/Y _17425_/X _18926_/S vssd1 vssd1 vccd1 vccd1 _18796_/X sky130_fd_sc_hd__mux2_1
XFILLER_208_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17747_ _19389_/Q vssd1 vssd1 vccd1 vccd1 _17747_/Y sky130_fd_sc_hd__inv_2
X_14959_ _20105_/Q _14967_/A _14958_/X _14883_/B vssd1 vssd1 vccd1 vccd1 _20105_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__13481__A _13481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_106_HCLK_A clkbuf_4_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17678_ _19716_/Q vssd1 vssd1 vccd1 vccd1 _17678_/Y sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_169_HCLK_A clkbuf_opt_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19417_ _19784_/CLK _19417_/D vssd1 vssd1 vccd1 vccd1 _19417_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_223_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16629_ _20250_/Q vssd1 vssd1 vccd1 vccd1 _16631_/A sky130_fd_sc_hd__inv_2
XANTENNA__18483__S _18904_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_2_0_HCLK_A clkbuf_3_3_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11236__C1 _19910_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19348_ _21453_/CLK _19348_/D vssd1 vssd1 vccd1 vccd1 _19348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19279_ _19733_/Q _19373_/Q _19789_/Q _19773_/Q _19280_/S0 _20122_/Q vssd1 vssd1
+ vccd1 vccd1 _19279_/X sky130_fd_sc_hd__mux4_1
XFILLER_248_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21310_ _21338_/CLK _21310_/D repeater222/X vssd1 vssd1 vccd1 vccd1 _21310_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__14725__B1 _13707_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11539__B1 _10900_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21241_ _21433_/CLK _21241_/D repeater236/X vssd1 vssd1 vccd1 vccd1 _21241_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_190_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21172_ _21182_/CLK _21172_/D repeater216/X vssd1 vssd1 vccd1 vccd1 _21172_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_105_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20123_ _21273_/CLK _20123_/D repeater246/X vssd1 vssd1 vccd1 vccd1 _20123_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__18219__A1 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09934_ _20890_/Q vssd1 vssd1 vccd1 vccd1 _13327_/A sky130_fd_sc_hd__buf_1
XANTENNA__15574__C _15574_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20054_ _20480_/CLK _20054_/D repeater183/X vssd1 vssd1 vccd1 vccd1 _20054_/Q sky130_fd_sc_hd__dfrtp_1
X_09865_ _09859_/A _09864_/X _09859_/Y vssd1 vssd1 vccd1 vccd1 _21443_/D sky130_fd_sc_hd__a21oi_1
XANTENNA_input8_A HADDR[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18658__S _18748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09796_ _09780_/A _09783_/A input74/X _09795_/Y vssd1 vssd1 vccd1 vccd1 _09804_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_133_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater150 _18884_/S vssd1 vssd1 vccd1 vccd1 _18908_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_246_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater161 _18617_/S vssd1 vssd1 vccd1 vccd1 _18841_/S sky130_fd_sc_hd__buf_8
Xrepeater172 _18775_/S vssd1 vssd1 vccd1 vccd1 _18891_/S sky130_fd_sc_hd__buf_6
XPHY_4304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater183 repeater280/X vssd1 vssd1 vccd1 vccd1 repeater183/X sky130_fd_sc_hd__buf_8
XFILLER_45_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13464__B1 _13272_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater194 repeater196/X vssd1 vssd1 vccd1 vccd1 repeater194/X sky130_fd_sc_hd__buf_4
XPHY_4326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20956_ _20981_/CLK _20956_/D repeater187/X vssd1 vssd1 vccd1 vccd1 _20956_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_4359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20887_ _21444_/CLK _20887_/D repeater246/X vssd1 vssd1 vccd1 vccd1 _20887_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__18393__S _18902_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_242_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13767__A1 _20601_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10640_ _10685_/A vssd1 vssd1 vccd1 vccd1 _10754_/B sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_28_HCLK_A clkbuf_4_9_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10571_ _21334_/Q vssd1 vssd1 vccd1 vccd1 _10663_/A sky130_fd_sc_hd__inv_2
XFILLER_42_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20098__RESET_B repeater259/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12310_ _12310_/A _12310_/B vssd1 vssd1 vccd1 vccd1 _12380_/A sky130_fd_sc_hd__or2_1
XFILLER_158_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14716__B1 _13586_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13290_ _20552_/Q _13286_/X _13209_/X _13288_/X vssd1 vssd1 vccd1 vccd1 _20552_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_213_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12241_ _20942_/Q _20522_/Q _20942_/Q _20522_/Q vssd1 vssd1 vccd1 vccd1 _12241_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_21439_ _21459_/CLK _21439_/D repeater245/X vssd1 vssd1 vccd1 vccd1 _21439_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_135_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12172_ _20357_/Q vssd1 vssd1 vccd1 vccd1 _12172_/Y sky130_fd_sc_hd__inv_2
XFILLER_122_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13566__A _13566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11123_ _21223_/Q vssd1 vssd1 vccd1 vccd1 _11123_/Y sky130_fd_sc_hd__inv_2
XFILLER_123_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16980_ _16980_/A vssd1 vssd1 vccd1 vccd1 _16980_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11054_ _11054_/A _11104_/A vssd1 vssd1 vccd1 vccd1 _11098_/A sky130_fd_sc_hd__or2_1
X_15931_ _19567_/Q _15927_/X _15793_/X _15928_/X vssd1 vssd1 vccd1 vccd1 _19567_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_110_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18568__S _18896_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10005_ _10005_/A vssd1 vssd1 vccd1 vccd1 _17033_/A sky130_fd_sc_hd__inv_2
XFILLER_77_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18650_ _18848_/A0 _18091_/Y _18666_/S vssd1 vssd1 vccd1 vccd1 _18650_/X sky130_fd_sc_hd__mux2_1
XFILLER_209_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15862_ _16405_/B vssd1 vssd1 vccd1 vccd1 _16150_/B sky130_fd_sc_hd__buf_1
XFILLER_236_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19963__RESET_B repeater185/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17601_ _19779_/Q vssd1 vssd1 vccd1 vccd1 _17601_/Y sky130_fd_sc_hd__inv_2
X_14813_ _21411_/Q _14813_/B _14813_/C _14813_/D vssd1 vssd1 vccd1 vccd1 _14819_/A
+ sky130_fd_sc_hd__or4_4
X_18581_ _18580_/X _14576_/A _18748_/S vssd1 vssd1 vccd1 vccd1 _18581_/X sky130_fd_sc_hd__mux2_2
XFILLER_18_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13455__B1 _13454_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output122_A _17061_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15793_ _15793_/A vssd1 vssd1 vccd1 vccd1 _15793_/X sky130_fd_sc_hd__buf_2
XFILLER_17_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17532_ _19337_/Q vssd1 vssd1 vccd1 vccd1 _17532_/Y sky130_fd_sc_hd__inv_2
X_14744_ _14744_/A vssd1 vssd1 vccd1 vccd1 _14747_/A sky130_fd_sc_hd__buf_1
X_11956_ _11951_/A _11136_/X _11127_/A vssd1 vssd1 vccd1 vccd1 _11956_/X sky130_fd_sc_hd__o21a_1
XANTENNA__20868__RESET_B repeater247/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17463_ _21139_/Q vssd1 vssd1 vccd1 vccd1 _17463_/Y sky130_fd_sc_hd__inv_2
X_10907_ _18993_/X _09919_/B _21248_/Q _17026_/B vssd1 vssd1 vccd1 vccd1 _21248_/D
+ sky130_fd_sc_hd__o22a_1
XANTENNA_repeater272_A repeater278/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11887_ _11874_/Y _11889_/B _11886_/A _19115_/S _11886_/Y vssd1 vssd1 vccd1 vccd1
+ _11887_/X sky130_fd_sc_hd__a32o_1
X_14675_ _10985_/A _14674_/X _14673_/Y vssd1 vssd1 vccd1 vccd1 _14679_/B sky130_fd_sc_hd__o21a_1
X_19202_ _17738_/Y _17739_/Y _17740_/Y _17741_/Y _19275_/S0 _21004_/Q vssd1 vssd1
+ vccd1 vccd1 _19202_/X sky130_fd_sc_hd__mux4_2
X_16414_ _16414_/A vssd1 vssd1 vccd1 vccd1 _16414_/X sky130_fd_sc_hd__buf_1
XFILLER_232_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10838_ _10756_/A _10756_/B _10827_/X _10836_/Y vssd1 vssd1 vccd1 vccd1 _21279_/D
+ sky130_fd_sc_hd__a211oi_2
X_13626_ _13626_/A vssd1 vssd1 vccd1 vccd1 _13626_/X sky130_fd_sc_hd__buf_1
X_17394_ _18824_/X vssd1 vssd1 vccd1 vccd1 _17394_/Y sky130_fd_sc_hd__inv_2
XFILLER_158_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19133_ _19759_/Q _19751_/Q _19743_/Q _19735_/Q _19285_/S0 _21017_/Q vssd1 vssd1
+ vccd1 vccd1 _19133_/X sky130_fd_sc_hd__mux4_2
X_16345_ _16352_/A vssd1 vssd1 vccd1 vccd1 _16345_/X sky130_fd_sc_hd__buf_1
X_10769_ _10769_/A _10769_/B vssd1 vssd1 vccd1 vccd1 _10811_/A sky130_fd_sc_hd__or2_1
X_13557_ input54/X vssd1 vssd1 vccd1 vccd1 _13557_/X sky130_fd_sc_hd__buf_4
XANTENNA__09938__B _10859_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12645__A _14304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12508_ _11545_/X _12525_/B _12507_/X _19908_/Q _19882_/Q vssd1 vssd1 vccd1 vccd1
+ _12512_/A sky130_fd_sc_hd__o32a_1
X_19064_ _21187_/Q _21129_/Q _19910_/Q vssd1 vssd1 vccd1 vccd1 _19064_/X sky130_fd_sc_hd__mux2_1
XANTENNA__14707__B1 _12849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13488_ _20450_/Q _13481_/X _13487_/X _13483_/X vssd1 vssd1 vccd1 vccd1 _20450_/D
+ sky130_fd_sc_hd__a22o_1
X_16276_ _16287_/A vssd1 vssd1 vccd1 vccd1 _16276_/X sky130_fd_sc_hd__buf_1
XFILLER_173_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18015_ _20456_/Q vssd1 vssd1 vccd1 vccd1 _18015_/Y sky130_fd_sc_hd__inv_2
X_15227_ _15226_/Y _20054_/Q _20475_/Q _15068_/A vssd1 vssd1 vccd1 vccd1 _15227_/X
+ sky130_fd_sc_hd__o22a_1
X_12439_ _20946_/Q _12437_/X _12438_/X _12434_/A vssd1 vssd1 vccd1 vccd1 _20946_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_172_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13179__C input73/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15158_ _15158_/A _15158_/B _15144_/X _15157_/X vssd1 vssd1 vccd1 vccd1 _15185_/A
+ sky130_fd_sc_hd__or4bb_4
XFILLER_153_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18051__B _18051_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14109_ _20544_/Q vssd1 vssd1 vccd1 vccd1 _17897_/A sky130_fd_sc_hd__inv_2
X_19966_ _20413_/CLK _19966_/D repeater185/X vssd1 vssd1 vccd1 vccd1 _19966_/Q sky130_fd_sc_hd__dfrtp_1
X_15089_ _15089_/A vssd1 vssd1 vccd1 vccd1 _15089_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18917_ _21431_/Q _21240_/Q _20871_/Q vssd1 vssd1 vccd1 vccd1 _18917_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19897_ _21185_/CLK _19897_/D repeater222/X vssd1 vssd1 vccd1 vccd1 _19897_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_67_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18478__S _18884_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09650_ _21476_/Q _09643_/X _09649_/X _09646_/X vssd1 vssd1 vccd1 vccd1 _21476_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_67_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18621__A1 _10631_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18848_ _18848_/A0 _14167_/Y _18902_/S vssd1 vssd1 vccd1 vccd1 _18848_/X sky130_fd_sc_hd__mux2_1
XFILLER_228_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18779_ _18778_/X _14569_/A _18898_/S vssd1 vssd1 vccd1 vccd1 _18779_/X sky130_fd_sc_hd__mux2_2
XFILLER_243_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20810_ _21242_/CLK _20810_/D repeater189/X vssd1 vssd1 vccd1 vccd1 _20810_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_63_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20741_ _21306_/CLK _20741_/D repeater207/X vssd1 vssd1 vccd1 vccd1 _20741_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20538__RESET_B repeater267/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19102__S _19870_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20672_ _21294_/CLK _20672_/D repeater209/X vssd1 vssd1 vccd1 vccd1 _20672_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_23_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20191__RESET_B repeater200/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18941__S _18946_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_opt_3_HCLK clkbuf_opt_3_HCLK/A vssd1 vssd1 vccd1 vccd1 _19985_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__20120__RESET_B repeater248/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15371__B1 _15355_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19559__CLK _19706_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21224_ _21235_/CLK _21224_/D repeater249/X vssd1 vssd1 vccd1 vccd1 _21224_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_117_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13386__A _13456_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21155_ _21429_/CLK _21155_/D repeater229/X vssd1 vssd1 vccd1 vccd1 _21155_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_160_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17663__A2 _17856_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20106_ _20107_/CLK _20106_/D repeater259/X vssd1 vssd1 vccd1 vccd1 _20106_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_104_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09917_ _11584_/B vssd1 vssd1 vccd1 vccd1 _09919_/B sky130_fd_sc_hd__buf_1
XFILLER_132_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21086_ _21087_/CLK _21086_/D repeater228/X vssd1 vssd1 vccd1 vccd1 _21086_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA__18388__S _18906_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20037_ _21183_/CLK _20037_/D repeater216/X vssd1 vssd1 vccd1 vccd1 _20037_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__18073__C1 _18072_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09848_ _14530_/C _10843_/C vssd1 vssd1 vccd1 vccd1 _09864_/A sky130_fd_sc_hd__or2_1
XFILLER_218_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09779_ _09775_/A _09777_/X _09781_/B _09778_/Y vssd1 vssd1 vccd1 vccd1 _21461_/D
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_46_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_233_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ _11810_/A _11841_/A vssd1 vssd1 vccd1 vccd1 _11837_/A sky130_fd_sc_hd__or2_1
XPHY_4134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12790_ _20785_/Q _12784_/X _09652_/X _12786_/X vssd1 vssd1 vccd1 vccd1 _20785_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20961__RESET_B repeater187/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11741_ _13171_/A vssd1 vssd1 vccd1 vccd1 _11741_/X sky130_fd_sc_hd__clkbuf_2
XPHY_4178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20939_ _20950_/CLK _20939_/D repeater278/X vssd1 vssd1 vccd1 vccd1 _20939_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_4189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20279__RESET_B repeater263/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19012__S _19019_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_152_HCLK_A clkbuf_opt_1_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14460_ _14460_/A _14460_/B _14460_/C _14460_/D vssd1 vssd1 vccd1 vccd1 _14462_/C
+ sky130_fd_sc_hd__or4_4
X_11672_ _11672_/A vssd1 vssd1 vccd1 vccd1 _21090_/D sky130_fd_sc_hd__inv_2
XANTENNA__18128__A0 _17079_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20208__RESET_B repeater248/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10623_ _20749_/Q vssd1 vssd1 vccd1 vccd1 _10623_/Y sky130_fd_sc_hd__inv_2
X_13411_ _13411_/A vssd1 vssd1 vccd1 vccd1 _13411_/X sky130_fd_sc_hd__buf_1
XPHY_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14391_ _14382_/A _14390_/Y _20239_/Q _20031_/Q vssd1 vssd1 vccd1 vccd1 _14391_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18851__S _18908_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16130_ _16141_/A vssd1 vssd1 vccd1 vccd1 _16130_/X sky130_fd_sc_hd__buf_1
XFILLER_10_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13342_ _20524_/Q _13339_/X _13280_/X _13340_/X vssd1 vssd1 vccd1 vccd1 _20524_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_210_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10554_ _21324_/Q vssd1 vssd1 vccd1 vccd1 _10653_/A sky130_fd_sc_hd__inv_2
XFILLER_194_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17975__B _17978_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14165__A1 _20538_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15362__B1 _14258_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16061_ _19502_/Q _16056_/X _15776_/X _16057_/X vssd1 vssd1 vccd1 vccd1 _19502_/D
+ sky130_fd_sc_hd__a22o_1
X_13273_ _20559_/Q _13264_/X _13272_/X _13268_/X vssd1 vssd1 vccd1 vccd1 _20559_/D
+ sky130_fd_sc_hd__a22o_1
X_10485_ _21277_/Q vssd1 vssd1 vccd1 vccd1 _10754_/A sky130_fd_sc_hd__inv_2
XFILLER_154_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12224_ _20930_/Q _12222_/Y _20923_/Q _12223_/Y vssd1 vssd1 vccd1 vccd1 _12224_/X
+ sky130_fd_sc_hd__o22a_1
X_15012_ _15012_/A vssd1 vssd1 vccd1 vccd1 _15012_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19820_ _19820_/CLK _19820_/D vssd1 vssd1 vccd1 vccd1 _19820_/Q sky130_fd_sc_hd__dfxtp_1
X_12155_ _20971_/Q _12153_/Y _20977_/Q _12154_/Y vssd1 vssd1 vccd1 vccd1 _12155_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_2_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11106_ _11099_/B _11105_/Y _11100_/X _11101_/X _11054_/A vssd1 vssd1 vccd1 vccd1
+ _11107_/A sky130_fd_sc_hd__o32a_1
X_19751_ _19765_/CLK _19751_/D vssd1 vssd1 vccd1 vccd1 _19751_/Q sky130_fd_sc_hd__dfxtp_1
X_16963_ _19969_/Q _16963_/B vssd1 vssd1 vccd1 vccd1 _16979_/B sky130_fd_sc_hd__or2_1
X_12086_ _12081_/X _20374_/Q _12320_/A _20381_/Q _12085_/X vssd1 vssd1 vccd1 vccd1
+ _12087_/D sky130_fd_sc_hd__o221a_1
XANTENNA__18298__S _18886_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18702_ _17705_/Y _16599_/Y _20870_/Q vssd1 vssd1 vccd1 vccd1 _18702_/X sky130_fd_sc_hd__mux2_1
XFILLER_204_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11037_ _19966_/Q _19969_/Q _19973_/Q vssd1 vssd1 vccd1 vccd1 _11039_/C sky130_fd_sc_hd__or3_2
X_15914_ _19576_/Q _15911_/X _15879_/X _15912_/X vssd1 vssd1 vccd1 vccd1 _19576_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17406__A2 _17384_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19682_ _19813_/CLK _19682_/D vssd1 vssd1 vccd1 vccd1 _19682_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_237_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16894_ _16894_/A _16894_/B vssd1 vssd1 vccd1 vccd1 _16894_/Y sky130_fd_sc_hd__nor2_1
XFILLER_49_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18633_ _18632_/X _14595_/A _18748_/S vssd1 vssd1 vccd1 vccd1 _18633_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15845_ _19607_/Q _15841_/X _09838_/X _15842_/X vssd1 vssd1 vccd1 vccd1 _19607_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_225_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18564_ _18563_/X _16927_/A _18680_/S vssd1 vssd1 vccd1 vccd1 _18564_/X sky130_fd_sc_hd__mux2_2
XFILLER_52_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15776_ _16127_/A vssd1 vssd1 vccd1 vccd1 _15776_/X sky130_fd_sc_hd__buf_1
XFILLER_220_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12988_ _20697_/Q _12983_/X _12984_/X _12987_/X vssd1 vssd1 vccd1 vccd1 _20697_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_206_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17515_ _19594_/Q vssd1 vssd1 vccd1 vccd1 _17515_/Y sky130_fd_sc_hd__inv_2
X_14727_ _20145_/Q _14723_/X _13712_/X _14724_/X vssd1 vssd1 vccd1 vccd1 _20145_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_91_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18495_ _18494_/X _12297_/Y _18910_/S vssd1 vssd1 vccd1 vccd1 _18495_/X sky130_fd_sc_hd__mux2_1
X_11939_ _11944_/A _11944_/B vssd1 vssd1 vccd1 vccd1 _11940_/B sky130_fd_sc_hd__and2_1
XFILLER_221_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17231__A _17231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17446_ _17446_/A vssd1 vssd1 vccd1 vccd1 _17446_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_221_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14658_ _14655_/Y _19124_/S _14657_/X _14656_/A vssd1 vssd1 vccd1 vccd1 _14659_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_220_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13609_ _20395_/Q _13605_/X _13538_/X _13608_/X vssd1 vssd1 vccd1 vccd1 _20395_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_11_HCLK_A clkbuf_opt_2_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17377_ _21058_/Q vssd1 vssd1 vccd1 vccd1 _17377_/Y sky130_fd_sc_hd__inv_2
X_14589_ _14589_/A _14589_/B vssd1 vssd1 vccd1 vccd1 _14609_/A sky130_fd_sc_hd__or2_1
XANTENNA__18761__S _18930_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_74_HCLK_A clkbuf_4_13_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19116_ _19117_/S _11916_/Y _19116_/S vssd1 vssd1 vccd1 vccd1 _19116_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16328_ _16336_/A vssd1 vssd1 vccd1 vccd1 _16328_/X sky130_fd_sc_hd__buf_1
XFILLER_185_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15353__B1 _15352_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19047_ _16796_/X _20822_/Q _19058_/S vssd1 vssd1 vccd1 vccd1 _19929_/D sky130_fd_sc_hd__mux2_1
X_16259_ _19407_/Q _16255_/X _16125_/X _16256_/X vssd1 vssd1 vccd1 vccd1 _19407_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__20559__CLK _20592_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09684__A input64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19095__A1 _21083_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19190__S1 _20122_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19949_ _21374_/CLK _19949_/D repeater255/X vssd1 vssd1 vccd1 vccd1 _19949_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_96_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09702_ _11743_/A vssd1 vssd1 vccd1 vccd1 _09702_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_228_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09633_ input47/X vssd1 vssd1 vccd1 vccd1 _09633_/X sky130_fd_sc_hd__buf_4
XFILLER_56_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18936__S _18946_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20719__RESET_B repeater264/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_215_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18358__A0 _17281_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10102__C1 _10101_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20372__RESET_B repeater186/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17141__A _17141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20724_ _20724_/CLK _20724_/D repeater264/X vssd1 vssd1 vccd1 vccd1 _20724_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20655_ _20657_/CLK _20655_/D repeater197/X vssd1 vssd1 vccd1 vccd1 _20655_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12716__C _12716_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20586_ _20946_/CLK _20586_/D repeater258/X vssd1 vssd1 vccd1 vccd1 _20586_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_99_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15596__A _15603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15344__B1 _15343_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09594__A _20890_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10270_ _10270_/A _10402_/A vssd1 vssd1 vccd1 vccd1 _10271_/B sky130_fd_sc_hd__or2_2
X_21207_ _21207_/CLK _21207_/D repeater256/X vssd1 vssd1 vccd1 vccd1 _21207_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__19181__S1 _20124_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18833__A1 _11916_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21138_ _21147_/CLK _21138_/D repeater215/X vssd1 vssd1 vccd1 vccd1 _21138_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_94_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19007__S _19019_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21069_ _21087_/CLK _21069_/D repeater227/X vssd1 vssd1 vccd1 vccd1 _21069_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_58_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13960_ _13957_/Y _20304_/Q _20647_/Q _13971_/D _13959_/X vssd1 vssd1 vccd1 vccd1
+ _13961_/D sky130_fd_sc_hd__o221a_1
XFILLER_58_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18597__A0 _18848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12911_ _20730_/Q _12909_/X _12663_/X _12910_/X vssd1 vssd1 vccd1 vccd1 _20730_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_235_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13891_ _13891_/A _13891_/B vssd1 vssd1 vccd1 vccd1 _13983_/A sky130_fd_sc_hd__or2_2
XANTENNA__18846__S _18897_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15630_ _19707_/Q _15625_/X _15550_/X _15627_/X vssd1 vssd1 vccd1 vccd1 _19707_/D
+ sky130_fd_sc_hd__a22o_1
X_12842_ _12842_/A vssd1 vssd1 vccd1 vccd1 _12842_/X sky130_fd_sc_hd__buf_1
XFILLER_74_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19888__D _19888_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_131_HCLK clkbuf_4_4_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20951_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_55_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15561_ _15568_/A vssd1 vssd1 vccd1 vccd1 _15561_/X sky130_fd_sc_hd__buf_1
XPHY_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12773_ _20796_/Q _12771_/X _12673_/X _12772_/X vssd1 vssd1 vccd1 vccd1 _20796_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_203_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17300_ _21128_/Q vssd1 vssd1 vccd1 vccd1 _17300_/Y sky130_fd_sc_hd__inv_2
XPHY_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14512_ _14500_/A _14500_/B _14510_/Y _14469_/X vssd1 vssd1 vccd1 vccd1 _20215_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_9_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11724_ _21065_/Q _11720_/X _11571_/X _11721_/X vssd1 vssd1 vccd1 vccd1 _21065_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18280_ _19191_/X _21275_/Q _18281_/S vssd1 vssd1 vccd1 vccd1 _18280_/X sky130_fd_sc_hd__mux2_1
XPHY_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15492_ _15499_/A vssd1 vssd1 vccd1 vccd1 _15492_/X sky130_fd_sc_hd__buf_1
XPHY_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17231_ _17231_/A vssd1 vssd1 vccd1 vccd1 _17474_/A sky130_fd_sc_hd__buf_1
XPHY_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14443_ _21468_/Q vssd1 vssd1 vccd1 vccd1 _14443_/Y sky130_fd_sc_hd__inv_2
X_11655_ _17549_/A _11726_/B vssd1 vssd1 vccd1 vccd1 _11667_/B sky130_fd_sc_hd__or2_1
XANTENNA__18581__S _18748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10606_ _20757_/Q vssd1 vssd1 vccd1 vccd1 _10606_/Y sky130_fd_sc_hd__inv_2
XFILLER_156_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17162_ _17162_/A _17162_/B vssd1 vssd1 vccd1 vccd1 _17162_/X sky130_fd_sc_hd__or2_1
XPHY_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14374_ _14463_/D _14374_/B vssd1 vssd1 vccd1 vccd1 _14476_/A sky130_fd_sc_hd__or2_1
XPHY_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11586_ _11586_/A vssd1 vssd1 vccd1 vccd1 _11596_/B sky130_fd_sc_hd__inv_2
XPHY_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16113_ _20330_/Q vssd1 vssd1 vccd1 vccd1 _16113_/X sky130_fd_sc_hd__clkbuf_2
X_10537_ _21313_/Q vssd1 vssd1 vccd1 vccd1 _10540_/A sky130_fd_sc_hd__inv_2
X_13325_ _20531_/Q _13321_/X _13171_/X _13322_/X vssd1 vssd1 vccd1 vccd1 _20531_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_116_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17093_ _19494_/Q vssd1 vssd1 vccd1 vccd1 _17093_/Y sky130_fd_sc_hd__inv_2
XFILLER_171_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16044_ _19513_/Q _16042_/X _16009_/X _16043_/X vssd1 vssd1 vccd1 vccd1 _19513_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_6_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10468_ _21297_/Q vssd1 vssd1 vccd1 vccd1 _10773_/A sky130_fd_sc_hd__inv_2
X_13256_ _13254_/X _20564_/Q _13256_/S vssd1 vssd1 vccd1 vccd1 _20564_/D sky130_fd_sc_hd__mux2_1
X_12207_ _12060_/X _12087_/X _12145_/X _20982_/Q _12206_/X vssd1 vssd1 vccd1 vccd1
+ _20982_/D sky130_fd_sc_hd__a32o_1
XANTENNA__19172__S1 _20122_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13187_ _16525_/A _13184_/S _16525_/B _13186_/Y vssd1 vssd1 vccd1 vccd1 _20597_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_123_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10399_ _10399_/A vssd1 vssd1 vccd1 vccd1 _10399_/Y sky130_fd_sc_hd__inv_2
XFILLER_215_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12138_ _20959_/Q vssd1 vssd1 vccd1 vccd1 _12313_/B sky130_fd_sc_hd__inv_2
X_19803_ _19811_/CLK _19803_/D vssd1 vssd1 vccd1 vccd1 _19803_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_229_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13649__B1 _13511_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17995_ _18064_/A vssd1 vssd1 vccd1 vccd1 _17995_/X sky130_fd_sc_hd__buf_1
XFILLER_150_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12069_ _20963_/Q vssd1 vssd1 vccd1 vccd1 _12316_/A sky130_fd_sc_hd__inv_2
X_16946_ _19964_/Q _16937_/A _19965_/Q vssd1 vssd1 vccd1 vccd1 _16946_/X sky130_fd_sc_hd__o21a_1
XFILLER_84_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19734_ _21011_/CLK _19734_/D vssd1 vssd1 vccd1 vccd1 _19734_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__18588__A0 _17079_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20883__RESET_B repeater243/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19665_ _19765_/CLK _19665_/D vssd1 vssd1 vccd1 vccd1 _19665_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16877_ _16877_/A _16877_/B vssd1 vssd1 vccd1 vccd1 _16877_/Y sky130_fd_sc_hd__nor2_1
X_18616_ _18082_/Y _20767_/Q _18891_/S vssd1 vssd1 vccd1 vccd1 _18616_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15828_ _19615_/Q _15824_/X _09838_/X _15825_/X vssd1 vssd1 vccd1 vccd1 _19615_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_37_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10883__B1 _09666_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_231_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19596_ _19626_/CLK _19596_/D vssd1 vssd1 vccd1 vccd1 _19596_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_240_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18547_ _18848_/A0 _14148_/Y _18902_/S vssd1 vssd1 vccd1 vccd1 _18547_/X sky130_fd_sc_hd__mux2_1
X_15759_ _15768_/A vssd1 vssd1 vccd1 vccd1 _15770_/A sky130_fd_sc_hd__inv_2
X_18478_ _18848_/A0 _14122_/Y _18884_/S vssd1 vssd1 vccd1 vccd1 _18478_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17429_ _19449_/Q vssd1 vssd1 vccd1 vccd1 _17429_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17896__A _17896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_221_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10618__A _20763_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18491__S _18784_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20440_ _20937_/CLK _20440_/D repeater279/X vssd1 vssd1 vccd1 vccd1 _20440_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_193_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15326__B1 _13545_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20371_ _20422_/CLK _20371_/D repeater271/X vssd1 vssd1 vccd1 vccd1 _20371_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_146_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19068__A1 _21142_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_12_HCLK clkbuf_opt_2_HCLK/A vssd1 vssd1 vccd1 vccd1 _21011_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_161_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19163__S1 _20122_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18815__A1 _13928_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18579__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_217_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_154_HCLK clkbuf_opt_1_HCLK/A vssd1 vssd1 vccd1 vccd1 _19626_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_84_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18666__S _18666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11184__A _17290_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09616_ _20875_/Q _12716_/B _12716_/C vssd1 vssd1 vccd1 vccd1 _12898_/A sky130_fd_sc_hd__or3_4
XANTENNA__10874__B1 _09693_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19747__CLK _19765_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_243_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15014__C1 _14970_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20707_ _21357_/CLK _20707_/D repeater210/X vssd1 vssd1 vccd1 vccd1 _20707_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15565__B1 _15548_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11440_ _19871_/Q vssd1 vssd1 vccd1 vccd1 _11459_/A sky130_fd_sc_hd__inv_2
XFILLER_211_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20638_ _20657_/CLK _20638_/D repeater198/X vssd1 vssd1 vccd1 vccd1 _20638_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_138_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11371_ _11371_/A _11371_/B vssd1 vssd1 vccd1 vccd1 _16595_/B sky130_fd_sc_hd__nand2_1
XFILLER_50_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20569_ _20590_/CLK _20569_/D repeater260/X vssd1 vssd1 vccd1 vccd1 _20569_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_153_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13110_ _13110_/A _13261_/A vssd1 vssd1 vccd1 vccd1 _13138_/A sky130_fd_sc_hd__or2_2
XFILLER_50_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10322_ _10277_/A _20721_/Q _21350_/Q _10320_/Y _10321_/X vssd1 vssd1 vccd1 vccd1
+ _10323_/D sky130_fd_sc_hd__o221a_1
X_14090_ _14090_/A _14195_/A vssd1 vssd1 vccd1 vccd1 _14091_/B sky130_fd_sc_hd__or2_1
XFILLER_137_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13041_ _13041_/A vssd1 vssd1 vccd1 vccd1 _13041_/X sky130_fd_sc_hd__buf_1
XANTENNA__19154__S1 _21017_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10253_ _21350_/Q vssd1 vssd1 vccd1 vccd1 _10266_/A sky130_fd_sc_hd__inv_2
XFILLER_106_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12551__B1 _12550_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input46_A HWDATA[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10184_ _21397_/Q _10182_/Y _10183_/X _10159_/B vssd1 vssd1 vccd1 vccd1 _21397_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_182_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16800_ _19931_/Q vssd1 vssd1 vccd1 vccd1 _16800_/Y sky130_fd_sc_hd__inv_2
XFILLER_120_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17780_ _21063_/Q vssd1 vssd1 vccd1 vccd1 _17780_/Y sky130_fd_sc_hd__inv_2
X_14992_ _20091_/Q _14991_/Y _14870_/B _14978_/X vssd1 vssd1 vccd1 vccd1 _20091_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_247_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16731_ _20993_/Q _11999_/B _12000_/B vssd1 vssd1 vccd1 vccd1 _16731_/X sky130_fd_sc_hd__a21bo_1
X_13943_ _20637_/Q vssd1 vssd1 vccd1 vccd1 _13943_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20294__RESET_B repeater262/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18576__S _18904_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19450_ _21453_/CLK _19450_/D vssd1 vssd1 vccd1 vccd1 _19450_/Q sky130_fd_sc_hd__dfxtp_1
X_16662_ _19865_/Q _15299_/B _18962_/S vssd1 vssd1 vccd1 vccd1 _16662_/X sky130_fd_sc_hd__a21o_1
XANTENNA__20223__RESET_B repeater202/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13874_ _20301_/Q vssd1 vssd1 vccd1 vccd1 _13875_/A sky130_fd_sc_hd__inv_2
XFILLER_235_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18401_ _18400_/X _10267_/A _18841_/S vssd1 vssd1 vccd1 vccd1 _18401_/X sky130_fd_sc_hd__mux2_1
X_15613_ _15619_/A vssd1 vssd1 vccd1 vccd1 _15613_/X sky130_fd_sc_hd__buf_1
X_12825_ _20769_/Q _12821_/X _12651_/X _12824_/X vssd1 vssd1 vccd1 vccd1 _20769_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19381_ _19776_/CLK _19381_/D vssd1 vssd1 vccd1 vccd1 _19381_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16593_ _16616_/A _16593_/B vssd1 vssd1 vccd1 vccd1 _19117_/S sky130_fd_sc_hd__nor2_2
XFILLER_201_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_repeater185_A repeater186/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12918__A input52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18332_ _18848_/A0 _18043_/Y _18666_/S vssd1 vssd1 vccd1 vccd1 _18332_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15544_ _15657_/A vssd1 vssd1 vccd1 vccd1 _15544_/X sky130_fd_sc_hd__clkbuf_2
XPHY_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12756_ _12783_/A vssd1 vssd1 vccd1 vccd1 _12777_/A sky130_fd_sc_hd__buf_1
XPHY_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11707_ _21074_/Q _11704_/X _11568_/X _11705_/X vssd1 vssd1 vccd1 vccd1 _21074_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18263_ _18262_/X _13900_/Y _18903_/S vssd1 vssd1 vccd1 vccd1 _18263_/X sky130_fd_sc_hd__mux2_1
X_15475_ _15764_/A vssd1 vssd1 vccd1 vccd1 _15475_/X sky130_fd_sc_hd__buf_1
X_12687_ _12687_/A vssd1 vssd1 vccd1 vccd1 _12708_/A sky130_fd_sc_hd__buf_2
XPHY_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17214_ _18045_/A vssd1 vssd1 vccd1 vccd1 _17214_/X sky130_fd_sc_hd__buf_2
X_14426_ _14397_/Y _20210_/Q _14463_/C _21486_/Q _14425_/X vssd1 vssd1 vccd1 vccd1
+ _14434_/B sky130_fd_sc_hd__o221a_1
XFILLER_187_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11638_ _11638_/A _18983_/S vssd1 vssd1 vccd1 vccd1 _11641_/A sky130_fd_sc_hd__nand2_1
XFILLER_30_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18194_ _18193_/X _10277_/A _18886_/S vssd1 vssd1 vccd1 vccd1 _18194_/X sky130_fd_sc_hd__mux2_1
XPHY_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17145_ _21080_/Q vssd1 vssd1 vccd1 vccd1 _17145_/Y sky130_fd_sc_hd__inv_2
X_14357_ _20218_/Q vssd1 vssd1 vccd1 vccd1 _14503_/A sky130_fd_sc_hd__inv_2
XFILLER_156_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11569_ _21129_/Q _11562_/X _11568_/X _11566_/X vssd1 vssd1 vccd1 vccd1 _21129_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_6_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12790__B1 _09652_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13308_ _13322_/A vssd1 vssd1 vccd1 vccd1 _13308_/X sky130_fd_sc_hd__buf_1
XANTENNA__21011__RESET_B repeater235/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17076_ _21135_/Q _20892_/Q _17076_/C vssd1 vssd1 vccd1 vccd1 _17076_/X sky130_fd_sc_hd__and3_1
X_14288_ _14288_/A vssd1 vssd1 vccd1 vccd1 _14288_/X sky130_fd_sc_hd__buf_1
XFILLER_171_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19145__S1 _21017_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16027_ _19522_/Q _16021_/X _15766_/X _16023_/X vssd1 vssd1 vccd1 vccd1 _19522_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13239_ _13248_/A vssd1 vssd1 vccd1 vccd1 _13239_/X sky130_fd_sc_hd__buf_1
XFILLER_69_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17481__B1 _18779_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17978_ _17978_/A _17978_/B vssd1 vssd1 vccd1 vccd1 _17978_/Y sky130_fd_sc_hd__nor2_1
X_16929_ _19961_/Q vssd1 vssd1 vccd1 vccd1 _16931_/A sky130_fd_sc_hd__inv_2
XFILLER_66_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19717_ _20432_/CLK _19717_/D vssd1 vssd1 vccd1 vccd1 _19717_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12845__A1 _20755_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18486__S _18907_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17233__B1 _17230_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19648_ _19821_/CLK _19648_/D vssd1 vssd1 vccd1 vccd1 _19648_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_225_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19579_ _19626_/CLK _19579_/D vssd1 vssd1 vccd1 vccd1 _19579_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_240_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10084__B2 _10081_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15547__B1 _15544_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21472_ _21476_/CLK _21472_/D repeater204/X vssd1 vssd1 vccd1 vccd1 _21472_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__10067__B _10154_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20423_ _20951_/CLK _20423_/D repeater271/X vssd1 vssd1 vccd1 vccd1 _20423_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__13659__A _13679_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12781__B1 _09636_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20354_ _20972_/CLK _20354_/D repeater280/X vssd1 vssd1 vccd1 vccd1 _20354_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_134_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11179__A _16342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20285_ _20293_/CLK _20285_/D repeater262/X vssd1 vssd1 vccd1 vccd1 _20285_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_248_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20734__RESET_B repeater257/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18396__S _18896_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10940_ _21198_/Q vssd1 vssd1 vccd1 vccd1 _10940_/Y sky130_fd_sc_hd__inv_2
XFILLER_71_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15786__B1 _15785_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10871_ _10871_/A vssd1 vssd1 vccd1 vccd1 _10871_/X sky130_fd_sc_hd__buf_1
XFILLER_44_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12610_ input16/X _11793_/X _20866_/Q _11797_/X vssd1 vssd1 vccd1 vccd1 _20866_/D
+ sky130_fd_sc_hd__o22a_1
XPHY_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13590_ _20404_/Q _13588_/X _13506_/X _13589_/X vssd1 vssd1 vccd1 vccd1 _20404_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_243_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_58_HCLK clkbuf_4_14_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _21321_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_169_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12541_ _12527_/A _12525_/Y _19990_/Q _11307_/C _12520_/X vssd1 vssd1 vccd1 vccd1
+ _20901_/D sky130_fd_sc_hd__a32o_1
XFILLER_200_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_opt_2_HCLK_A clkbuf_opt_2_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19020__S _19026_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19988__RESET_B repeater218/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15260_ _20476_/Q vssd1 vssd1 vccd1 vccd1 _15260_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12472_ _12472_/A _12472_/B vssd1 vssd1 vccd1 vccd1 _12483_/A sky130_fd_sc_hd__or2_1
X_14211_ _14081_/A _14081_/B _14209_/Y _14207_/X vssd1 vssd1 vccd1 vccd1 _20271_/D
+ sky130_fd_sc_hd__a211oi_2
X_11423_ _11363_/B _11418_/X _11376_/C _11403_/A vssd1 vssd1 vccd1 vccd1 _21178_/D
+ sky130_fd_sc_hd__o22ai_1
XANTENNA__19917__RESET_B repeater220/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15191_ _15191_/A vssd1 vssd1 vccd1 vccd1 _15191_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11354_ _16595_/A _18968_/X vssd1 vssd1 vccd1 vccd1 _11409_/C sky130_fd_sc_hd__or2b_1
X_14142_ _20535_/Q vssd1 vssd1 vccd1 vccd1 _14142_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17983__B _18007_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10305_ _10288_/A _20732_/Q _21351_/Q _10304_/Y vssd1 vssd1 vccd1 vccd1 _10305_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_180_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19127__S1 _21017_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11285_ _20910_/Q vssd1 vssd1 vccd1 vccd1 _11313_/C sky130_fd_sc_hd__inv_2
X_18950_ _16660_/X _21086_/Q _18962_/S vssd1 vssd1 vccd1 vccd1 _18950_/X sky130_fd_sc_hd__mux2_1
X_14073_ _14073_/A _14225_/A vssd1 vssd1 vccd1 vccd1 _14074_/B sky130_fd_sc_hd__or2_2
XANTENNA__20899__SET_B repeater212/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10236_ _21367_/Q vssd1 vssd1 vccd1 vccd1 _10282_/A sky130_fd_sc_hd__inv_2
X_17901_ _17901_/A _17938_/B vssd1 vssd1 vccd1 vccd1 _17901_/Y sky130_fd_sc_hd__nor2_1
X_13024_ _20679_/Q _13019_/X _12855_/X _13021_/X vssd1 vssd1 vccd1 vccd1 _20679_/D
+ sky130_fd_sc_hd__a22o_1
X_18881_ _17187_/Y _10221_/B _18899_/S vssd1 vssd1 vccd1 vccd1 _18881_/X sky130_fd_sc_hd__mux2_1
X_17832_ _20406_/Q vssd1 vssd1 vccd1 vccd1 _17832_/Y sky130_fd_sc_hd__inv_2
XFILLER_239_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10167_ _21405_/Q _10164_/Y _10076_/C _10164_/A _10166_/X vssd1 vssd1 vccd1 vccd1
+ _21405_/D sky130_fd_sc_hd__o221a_1
XFILLER_120_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17763_ _19597_/Q vssd1 vssd1 vccd1 vccd1 _17763_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12827__A1 _20767_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14975_ _14989_/A vssd1 vssd1 vccd1 vccd1 _14975_/X sky130_fd_sc_hd__clkbuf_2
X_10098_ _10098_/A _10098_/B _10098_/C _10098_/D vssd1 vssd1 vccd1 vccd1 _10137_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_47_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16714_ _16718_/A _18936_/X vssd1 vssd1 vccd1 vccd1 _19900_/D sky130_fd_sc_hd__and2_1
X_19502_ _20326_/CLK _19502_/D vssd1 vssd1 vccd1 vccd1 _19502_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_212_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13926_ _20663_/Q _20320_/Q _20663_/Q _20320_/Q vssd1 vssd1 vccd1 vccd1 _13926_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_17694_ _19492_/Q vssd1 vssd1 vccd1 vccd1 _17694_/Y sky130_fd_sc_hd__inv_2
X_19433_ _21449_/CLK _19433_/D vssd1 vssd1 vccd1 vccd1 _19433_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_207_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16645_ _16663_/A vssd1 vssd1 vccd1 vccd1 _16652_/A sky130_fd_sc_hd__buf_1
XFILLER_74_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13857_ _13857_/A vssd1 vssd1 vccd1 vccd1 _13971_/C sky130_fd_sc_hd__buf_1
XANTENNA__12648__A _17083_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19364_ _21001_/CLK _19364_/D vssd1 vssd1 vccd1 vccd1 _19364_/Q sky130_fd_sc_hd__dfxtp_1
X_12808_ _20773_/Q _12803_/X _11743_/X _12804_/X vssd1 vssd1 vccd1 vccd1 _20773_/D
+ sky130_fd_sc_hd__a22o_1
X_16576_ _21095_/Q _16576_/B _19875_/Q _19841_/D vssd1 vssd1 vccd1 vccd1 _16576_/X
+ sky130_fd_sc_hd__or4_4
XFILLER_222_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13788_ _20193_/Q vssd1 vssd1 vccd1 vccd1 _14582_/A sky130_fd_sc_hd__inv_2
XFILLER_50_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18315_ _18030_/Y _20457_/Q _18906_/S vssd1 vssd1 vccd1 vccd1 _18315_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15527_ _19758_/Q _15516_/X _15526_/X _15519_/X vssd1 vssd1 vccd1 vccd1 _19758_/D
+ sky130_fd_sc_hd__a22o_1
X_19295_ _19813_/CLK _19295_/D vssd1 vssd1 vccd1 vccd1 _19295_/Q sky130_fd_sc_hd__dfxtp_1
X_12739_ _12746_/B vssd1 vssd1 vccd1 vccd1 _12739_/Y sky130_fd_sc_hd__inv_2
XFILLER_188_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09957__A _09957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18246_ _19146_/X _20164_/Q _18249_/S vssd1 vssd1 vccd1 vccd1 _18246_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13004__A1 _20690_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15458_ _19786_/Q _15449_/X _15421_/X _15452_/X vssd1 vssd1 vccd1 vccd1 _19786_/D
+ sky130_fd_sc_hd__a22o_1
X_14409_ _21465_/Q vssd1 vssd1 vccd1 vccd1 _14409_/Y sky130_fd_sc_hd__inv_2
XFILLER_163_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13479__A input50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18177_ _18176_/X _14439_/Y _18897_/S vssd1 vssd1 vccd1 vccd1 _18177_/X sky130_fd_sc_hd__mux2_1
X_15389_ _15389_/A vssd1 vssd1 vccd1 vccd1 _15389_/X sky130_fd_sc_hd__buf_1
XFILLER_117_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12763__B1 _12658_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17128_ _19454_/Q vssd1 vssd1 vccd1 vccd1 _17128_/Y sky130_fd_sc_hd__inv_2
XFILLER_116_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17059_ _17057_/Y _19847_/Q _11376_/D _17058_/X vssd1 vssd1 vccd1 vccd1 _19844_/D
+ sky130_fd_sc_hd__a31o_1
X_09950_ _09957_/A vssd1 vssd1 vccd1 vccd1 _09950_/X sky130_fd_sc_hd__buf_1
XFILLER_143_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_129_HCLK_A clkbuf_4_4_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09692__A _16338_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20070_ _20070_/CLK _20070_/D repeater276/X vssd1 vssd1 vccd1 vccd1 _20070_/Q sky130_fd_sc_hd__dfrtp_1
X_09881_ _09878_/A _09870_/X _09878_/Y vssd1 vssd1 vccd1 vccd1 _21439_/D sky130_fd_sc_hd__a21oi_1
XFILLER_106_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20145__RESET_B repeater250/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_239_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19105__S _19870_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20972_ _20972_/CLK _20972_/D repeater187/X vssd1 vssd1 vccd1 vccd1 _20972_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_122_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09695__B1 _09693_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18944__S _18946_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18182__A1 _21471_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21455_ _21457_/CLK _21455_/D repeater245/X vssd1 vssd1 vccd1 vccd1 _21455_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__15940__B1 _15893_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20406_ _20408_/CLK _20406_/D repeater184/X vssd1 vssd1 vccd1 vccd1 _20406_/Q sky130_fd_sc_hd__dfrtp_1
X_21386_ _21405_/CLK _21386_/D repeater252/X vssd1 vssd1 vccd1 vccd1 _21386_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__20915__RESET_B repeater218/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20337_ _20422_/CLK _20337_/D repeater271/X vssd1 vssd1 vccd1 vccd1 _20337_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11070_ _11063_/A _11067_/X _11063_/B _11067_/B vssd1 vssd1 vccd1 vccd1 _21238_/D
+ sky130_fd_sc_hd__o22ai_1
X_20268_ _20293_/CLK _20268_/D repeater263/X vssd1 vssd1 vccd1 vccd1 _20268_/Q sky130_fd_sc_hd__dfrtp_1
Xoutput79 _17235_/Y vssd1 vssd1 vccd1 vccd1 HRDATA[0] sky130_fd_sc_hd__clkbuf_2
X_10021_ _11621_/A _17031_/A vssd1 vssd1 vccd1 vccd1 _11614_/B sky130_fd_sc_hd__and2_1
XFILLER_49_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_248_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20199_ _20626_/CLK _20199_/D repeater193/X vssd1 vssd1 vccd1 vccd1 _20199_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_193_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_236_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19015__S _19019_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14760_ _14753_/A _14548_/X _14751_/A vssd1 vssd1 vccd1 vccd1 _14760_/X sky130_fd_sc_hd__o21a_1
XANTENNA__09686__B1 _09685_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11972_ _11972_/A vssd1 vssd1 vccd1 vccd1 _11972_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13711_ _20334_/Q _13706_/X _13710_/X _13708_/X vssd1 vssd1 vccd1 vccd1 _20334_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_244_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10923_ _21028_/Q vssd1 vssd1 vccd1 vccd1 _11805_/A sky130_fd_sc_hd__inv_2
X_14691_ _19286_/X _16490_/B _14688_/X _20167_/Q _14690_/X vssd1 vssd1 vccd1 vccd1
+ _20167_/D sky130_fd_sc_hd__a32o_1
XANTENNA__18854__S _18908_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16430_ _19319_/Q _16427_/X _15879_/A _16428_/X vssd1 vssd1 vccd1 vccd1 _19319_/D
+ sky130_fd_sc_hd__a22o_1
X_13642_ _20374_/Q _13639_/X _13432_/X _13640_/X vssd1 vssd1 vccd1 vccd1 _20374_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_232_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17978__B _17978_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10854_ _18278_/X _10853_/X _21272_/Q _10849_/X vssd1 vssd1 vccd1 vccd1 _21272_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_198_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16361_ _17072_/B _12006_/C _19889_/D _19357_/Q _16360_/X vssd1 vssd1 vccd1 vccd1
+ _19357_/D sky130_fd_sc_hd__a32o_1
XFILLER_188_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13573_ _13594_/A vssd1 vssd1 vccd1 vccd1 _13573_/X sky130_fd_sc_hd__buf_1
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10785_ _10785_/A vssd1 vssd1 vccd1 vccd1 _10830_/A sky130_fd_sc_hd__inv_2
X_18100_ _20428_/Q vssd1 vssd1 vccd1 vccd1 _18100_/Y sky130_fd_sc_hd__inv_2
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15312_ _15312_/A _17133_/B _17133_/A _15312_/D vssd1 vssd1 vccd1 vccd1 _15313_/S
+ sky130_fd_sc_hd__or4_4
X_12524_ _12527_/A vssd1 vssd1 vccd1 vccd1 _12524_/X sky130_fd_sc_hd__buf_1
XFILLER_169_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19080_ _16723_/X _20895_/Q _19908_/D vssd1 vssd1 vccd1 vccd1 _19080_/X sky130_fd_sc_hd__mux2_1
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16292_ _19392_/Q _16287_/X _16291_/X _16289_/X vssd1 vssd1 vccd1 vccd1 _19392_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18031_ _18031_/A _18032_/B vssd1 vssd1 vccd1 vccd1 _18031_/Y sky130_fd_sc_hd__nor2_1
XFILLER_200_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15243_ _20468_/Q vssd1 vssd1 vccd1 vccd1 _15243_/Y sky130_fd_sc_hd__inv_2
X_12455_ _12455_/A vssd1 vssd1 vccd1 vccd1 _12455_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15931__B1 _15793_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater148_A _18848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11406_ _21182_/Q _11401_/X _11409_/A _11404_/X vssd1 vssd1 vccd1 vccd1 _21182_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_138_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15174_ _20069_/Q _15173_/Y _15166_/X _15084_/B vssd1 vssd1 vccd1 vccd1 _20069_/D
+ sky130_fd_sc_hd__o211a_1
X_12386_ _12386_/A vssd1 vssd1 vccd1 vccd1 _12386_/Y sky130_fd_sc_hd__inv_2
X_14125_ _20560_/Q vssd1 vssd1 vccd1 vccd1 _14125_/Y sky130_fd_sc_hd__inv_2
X_11337_ _21180_/Q _11783_/D vssd1 vssd1 vccd1 vccd1 _11357_/D sky130_fd_sc_hd__or2_1
XFILLER_207_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19982_ _20075_/CLK _19982_/D repeater276/X vssd1 vssd1 vccd1 vccd1 _19982_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_140_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20592__CLK _20592_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18933_ _16719_/X _21143_/Q _18946_/S vssd1 vssd1 vccd1 vccd1 _18933_/X sky130_fd_sc_hd__mux2_1
X_14056_ _20272_/Q vssd1 vssd1 vccd1 vccd1 _14082_/A sky130_fd_sc_hd__inv_2
X_11268_ _11283_/C _11302_/A vssd1 vssd1 vccd1 vccd1 _12505_/A sky130_fd_sc_hd__or2_1
XFILLER_106_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13170__B1 _13169_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13007_ _13013_/A vssd1 vssd1 vccd1 vccd1 _13007_/X sky130_fd_sc_hd__buf_1
X_10219_ _21380_/Q _10223_/A _10216_/A _10140_/X vssd1 vssd1 vccd1 vccd1 _21380_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_228_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18864_ _18863_/X _14275_/Y _18929_/S vssd1 vssd1 vccd1 vccd1 _18864_/X sky130_fd_sc_hd__mux2_1
X_11199_ _11199_/A _12725_/B vssd1 vssd1 vccd1 vccd1 _17838_/A sky130_fd_sc_hd__or2_4
XFILLER_223_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17815_ _18085_/B vssd1 vssd1 vccd1 vccd1 _17944_/B sky130_fd_sc_hd__buf_2
XFILLER_39_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18795_ _18794_/X _19241_/X _18930_/S vssd1 vssd1 vccd1 vccd1 _18795_/X sky130_fd_sc_hd__mux2_2
XFILLER_67_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17746_ _19525_/Q vssd1 vssd1 vccd1 vccd1 _17746_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14958_ _14978_/A vssd1 vssd1 vccd1 vccd1 _14958_/X sky130_fd_sc_hd__buf_1
XFILLER_63_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19284__S0 _19285_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13909_ _20655_/Q _13971_/A _13908_/Y _20318_/Q vssd1 vssd1 vccd1 vccd1 _13909_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__21444__RESET_B repeater243/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17677_ _19724_/Q vssd1 vssd1 vccd1 vccd1 _17677_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14889_ _20591_/Q vssd1 vssd1 vccd1 vccd1 _14889_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18764__S _18928_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16628_ _16628_/A _17143_/A vssd1 vssd1 vccd1 vccd1 _19838_/D sky130_fd_sc_hd__nor2_2
X_19416_ _19784_/CLK _19416_/D vssd1 vssd1 vccd1 vccd1 _19416_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14422__B1 _21480_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16559_ _16689_/B _16535_/X _19994_/Q _16689_/B _16558_/X vssd1 vssd1 vccd1 vccd1
+ _19994_/D sky130_fd_sc_hd__a32o_1
X_19347_ _21453_/CLK _19347_/D vssd1 vssd1 vccd1 vccd1 _19347_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09687__A input63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19278_ _19549_/Q _19541_/Q _19533_/Q _19517_/Q _19280_/S0 _20122_/Q vssd1 vssd1
+ vccd1 vccd1 _19278_/X sky130_fd_sc_hd__mux4_2
X_18229_ _20853_/Q input2/X _18236_/S vssd1 vssd1 vccd1 vccd1 _18229_/X sky130_fd_sc_hd__mux2_1
XFILLER_164_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15201__B _15201_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11539__A1 _21136_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21240_ _21433_/CLK _21240_/D repeater236/X vssd1 vssd1 vccd1 vccd1 _21240_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_190_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20397__RESET_B repeater270/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21171_ _21182_/CLK _21171_/D repeater216/X vssd1 vssd1 vccd1 vccd1 _21171_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_132_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12841__A _12841_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16313__A _16319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20326__RESET_B repeater250/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20122_ _21273_/CLK _20122_/D repeater247/X vssd1 vssd1 vccd1 vccd1 _20122_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_104_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09933_ _14304_/A vssd1 vssd1 vccd1 vccd1 _11654_/A sky130_fd_sc_hd__buf_1
XFILLER_120_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18939__S _18946_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13161__B1 _12954_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20053_ _20066_/CLK _20053_/D repeater281/X vssd1 vssd1 vccd1 vccd1 _20053_/Q sky130_fd_sc_hd__dfrtp_1
X_09864_ _09864_/A _15314_/A vssd1 vssd1 vccd1 vccd1 _09864_/X sky130_fd_sc_hd__or2_1
XFILLER_133_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09795_ _09795_/A vssd1 vssd1 vccd1 vccd1 _09795_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater151 _18902_/S vssd1 vssd1 vccd1 vccd1 _18884_/S sky130_fd_sc_hd__clkbuf_16
Xrepeater162 _18880_/S vssd1 vssd1 vccd1 vccd1 _18617_/S sky130_fd_sc_hd__buf_8
XFILLER_73_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater173 _18879_/S vssd1 vssd1 vccd1 vccd1 _18775_/S sky130_fd_sc_hd__buf_6
XPHY_4305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19275__S0 _19275_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater184 repeater185/X vssd1 vssd1 vccd1 vccd1 repeater184/X sky130_fd_sc_hd__buf_6
Xrepeater195 repeater196/X vssd1 vssd1 vccd1 vccd1 repeater195/X sky130_fd_sc_hd__buf_6
XFILLER_66_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20955_ _20981_/CLK _20955_/D repeater187/X vssd1 vssd1 vccd1 vccd1 _20955_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__18674__S _18928_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21114__RESET_B repeater233/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_242_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_214_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20886_ _21444_/CLK _20886_/D repeater246/X vssd1 vssd1 vccd1 vccd1 _20886_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11227__B1 _10894_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18155__A1 _10588_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10570_ _21335_/Q vssd1 vssd1 vccd1 vccd1 _10664_/A sky130_fd_sc_hd__inv_2
XFILLER_21_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12240_ _20926_/Q vssd1 vssd1 vccd1 vccd1 _12474_/A sky130_fd_sc_hd__inv_2
XFILLER_107_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21438_ _21438_/CLK _21438_/D repeater239/X vssd1 vssd1 vccd1 vccd1 _21438_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_182_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12171_ _20980_/Q _12168_/Y _20961_/Q _12169_/Y _12170_/X vssd1 vssd1 vccd1 vccd1
+ _12175_/C sky130_fd_sc_hd__a221o_1
X_21369_ _21374_/CLK _21369_/D repeater254/X vssd1 vssd1 vccd1 vccd1 _21369_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__20067__RESET_B repeater276/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10753__A2 _10752_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11122_ _09744_/X _11066_/B _11050_/A _11113_/X vssd1 vssd1 vccd1 vccd1 _21224_/D
+ sky130_fd_sc_hd__o22a_1
XANTENNA_clkbuf_leaf_112_HCLK_A clkbuf_opt_3_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18849__S _18849_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11053_ _11053_/A _11108_/A vssd1 vssd1 vccd1 vccd1 _11104_/A sky130_fd_sc_hd__or2_1
X_15930_ _19568_/Q _15927_/X _15791_/X _15928_/X vssd1 vssd1 vccd1 vccd1 _19568_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_49_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10004_ _09999_/X _10000_/X _09999_/X _10000_/X vssd1 vssd1 vccd1 vccd1 _10005_/A
+ sky130_fd_sc_hd__o2bb2a_1
X_15861_ _19598_/Q _15856_/X _15795_/X _15857_/X vssd1 vssd1 vccd1 vccd1 _19598_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_190_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17600_ _19715_/Q vssd1 vssd1 vccd1 vccd1 _17600_/Y sky130_fd_sc_hd__inv_2
XFILLER_218_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14812_ _14800_/A _14807_/X _14800_/A _14807_/X vssd1 vssd1 vccd1 vccd1 _20117_/D
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_190_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18580_ _18579_/X _14435_/Y _18669_/S vssd1 vssd1 vccd1 vccd1 _18580_/X sky130_fd_sc_hd__mux2_1
XANTENNA__19266__S0 _21005_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15792_ _19632_/Q _15787_/X _15791_/X _15789_/X vssd1 vssd1 vccd1 vccd1 _19632_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_92_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17531_ _20143_/Q vssd1 vssd1 vccd1 vccd1 _17531_/Y sky130_fd_sc_hd__inv_2
X_14743_ _15816_/A _14536_/X _14541_/Y _19122_/X _14742_/X vssd1 vssd1 vccd1 vccd1
+ _20137_/D sky130_fd_sc_hd__a41o_1
X_11955_ _11955_/A _11955_/B vssd1 vssd1 vccd1 vccd1 _21005_/D sky130_fd_sc_hd__nor2_1
XANTENNA__18394__A1 _13919_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18584__S _18841_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17462_ _20896_/Q vssd1 vssd1 vccd1 vccd1 _17462_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10906_ _17019_/A vssd1 vssd1 vccd1 vccd1 _17026_/B sky130_fd_sc_hd__buf_1
XFILLER_178_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14674_ _14674_/A vssd1 vssd1 vccd1 vccd1 _14674_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_60_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11886_ _11886_/A vssd1 vssd1 vccd1 vccd1 _11886_/Y sky130_fd_sc_hd__inv_2
XFILLER_220_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16413_ _16413_/A vssd1 vssd1 vccd1 vccd1 _16413_/X sky130_fd_sc_hd__buf_1
X_19201_ _19197_/X _19198_/X _19199_/X _19200_/X _20132_/Q _20133_/Q vssd1 vssd1 vccd1
+ vccd1 _19201_/X sky130_fd_sc_hd__mux4_2
X_13625_ _13625_/A vssd1 vssd1 vccd1 vccd1 _13625_/X sky130_fd_sc_hd__buf_1
XANTENNA__11218__B1 _09666_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17393_ _16690_/Y _17286_/X _17385_/Y _17147_/X _17392_/X vssd1 vssd1 vccd1 vccd1
+ _17393_/X sky130_fd_sc_hd__o221a_2
X_10837_ _21280_/Q _10836_/Y _10830_/X _10758_/B vssd1 vssd1 vccd1 vccd1 _21280_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA_repeater265_A repeater267/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19132_ _19679_/Q _19807_/Q _19799_/Q _19791_/Q _19285_/S0 _21017_/Q vssd1 vssd1
+ vccd1 vccd1 _19132_/X sky130_fd_sc_hd__mux4_2
XFILLER_186_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16344_ _16344_/A _16344_/B _16344_/C vssd1 vssd1 vccd1 vccd1 _16352_/A sky130_fd_sc_hd__or3_4
X_13556_ _20422_/Q _13549_/X _13555_/X _13551_/X vssd1 vssd1 vccd1 vccd1 _20422_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_13_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10768_ _10768_/A _10815_/A vssd1 vssd1 vccd1 vccd1 _10769_/B sky130_fd_sc_hd__or2_2
XANTENNA__20837__RESET_B repeater257/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12507_ _12507_/A _16569_/A _16689_/C _12506_/X vssd1 vssd1 vccd1 vccd1 _12507_/X
+ sky130_fd_sc_hd__or4b_4
X_19063_ _21188_/Q _21130_/Q _19910_/Q vssd1 vssd1 vccd1 vccd1 _19063_/X sky130_fd_sc_hd__mux2_1
X_16275_ _16344_/A _16344_/B _16465_/C vssd1 vssd1 vccd1 vccd1 _16287_/A sky130_fd_sc_hd__or3_4
X_13487_ input46/X vssd1 vssd1 vccd1 vccd1 _13487_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_139_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10699_ _10651_/A _10651_/B _10697_/Y _10729_/C vssd1 vssd1 vccd1 vccd1 _21322_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_9_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12718__A0 _11179_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18014_ _18014_/A _18014_/B _18014_/C _18014_/D vssd1 vssd1 vccd1 vccd1 _18014_/X
+ sky130_fd_sc_hd__or4_4
X_15226_ _20475_/Q vssd1 vssd1 vccd1 vccd1 _15226_/Y sky130_fd_sc_hd__inv_2
XFILLER_172_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12438_ _12462_/A vssd1 vssd1 vccd1 vccd1 _12438_/X sky130_fd_sc_hd__buf_1
XFILLER_161_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17657__B1 _18710_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15157_ _15157_/A _15157_/B _15157_/C _15157_/D vssd1 vssd1 vccd1 vccd1 _15157_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_126_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12369_ _12369_/A vssd1 vssd1 vccd1 vccd1 _12369_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14108_ _20553_/Q vssd1 vssd1 vccd1 vccd1 _14108_/Y sky130_fd_sc_hd__inv_2
X_19965_ _20413_/CLK _19965_/D repeater184/X vssd1 vssd1 vccd1 vccd1 _19965_/Q sky130_fd_sc_hd__dfrtp_1
X_15088_ _15088_/A _15088_/B vssd1 vssd1 vccd1 vccd1 _15089_/A sky130_fd_sc_hd__or2_1
XFILLER_102_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18759__S _18928_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13143__B1 _13140_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14039_ _20289_/Q vssd1 vssd1 vccd1 vccd1 _14099_/A sky130_fd_sc_hd__inv_2
X_18916_ _18915_/X _21430_/Q _18920_/S vssd1 vssd1 vccd1 vccd1 _18916_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19896_ _21191_/CLK _19896_/D repeater222/X vssd1 vssd1 vccd1 vccd1 _19896_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_68_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18847_ _18846_/X _14567_/A _18898_/S vssd1 vssd1 vccd1 vccd1 _18847_/X sky130_fd_sc_hd__mux2_2
XANTENNA_clkbuf_leaf_34_HCLK_A clkbuf_opt_4_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_97_HCLK_A clkbuf_4_13_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_243_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19257__S0 _20130_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18778_ _18777_/X _14438_/Y _18897_/S vssd1 vssd1 vccd1 vccd1 _18778_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17729_ _18702_/X _17472_/X _18701_/X _17474_/X vssd1 vssd1 vccd1 vccd1 _17729_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__18494__S _18787_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20740_ _21306_/CLK _20740_/D repeater207/X vssd1 vssd1 vccd1 vccd1 _20740_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__16396__B1 _16235_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11209__B1 _09641_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20671_ _21294_/CLK _20671_/D repeater211/X vssd1 vssd1 vccd1 vccd1 _20671_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12836__A _12842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12709__B1 _11736_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13382__B1 _13173_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21223_ _21223_/CLK _21223_/D repeater241/X vssd1 vssd1 vccd1 vccd1 _21223_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__13667__A _13679_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21154_ _21429_/CLK _21154_/D repeater229/X vssd1 vssd1 vccd1 vccd1 _21154_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__13386__B _17174_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18669__S _18669_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13134__B1 _12925_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20105_ _20107_/CLK _20105_/D repeater259/X vssd1 vssd1 vccd1 vccd1 _20105_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_160_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09916_ _09916_/A _09916_/B _20013_/D _09915_/X vssd1 vssd1 vccd1 vccd1 _11584_/B
+ sky130_fd_sc_hd__or4b_4
X_21085_ _21087_/CLK _21085_/D repeater227/X vssd1 vssd1 vccd1 vccd1 _21085_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_247_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20036_ _21184_/CLK _20036_/D repeater220/X vssd1 vssd1 vccd1 vccd1 _20036_/Q sky130_fd_sc_hd__dfrtp_1
X_09847_ _09847_/A _09871_/A vssd1 vssd1 vccd1 vccd1 _10843_/C sky130_fd_sc_hd__or2_1
XFILLER_112_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21366__RESET_B repeater254/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09778_ _21461_/Q _21460_/Q _16617_/A vssd1 vssd1 vccd1 vccd1 _09778_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__19248__S0 _20130_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_233_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_233_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ _21058_/Q _11735_/X _11739_/X _11737_/X vssd1 vssd1 vccd1 vccd1 _21058_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_15_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20938_ _20950_/CLK _20938_/D repeater278/X vssd1 vssd1 vccd1 vccd1 _20938_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_202_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11671_ _16654_/A _11657_/A _11670_/Y _11516_/Y _11676_/S vssd1 vssd1 vccd1 vccd1
+ _11672_/A sky130_fd_sc_hd__o32a_1
XPHY_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20869_ _21431_/CLK _20869_/D repeater237/X vssd1 vssd1 vccd1 vccd1 _20869_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13410_ _13410_/A vssd1 vssd1 vccd1 vccd1 _13410_/X sky130_fd_sc_hd__buf_1
XPHY_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10622_ _10608_/X _10622_/B _10622_/C _10622_/D vssd1 vssd1 vccd1 vccd1 _10639_/C
+ sky130_fd_sc_hd__and4b_1
X_14390_ _20031_/Q vssd1 vssd1 vccd1 vccd1 _14390_/Y sky130_fd_sc_hd__inv_2
XPHY_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13341_ _20525_/Q _13339_/X _13277_/X _13340_/X vssd1 vssd1 vccd1 vccd1 _20525_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17887__B1 _18489_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10553_ _21325_/Q vssd1 vssd1 vccd1 vccd1 _10654_/A sky130_fd_sc_hd__inv_2
X_16060_ _19503_/Q _16056_/X _15774_/X _16057_/X vssd1 vssd1 vccd1 vccd1 _19503_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_input76_A scl_i_S5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13272_ input59/X vssd1 vssd1 vccd1 vccd1 _13272_/X sky130_fd_sc_hd__clkbuf_2
X_10484_ _20692_/Q vssd1 vssd1 vccd1 vccd1 _10484_/Y sky130_fd_sc_hd__inv_2
XFILLER_154_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15011_ _15004_/A _15004_/B _15009_/Y _14970_/X vssd1 vssd1 vccd1 vccd1 _20084_/D
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__13373__B1 _13240_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12223_ _20503_/Q vssd1 vssd1 vccd1 vccd1 _12223_/Y sky130_fd_sc_hd__inv_2
XFILLER_136_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15114__A1 _20451_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12154_ _20359_/Q vssd1 vssd1 vccd1 vccd1 _12154_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18579__S _18896_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13125__B1 _13003_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11105_ _21229_/Q _11105_/B vssd1 vssd1 vccd1 vccd1 _11105_/Y sky130_fd_sc_hd__nor2_1
XFILLER_2_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19750_ _21009_/CLK _19750_/D vssd1 vssd1 vccd1 vccd1 _19750_/Q sky130_fd_sc_hd__dfxtp_1
X_16962_ _19969_/Q vssd1 vssd1 vccd1 vccd1 _16966_/A sky130_fd_sc_hd__inv_2
X_12085_ _20960_/Q _12083_/Y _20954_/Q _17539_/A vssd1 vssd1 vccd1 vccd1 _12085_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_150_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18701_ _17706_/Y _16598_/Y _20870_/Q vssd1 vssd1 vccd1 vccd1 _18701_/X sky130_fd_sc_hd__mux2_1
X_15913_ _19577_/Q _15911_/X _15876_/X _15912_/X vssd1 vssd1 vccd1 vccd1 _19577_/D
+ sky130_fd_sc_hd__a22o_1
X_11036_ _19965_/Q _19964_/Q _16937_/A vssd1 vssd1 vccd1 vccd1 _16949_/B sky130_fd_sc_hd__or3_4
XFILLER_110_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16893_ _19952_/Q _16892_/A _16891_/Y _16892_/Y vssd1 vssd1 vccd1 vccd1 _16894_/B
+ sky130_fd_sc_hd__o22a_1
X_19681_ _19820_/CLK _19681_/D vssd1 vssd1 vccd1 vccd1 _19681_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_237_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18632_ _18631_/X _14390_/Y _18669_/S vssd1 vssd1 vccd1 vccd1 _18632_/X sky130_fd_sc_hd__mux2_1
X_15844_ _19608_/Q _15841_/X _09835_/X _15842_/X vssd1 vssd1 vccd1 vccd1 _19608_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_225_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19239__S0 _20130_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21036__RESET_B repeater242/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18563_ _17281_/X _17851_/Y _18835_/S vssd1 vssd1 vccd1 vccd1 _18563_/X sky130_fd_sc_hd__mux2_1
X_15775_ _19639_/Q _15768_/X _15774_/X _15770_/X vssd1 vssd1 vccd1 vccd1 _19639_/D
+ sky130_fd_sc_hd__a22o_1
X_12987_ _13013_/A vssd1 vssd1 vccd1 vccd1 _12987_/X sky130_fd_sc_hd__buf_1
XANTENNA__18367__A1 _20758_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17514_ _19610_/Q vssd1 vssd1 vccd1 vccd1 _17514_/Y sky130_fd_sc_hd__inv_2
X_14726_ _20146_/Q _14723_/X _13710_/X _14724_/X vssd1 vssd1 vccd1 vccd1 _20146_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_206_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18494_ _18493_/X _12164_/Y _18787_/S vssd1 vssd1 vccd1 vccd1 _18494_/X sky130_fd_sc_hd__mux2_2
X_11938_ _11936_/Y _19116_/S _11940_/A _11165_/X vssd1 vssd1 vccd1 vccd1 _11944_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_32_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_221_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17445_ _19336_/Q vssd1 vssd1 vccd1 vccd1 _17446_/A sky130_fd_sc_hd__inv_2
X_14657_ _20173_/Q vssd1 vssd1 vccd1 vccd1 _14657_/X sky130_fd_sc_hd__buf_1
XANTENNA__12656__A input61/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11869_ _21025_/Q _10934_/X _21026_/Q _11868_/X vssd1 vssd1 vccd1 vccd1 _11869_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_221_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11560__A _13163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12939__B1 _12853_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13608_ _13626_/A vssd1 vssd1 vccd1 vccd1 _13608_/X sky130_fd_sc_hd__buf_1
X_17376_ _17376_/A vssd1 vssd1 vccd1 vccd1 _17376_/X sky130_fd_sc_hd__buf_1
X_14588_ _14588_/A _14613_/A vssd1 vssd1 vccd1 vccd1 _14589_/B sky130_fd_sc_hd__or2_2
XANTENNA__20671__RESET_B repeater211/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16327_ _16334_/A vssd1 vssd1 vccd1 vccd1 _16336_/A sky130_fd_sc_hd__inv_2
X_19115_ _16594_/Y _11986_/Y _19115_/S vssd1 vssd1 vccd1 vccd1 _19115_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13539_ _13572_/A vssd1 vssd1 vccd1 vccd1 _13574_/A sky130_fd_sc_hd__inv_2
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19046_ _16799_/Y _20823_/Q _19046_/S vssd1 vssd1 vccd1 vccd1 _19930_/D sky130_fd_sc_hd__mux2_1
X_16258_ _19408_/Q _16255_/X _16123_/X _16256_/X vssd1 vssd1 vccd1 vccd1 _19408_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_173_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15209_ _20049_/Q _15208_/Y _15065_/B _15177_/X vssd1 vssd1 vccd1 vccd1 _20049_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12167__B2 _20347_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13487__A input46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13364__B1 _13148_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16189_ _19441_/Q _16187_/X _16142_/X _16188_/X vssd1 vssd1 vccd1 vccd1 _19441_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_142_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18489__S _18907_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13116__B1 _12984_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19948_ _20841_/CLK _19948_/D repeater256/X vssd1 vssd1 vccd1 vccd1 _19948_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_229_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09701_ _15354_/A vssd1 vssd1 vccd1 vccd1 _11743_/A sky130_fd_sc_hd__buf_1
X_19879_ _21193_/CLK _19879_/D repeater224/X vssd1 vssd1 vccd1 vccd1 _19879_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_56_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09632_ _09657_/A vssd1 vssd1 vccd1 vccd1 _09632_/X sky130_fd_sc_hd__buf_1
XFILLER_55_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17802__B1 _18392_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_215_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20723_ _21366_/CLK _20723_/D repeater264/X vssd1 vssd1 vccd1 vccd1 _20723_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_23_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18952__S _18962_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17318__C1 _17317_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20654_ _20657_/CLK _20654_/D repeater197/X vssd1 vssd1 vccd1 vccd1 _20654_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_23_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_91_HCLK clkbuf_4_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _21366_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_183_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20585_ _20946_/CLK _20585_/D repeater258/X vssd1 vssd1 vccd1 vccd1 _20585_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_139_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18530__A1 _20790_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21206_ _21401_/CLK _21206_/D repeater256/X vssd1 vssd1 vccd1 vccd1 _21206_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__18399__S _18884_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21137_ _21147_/CLK _21137_/D repeater215/X vssd1 vssd1 vccd1 vccd1 _21137_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_78_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21068_ _21087_/CLK _21068_/D repeater228/X vssd1 vssd1 vccd1 vccd1 _21068_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_48_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20019_ _21417_/CLK _20019_/D repeater230/X vssd1 vssd1 vccd1 vccd1 _20019_/Q sky130_fd_sc_hd__dfrtp_1
X_12910_ _12926_/A vssd1 vssd1 vccd1 vccd1 _12910_/X sky130_fd_sc_hd__buf_1
XFILLER_207_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__21009__CLK _21009_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13890_ _13974_/C _13986_/A vssd1 vssd1 vccd1 vccd1 _13891_/B sky130_fd_sc_hd__or2_2
XFILLER_235_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12841_ _12841_/A vssd1 vssd1 vccd1 vccd1 _12841_/X sky130_fd_sc_hd__buf_1
XANTENNA_clkbuf_leaf_80_HCLK_A clkbuf_opt_7_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19023__S _19026_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15560_ _15673_/A _15778_/B _15708_/C vssd1 vssd1 vccd1 vccd1 _15568_/A sky130_fd_sc_hd__or3_4
XPHY_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12772_ _12778_/A vssd1 vssd1 vccd1 vccd1 _12772_/X sky130_fd_sc_hd__buf_1
XPHY_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14511_ _20216_/Q _14510_/Y _14502_/B _14453_/X vssd1 vssd1 vccd1 vccd1 _20216_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ _21066_/Q _11720_/X _11568_/X _11721_/X vssd1 vssd1 vccd1 vccd1 _21066_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_202_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15491_ _16325_/A _15624_/B _16229_/C vssd1 vssd1 vccd1 vccd1 _15499_/A sky130_fd_sc_hd__or3_4
XFILLER_9_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18862__S _18927_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20429__RESET_B repeater190/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17230_ _18916_/X vssd1 vssd1 vccd1 vccd1 _17230_/Y sky130_fd_sc_hd__inv_2
X_14442_ _20029_/Q vssd1 vssd1 vccd1 vccd1 _14442_/Y sky130_fd_sc_hd__inv_2
XPHY_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11654_ _11654_/A _17157_/D vssd1 vssd1 vccd1 vccd1 _11726_/B sky130_fd_sc_hd__or2_2
XANTENNA__16780__B1 _16779_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10605_ _10605_/A _10605_/B _10605_/C _10605_/D vssd1 vssd1 vccd1 vccd1 _10639_/B
+ sky130_fd_sc_hd__and4_1
X_17161_ _21127_/Q vssd1 vssd1 vccd1 vccd1 _17161_/Y sky130_fd_sc_hd__inv_2
XPHY_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14373_ _14460_/A _14480_/A vssd1 vssd1 vccd1 vccd1 _14374_/B sky130_fd_sc_hd__or2_2
XFILLER_155_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11585_ _11590_/B _11591_/A vssd1 vssd1 vccd1 vccd1 _11586_/A sky130_fd_sc_hd__or2b_1
XFILLER_167_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16112_ _19477_/Q _16108_/X _16109_/X _16111_/X vssd1 vssd1 vccd1 vccd1 _19477_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09785__A _14309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13324_ _20532_/Q _13321_/X _13169_/X _13322_/X vssd1 vssd1 vccd1 vccd1 _20532_/D
+ sky130_fd_sc_hd__a22o_1
X_10536_ _21314_/Q vssd1 vssd1 vccd1 vccd1 _10702_/A sky130_fd_sc_hd__inv_2
X_17092_ _21242_/Q _20810_/Q vssd1 vssd1 vccd1 vccd1 _17092_/X sky130_fd_sc_hd__and2_4
XFILLER_171_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16043_ _16043_/A vssd1 vssd1 vccd1 vccd1 _16043_/X sky130_fd_sc_hd__buf_1
X_13255_ _17178_/A _13259_/B vssd1 vssd1 vccd1 vccd1 _13256_/S sky130_fd_sc_hd__or2_1
X_10467_ _21287_/Q vssd1 vssd1 vccd1 vccd1 _10763_/A sky130_fd_sc_hd__inv_2
XFILLER_182_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18285__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12206_ _12373_/A vssd1 vssd1 vccd1 vccd1 _12206_/X sky130_fd_sc_hd__buf_1
XANTENNA__21288__RESET_B repeater207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13186_ _12968_/A _13185_/X _13184_/S vssd1 vssd1 vccd1 vccd1 _13186_/Y sky130_fd_sc_hd__a21oi_1
X_10398_ _10273_/A _10273_/B _10394_/Y _10397_/X vssd1 vssd1 vccd1 vccd1 _21358_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_123_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19802_ _19811_/CLK _19802_/D vssd1 vssd1 vccd1 vccd1 _19802_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_215_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12137_ _20366_/Q vssd1 vssd1 vccd1 vccd1 _12137_/Y sky130_fd_sc_hd__inv_2
XFILLER_111_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17994_ _18344_/X _17926_/X _18216_/X _17927_/X _17993_/X vssd1 vssd1 vccd1 vccd1
+ _17999_/B sky130_fd_sc_hd__o221a_2
X_19733_ _19777_/CLK _19733_/D vssd1 vssd1 vccd1 vccd1 _19733_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12068_ _20979_/Q vssd1 vssd1 vccd1 vccd1 _12332_/A sky130_fd_sc_hd__inv_2
X_16945_ _16949_/B vssd1 vssd1 vccd1 vccd1 _16951_/B sky130_fd_sc_hd__inv_2
XFILLER_237_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11019_ _17027_/A _20005_/Q vssd1 vssd1 vccd1 vccd1 _18992_/S sky130_fd_sc_hd__or2_4
XFILLER_237_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19664_ _19811_/CLK _19664_/D vssd1 vssd1 vccd1 vccd1 _19664_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16876_ _19948_/Q _16872_/A _16875_/Y _16872_/Y vssd1 vssd1 vccd1 vccd1 _16877_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_231_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18615_ _17830_/X _09747_/Y _18928_/S vssd1 vssd1 vccd1 vccd1 _18615_/X sky130_fd_sc_hd__mux2_1
X_15827_ _19616_/Q _15824_/X _09835_/X _15825_/X vssd1 vssd1 vccd1 vccd1 _19616_/D
+ sky130_fd_sc_hd__a22o_1
X_19595_ _19626_/CLK _19595_/D vssd1 vssd1 vccd1 vccd1 _19595_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18546_ _18545_/X _10763_/A _18617_/S vssd1 vssd1 vccd1 vccd1 _18546_/X sky130_fd_sc_hd__mux2_1
X_15758_ _15758_/A vssd1 vssd1 vccd1 vccd1 _15758_/X sky130_fd_sc_hd__buf_1
XFILLER_240_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20852__RESET_B repeater243/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14709_ _20157_/Q _14704_/X _12855_/A _14706_/X vssd1 vssd1 vccd1 vccd1 _20157_/D
+ sky130_fd_sc_hd__a22o_1
X_15689_ _15696_/A vssd1 vssd1 vccd1 vccd1 _15698_/A sky130_fd_sc_hd__inv_2
XFILLER_100_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18477_ _18476_/X _14084_/A _18904_/S vssd1 vssd1 vccd1 vccd1 _18477_/X sky130_fd_sc_hd__mux2_1
XANTENNA__18772__S _18879_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_221_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17428_ _19481_/Q vssd1 vssd1 vccd1 vccd1 _17428_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17896__B _17898_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13585__B1 _13584_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19699__CLK _21009_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17359_ _19432_/Q vssd1 vssd1 vccd1 vccd1 _17359_/Y sky130_fd_sc_hd__inv_2
X_20370_ _20957_/CLK _20370_/D repeater187/X vssd1 vssd1 vccd1 vccd1 _20370_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_118_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15326__A1 _20030_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13337__B1 _13272_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19029_ _16874_/X _20840_/Q _19046_/S vssd1 vssd1 vccd1 vccd1 _19947_/D sky130_fd_sc_hd__mux2_1
XFILLER_133_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09615_ _20880_/Q _20879_/Q _09615_/C _09615_/D vssd1 vssd1 vccd1 vccd1 _12716_/C
+ sky130_fd_sc_hd__or4_4
XFILLER_28_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13680__A _13680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20593__RESET_B repeater259/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_221_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18200__A0 _17281_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18682__S _18880_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20706_ _21349_/CLK _20706_/D repeater210/X vssd1 vssd1 vccd1 vccd1 _20706_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__21451__CLK _21452_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13576__B1 _13418_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20637_ _21486_/CLK _20637_/D repeater198/X vssd1 vssd1 vccd1 vccd1 _20637_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__18503__A1 _10609_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11370_ _11387_/B _11379_/B _11387_/A vssd1 vssd1 vccd1 vccd1 _11371_/B sky130_fd_sc_hd__or3b_4
XFILLER_153_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20568_ _20590_/CLK _20568_/D repeater260/X vssd1 vssd1 vccd1 vccd1 _20568_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10321_ _10269_/A _20713_/Q _10279_/A _20723_/Q vssd1 vssd1 vccd1 vccd1 _10321_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_166_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20499_ _20929_/CLK _20499_/D repeater267/X vssd1 vssd1 vccd1 vccd1 _20499_/Q sky130_fd_sc_hd__dfrtp_2
X_13040_ _13040_/A vssd1 vssd1 vccd1 vccd1 _13040_/X sky130_fd_sc_hd__buf_1
X_10252_ _21351_/Q vssd1 vssd1 vccd1 vccd1 _10267_/A sky130_fd_sc_hd__inv_2
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19018__S _19019_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10183_ _10183_/A vssd1 vssd1 vccd1 vccd1 _10183_/X sky130_fd_sc_hd__buf_1
XANTENNA__16231__A _16231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17046__B _17046_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input39_A HWDATA[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14991_ _14991_/A vssd1 vssd1 vccd1 vccd1 _14991_/Y sky130_fd_sc_hd__inv_2
XFILLER_219_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16730_ _20992_/Q _11998_/B _11999_/B vssd1 vssd1 vccd1 vccd1 _16730_/X sky130_fd_sc_hd__a21bo_1
X_13942_ _20635_/Q vssd1 vssd1 vccd1 vccd1 _13942_/Y sky130_fd_sc_hd__inv_2
XFILLER_247_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16661_ _16661_/A _18950_/X vssd1 vssd1 vccd1 vccd1 _19864_/D sky130_fd_sc_hd__and2_1
XFILLER_207_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13873_ _20302_/Q vssd1 vssd1 vccd1 vccd1 _13876_/C sky130_fd_sc_hd__inv_2
XFILLER_47_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15612_ _15618_/A vssd1 vssd1 vccd1 vccd1 _15619_/A sky130_fd_sc_hd__inv_2
X_18400_ _18399_/X _10109_/Y _18879_/S vssd1 vssd1 vccd1 vccd1 _18400_/X sky130_fd_sc_hd__mux2_1
X_12824_ _12842_/A vssd1 vssd1 vccd1 vccd1 _12824_/X sky130_fd_sc_hd__buf_1
X_19380_ _19776_/CLK _19380_/D vssd1 vssd1 vccd1 vccd1 _19380_/Q sky130_fd_sc_hd__dfxtp_1
X_16592_ _16592_/A vssd1 vssd1 vccd1 vccd1 _19118_/S sky130_fd_sc_hd__inv_2
XFILLER_62_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18331_ _18330_/X _14590_/A _18748_/S vssd1 vssd1 vccd1 vccd1 _18331_/X sky130_fd_sc_hd__mux2_1
X_15543_ _15553_/A vssd1 vssd1 vccd1 vccd1 _15543_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__10617__B2 _20742_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12755_ _17083_/A _12887_/A vssd1 vssd1 vccd1 vccd1 _12783_/A sky130_fd_sc_hd__or2_1
XANTENNA__18592__S _18879_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_repeater178_A _18874_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20263__RESET_B repeater264/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11706_ _21075_/Q _11704_/X _11565_/X _11705_/X vssd1 vssd1 vccd1 vccd1 _21075_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18262_ _18848_/A0 _14147_/Y _18902_/S vssd1 vssd1 vccd1 vccd1 _18262_/X sky130_fd_sc_hd__mux2_1
XFILLER_203_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15474_ _19780_/Q _15468_/X _15473_/X _15471_/X vssd1 vssd1 vccd1 vccd1 _19780_/D
+ sky130_fd_sc_hd__a22o_1
X_12686_ _12707_/A vssd1 vssd1 vccd1 vccd1 _12686_/X sky130_fd_sc_hd__buf_1
XPHY_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14425_ _14424_/Y _20215_/Q _14378_/A _14425_/B2 vssd1 vssd1 vccd1 vccd1 _14425_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__20699__CLK _21342_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17213_ _17573_/A vssd1 vssd1 vccd1 vccd1 _18045_/A sky130_fd_sc_hd__clkbuf_2
X_11637_ _11637_/A vssd1 vssd1 vccd1 vccd1 _18983_/S sky130_fd_sc_hd__clkbuf_4
X_18193_ _18192_/X _10099_/Y _18644_/S vssd1 vssd1 vccd1 vccd1 _18193_/X sky130_fd_sc_hd__mux2_1
XPHY_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17144_ _17134_/Y _17175_/B _17137_/Y _17177_/B _17143_/X vssd1 vssd1 vccd1 vccd1
+ _17144_/X sky130_fd_sc_hd__o221a_1
XFILLER_11_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14356_ _14501_/A _14500_/A _14499_/A _14496_/A vssd1 vssd1 vccd1 vccd1 _14362_/C
+ sky130_fd_sc_hd__or4_4
XPHY_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21469__RESET_B repeater204/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11568_ _11739_/A vssd1 vssd1 vccd1 vccd1 _11568_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13319__B1 _13245_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13307_ _13321_/A vssd1 vssd1 vccd1 vccd1 _13307_/X sky130_fd_sc_hd__buf_1
X_17075_ _20252_/Q vssd1 vssd1 vccd1 vccd1 _17075_/Y sky130_fd_sc_hd__inv_2
X_10519_ _20690_/Q vssd1 vssd1 vccd1 vccd1 _18034_/A sky130_fd_sc_hd__inv_2
XANTENNA__10454__A _20696_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14287_ _15357_/B vssd1 vssd1 vccd1 vccd1 _14779_/B sky130_fd_sc_hd__buf_1
X_11499_ _21151_/Q vssd1 vssd1 vccd1 vccd1 _16548_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_226_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16026_ _19523_/Q _16021_/X _15764_/X _16023_/X vssd1 vssd1 vccd1 vccd1 _19523_/D
+ sky130_fd_sc_hd__a22o_1
X_13238_ _20573_/Q _13233_/X _13032_/X _13234_/X vssd1 vssd1 vccd1 vccd1 _20573_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_124_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21051__RESET_B repeater226/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13169_ _13710_/A vssd1 vssd1 vccd1 vccd1 _13169_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18767__S _18835_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17977_ _17977_/A _17978_/B vssd1 vssd1 vccd1 vccd1 _17977_/Y sky130_fd_sc_hd__nor2_1
X_19716_ _20432_/CLK _19716_/D vssd1 vssd1 vccd1 vccd1 _19716_/Q sky130_fd_sc_hd__dfxtp_1
X_16928_ _16931_/B _16927_/Y _16915_/X vssd1 vssd1 vccd1 vccd1 _16928_/X sky130_fd_sc_hd__o21a_1
XANTENNA__17233__A1 _18907_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17233__B2 _17232_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19647_ _21021_/CLK _19647_/D vssd1 vssd1 vccd1 vccd1 _19647_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16859_ _16863_/B _16858_/Y _16831_/X vssd1 vssd1 vccd1 vccd1 _16859_/X sky130_fd_sc_hd__o21a_1
XFILLER_81_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19578_ _21449_/CLK _19578_/D vssd1 vssd1 vccd1 vccd1 _19578_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_240_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10608__B2 _20758_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18529_ _18528_/X _20193_/Q _18748_/S vssd1 vssd1 vccd1 vccd1 _18529_/X sky130_fd_sc_hd__mux2_1
XFILLER_179_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13005__A _13012_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13558__B1 _13557_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21471_ _21477_/CLK _21471_/D repeater204/X vssd1 vssd1 vccd1 vccd1 _21471_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_193_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20422_ _20422_/CLK _20422_/D repeater271/X vssd1 vssd1 vccd1 vccd1 _20422_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_135_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12781__A1 _20790_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20353_ _20476_/CLK _20353_/D repeater279/X vssd1 vssd1 vccd1 vccd1 _20353_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_162_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_121_HCLK clkbuf_opt_3_HCLK/A vssd1 vssd1 vccd1 vccd1 _20972_/CLK sky130_fd_sc_hd__clkbuf_16
X_20284_ _20661_/CLK _20284_/D repeater263/X vssd1 vssd1 vccd1 vccd1 _20284_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_162_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18677__S _18928_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18421__A0 _18848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20703__RESET_B repeater210/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_232_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10870_ _21264_/Q _10864_/X _09685_/X _10866_/X vssd1 vssd1 vccd1 vccd1 _21264_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_232_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12540_ _11307_/B _12524_/X _11544_/B _12528_/A vssd1 vssd1 vccd1 vccd1 _20902_/D
+ sky130_fd_sc_hd__o22ai_1
XPHY_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12471_ _12471_/A _12486_/A vssd1 vssd1 vccd1 vccd1 _12472_/B sky130_fd_sc_hd__or2_1
XFILLER_200_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14210_ _20272_/Q _14209_/Y _14205_/X _14083_/B vssd1 vssd1 vccd1 vccd1 _20272_/D
+ sky130_fd_sc_hd__o211a_1
X_11422_ _11363_/A _11420_/X _11365_/A _11421_/X vssd1 vssd1 vccd1 vccd1 _21179_/D
+ sky130_fd_sc_hd__o22a_1
X_15190_ _15074_/A _15074_/B _15188_/Y _15179_/X vssd1 vssd1 vccd1 vccd1 _20060_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_193_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14141_ _20551_/Q _14090_/A _20547_/Q _14086_/A _14140_/X vssd1 vssd1 vccd1 vccd1
+ _14155_/A sky130_fd_sc_hd__o221a_1
X_11353_ _11375_/A _11390_/D _11390_/C _11390_/B vssd1 vssd1 vccd1 vccd1 _16595_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_152_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10304_ _20710_/Q vssd1 vssd1 vccd1 vccd1 _10304_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19957__RESET_B repeater184/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14072_ _14072_/A _14072_/B vssd1 vssd1 vccd1 vccd1 _14225_/A sky130_fd_sc_hd__or2_1
X_11284_ _20905_/Q _11284_/B _11290_/C _11299_/D vssd1 vssd1 vccd1 vccd1 _12500_/A
+ sky130_fd_sc_hd__nor4_2
XFILLER_152_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13023_ _20680_/Q _13019_/X _12853_/X _13021_/X vssd1 vssd1 vccd1 vccd1 _20680_/D
+ sky130_fd_sc_hd__a22o_1
X_17900_ _17900_/A _17938_/B vssd1 vssd1 vccd1 vccd1 _17900_/Y sky130_fd_sc_hd__nor2_1
X_10235_ _21368_/Q vssd1 vssd1 vccd1 vccd1 _10283_/A sky130_fd_sc_hd__inv_2
X_18880_ _18879_/X _16753_/B _18880_/S vssd1 vssd1 vccd1 vccd1 _18880_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17831_ _20820_/Q vssd1 vssd1 vccd1 vccd1 _17831_/Y sky130_fd_sc_hd__inv_2
X_10166_ _10166_/A vssd1 vssd1 vccd1 vccd1 _10166_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_output145_A _21135_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18587__S _18907_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17762_ _19613_/Q vssd1 vssd1 vccd1 vccd1 _17762_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14974_ _20101_/Q _14972_/Y _14973_/X _14880_/B vssd1 vssd1 vccd1 vccd1 _20101_/D
+ sky130_fd_sc_hd__o211a_1
X_10097_ _21402_/Q _10093_/Y _21386_/Q _10094_/Y _10096_/X vssd1 vssd1 vccd1 vccd1
+ _10098_/D sky130_fd_sc_hd__o221a_1
X_19501_ _20327_/CLK _19501_/D vssd1 vssd1 vccd1 vccd1 _19501_/Q sky130_fd_sc_hd__dfxtp_1
X_16713_ _19900_/Q _14240_/B _14241_/B vssd1 vssd1 vccd1 vccd1 _16713_/X sky130_fd_sc_hd__a21bo_1
XFILLER_47_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13925_ _20643_/Q vssd1 vssd1 vccd1 vccd1 _13925_/Y sky130_fd_sc_hd__inv_2
X_17693_ _19580_/Q vssd1 vssd1 vccd1 vccd1 _17693_/Y sky130_fd_sc_hd__inv_2
XFILLER_208_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19432_ _20137_/CLK _19432_/D vssd1 vssd1 vccd1 vccd1 _19432_/Q sky130_fd_sc_hd__dfxtp_1
X_16644_ _19857_/Q _15291_/B _15292_/B vssd1 vssd1 vccd1 vccd1 _16644_/X sky130_fd_sc_hd__a21bo_1
X_13856_ _20305_/Q vssd1 vssd1 vccd1 vccd1 _13857_/A sky130_fd_sc_hd__inv_2
XANTENNA__12648__B _12815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12807_ _20774_/Q _12803_/X _11741_/X _12804_/X vssd1 vssd1 vccd1 vccd1 _20774_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_222_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19363_ _21001_/CLK _19363_/D vssd1 vssd1 vccd1 vccd1 _19363_/Q sky130_fd_sc_hd__dfxtp_1
X_16575_ _16683_/A _19997_/Q _16521_/B _16574_/X vssd1 vssd1 vccd1 vccd1 _16575_/Y
+ sky130_fd_sc_hd__a31oi_4
X_13787_ _20197_/Q vssd1 vssd1 vccd1 vccd1 _14586_/A sky130_fd_sc_hd__inv_2
X_10999_ _11008_/B vssd1 vssd1 vccd1 vccd1 _15396_/B sky130_fd_sc_hd__buf_1
X_18314_ _18313_/X _10778_/A _18898_/S vssd1 vssd1 vccd1 vccd1 _18314_/X sky130_fd_sc_hd__mux2_1
X_15526_ _15592_/A vssd1 vssd1 vccd1 vccd1 _15526_/X sky130_fd_sc_hd__buf_1
X_12738_ _14685_/A _12738_/B vssd1 vssd1 vccd1 vccd1 _12746_/B sky130_fd_sc_hd__or2_1
X_19294_ _19776_/CLK _19294_/D vssd1 vssd1 vccd1 vccd1 _19294_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_230_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15457_ _19787_/Q _15449_/X _15456_/X _15452_/X vssd1 vssd1 vccd1 vccd1 _19787_/D
+ sky130_fd_sc_hd__a22o_1
X_18245_ _19141_/X _20163_/Q _18249_/S vssd1 vssd1 vccd1 vccd1 _18245_/X sky130_fd_sc_hd__mux2_1
XPHY_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12669_ _20836_/Q _12662_/X _12668_/X _12664_/X vssd1 vssd1 vccd1 vccd1 _20836_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_187_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14408_ _21471_/Q _14502_/A _14406_/Y _20217_/Q _14407_/X vssd1 vssd1 vccd1 vccd1
+ _14420_/B sky130_fd_sc_hd__o221a_1
XANTENNA__15040__A _20062_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18176_ _18845_/A0 _13780_/Y _18896_/S vssd1 vssd1 vccd1 vccd1 _18176_/X sky130_fd_sc_hd__mux2_1
X_15388_ _19818_/Q _15376_/X _15343_/X _15380_/X vssd1 vssd1 vccd1 vccd1 _19818_/D
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_144_HCLK clkbuf_4_3_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20142_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_117_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14339_ _20226_/Q vssd1 vssd1 vccd1 vccd1 _14461_/B sky130_fd_sc_hd__inv_2
XANTENNA__15975__A _16237_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17127_ _19438_/Q vssd1 vssd1 vccd1 vccd1 _17127_/Y sky130_fd_sc_hd__inv_2
XFILLER_156_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21232__RESET_B repeater249/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_237_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17058_ _21042_/Q _21041_/Q _17058_/C vssd1 vssd1 vccd1 vccd1 _17058_/X sky130_fd_sc_hd__and3_1
XFILLER_116_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16009_ _16335_/A vssd1 vssd1 vccd1 vccd1 _16009_/X sky130_fd_sc_hd__clkbuf_2
X_09880_ _21440_/Q _09878_/Y _09878_/B _09879_/Y vssd1 vssd1 vccd1 vccd1 _21440_/D
+ sky130_fd_sc_hd__o22a_1
Xclkbuf_4_7_0_HCLK clkbuf_4_7_0_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_7_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__18497__S _18787_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20971_ _20971_/CLK _20971_/D repeater187/X vssd1 vssd1 vccd1 vccd1 _20971_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__18954__A1 _21082_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_214_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_214_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18706__A1 _19216_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18960__S _18962_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21454_ _21457_/CLK _21454_/D repeater245/X vssd1 vssd1 vccd1 vccd1 _21454_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_31_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20405_ _20408_/CLK _20405_/D repeater184/X vssd1 vssd1 vccd1 vccd1 _20405_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_147_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21385_ _21390_/CLK _21385_/D repeater239/X vssd1 vssd1 vccd1 vccd1 _21385_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_190_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20336_ _20951_/CLK _20336_/D repeater271/X vssd1 vssd1 vccd1 vccd1 _20336_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_134_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13703__B1 _13511_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20267_ _20293_/CLK _20267_/D repeater263/X vssd1 vssd1 vccd1 vccd1 _20267_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__20955__RESET_B repeater187/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10020_ _14813_/D vssd1 vssd1 vccd1 vccd1 _17031_/A sky130_fd_sc_hd__inv_2
XANTENNA__18642__A0 _18641_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20198_ _20626_/CLK _20198_/D repeater193/X vssd1 vssd1 vccd1 vccd1 _20198_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__13926__A1_N _20663_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18200__S _18835_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_25_HCLK clkbuf_4_9_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _21419_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_57_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11971_ _16515_/A _11978_/B vssd1 vssd1 vccd1 vccd1 _11972_/A sky130_fd_sc_hd__or2_1
XANTENNA__09686__A1 _21467_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13710_ _13710_/A vssd1 vssd1 vccd1 vccd1 _13710_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_244_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10922_ _21201_/Q vssd1 vssd1 vccd1 vccd1 _10922_/Y sky130_fd_sc_hd__inv_2
X_14690_ _14696_/A vssd1 vssd1 vccd1 vccd1 _14690_/X sky130_fd_sc_hd__buf_1
XANTENNA__12690__B1 _09645_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13641_ _20375_/Q _13639_/X _13429_/X _13640_/X vssd1 vssd1 vccd1 vccd1 _20375_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_16_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10853_ _10853_/A vssd1 vssd1 vccd1 vccd1 _10853_/X sky130_fd_sc_hd__buf_1
XANTENNA__14964__A _20497_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_232_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19031__S _19046_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16360_ _17073_/B _19888_/Q vssd1 vssd1 vccd1 vccd1 _16360_/X sky130_fd_sc_hd__or2_1
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13572_ _13572_/A vssd1 vssd1 vccd1 vccd1 _13594_/A sky130_fd_sc_hd__clkbuf_2
X_10784_ _10784_/A vssd1 vssd1 vccd1 vccd1 _10784_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_167_HCLK clkbuf_opt_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20857_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_135_HCLK_A clkbuf_4_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15311_ _19916_/Q _16632_/A _20036_/Q _15310_/A vssd1 vssd1 vccd1 vccd1 _20036_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_212_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12523_ _12523_/A vssd1 vssd1 vccd1 vccd1 _12527_/A sky130_fd_sc_hd__buf_1
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16291_ _20326_/Q vssd1 vssd1 vccd1 vccd1 _16291_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_200_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18870__S _18930_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15242_ _20485_/Q vssd1 vssd1 vccd1 vccd1 _17976_/A sky130_fd_sc_hd__inv_2
X_18030_ _18030_/A _18032_/B vssd1 vssd1 vccd1 vccd1 _18030_/Y sky130_fd_sc_hd__nor2_1
XFILLER_145_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12454_ _12427_/A _12427_/B _12453_/X _12451_/Y vssd1 vssd1 vccd1 vccd1 _20938_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_185_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11405_ _21183_/Q _11401_/X _11411_/A _11404_/X vssd1 vssd1 vccd1 vccd1 _21183_/D
+ sky130_fd_sc_hd__a22o_1
X_15173_ _15173_/A vssd1 vssd1 vccd1 vccd1 _15173_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15795__A _16016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12385_ _12109_/X _12308_/B _12350_/A _12383_/Y vssd1 vssd1 vccd1 vccd1 _20954_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_125_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20737__CLK _21342_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14124_ _20532_/Q _14072_/A _14121_/Y _20261_/Q _14123_/X vssd1 vssd1 vccd1 vccd1
+ _14124_/X sky130_fd_sc_hd__a221o_1
XFILLER_125_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11336_ _21177_/Q _21176_/Q _11346_/C vssd1 vssd1 vccd1 vccd1 _11783_/D sky130_fd_sc_hd__or3_1
X_19981_ _21242_/CLK _19981_/D repeater189/X vssd1 vssd1 vccd1 vccd1 _19981_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_180_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18932_ _21193_/Q _21144_/Q _19881_/Q vssd1 vssd1 vccd1 vccd1 _18932_/X sky130_fd_sc_hd__mux2_1
XANTENNA_repeater210_A repeater211/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14055_ _20273_/Q vssd1 vssd1 vccd1 vccd1 _14083_/A sky130_fd_sc_hd__inv_2
XFILLER_125_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11267_ _11541_/A _20913_/Q _11299_/C _11294_/A vssd1 vssd1 vccd1 vccd1 _11302_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_4_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20696__RESET_B repeater193/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13170__A1 _20601_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13006_ input53/X vssd1 vssd1 vccd1 vccd1 _13006_/X sky130_fd_sc_hd__clkbuf_4
X_10218_ _10218_/A vssd1 vssd1 vccd1 vccd1 _10223_/A sky130_fd_sc_hd__inv_2
X_18863_ _18862_/X _09746_/Y _18928_/S vssd1 vssd1 vccd1 vccd1 _18863_/X sky130_fd_sc_hd__mux2_1
X_11198_ _21213_/Q _11192_/A _10900_/X _11193_/A vssd1 vssd1 vccd1 vccd1 _21213_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_121_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20625__RESET_B repeater193/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17814_ _17814_/A vssd1 vssd1 vccd1 vccd1 _18085_/B sky130_fd_sc_hd__buf_1
X_10149_ _10149_/A _10149_/B vssd1 vssd1 vccd1 vccd1 _10196_/A sky130_fd_sc_hd__or2_1
X_18794_ _18793_/X _16483_/Y _18929_/S vssd1 vssd1 vccd1 vccd1 _18794_/X sky130_fd_sc_hd__mux2_1
X_17745_ _19413_/Q vssd1 vssd1 vccd1 vccd1 _17745_/Y sky130_fd_sc_hd__inv_2
XFILLER_236_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14957_ _14957_/A vssd1 vssd1 vccd1 vccd1 _14967_/A sky130_fd_sc_hd__inv_2
XANTENNA__19284__S1 _21017_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11563__A input63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13908_ _20661_/Q vssd1 vssd1 vccd1 vccd1 _13908_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12681__B1 _09630_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17676_ _19508_/Q vssd1 vssd1 vccd1 vccd1 _17676_/Y sky130_fd_sc_hd__inv_2
X_14888_ _20585_/Q _14838_/A _20594_/Q _14882_/A vssd1 vssd1 vccd1 vccd1 _14894_/A
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_4_15_0_HCLK clkbuf_3_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_7_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_19415_ _21273_/CLK _19415_/D vssd1 vssd1 vccd1 vccd1 _19415_/Q sky130_fd_sc_hd__dfxtp_1
X_16627_ _19842_/Q vssd1 vssd1 vccd1 vccd1 _17143_/A sky130_fd_sc_hd__inv_2
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13839_ _14639_/A vssd1 vssd1 vccd1 vccd1 _14636_/A sky130_fd_sc_hd__buf_2
XANTENNA__14422__A1 _21467_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19346_ _21453_/CLK _19346_/D vssd1 vssd1 vccd1 vccd1 _19346_/Q sky130_fd_sc_hd__dfxtp_1
X_16558_ _16738_/B _19994_/Q _16561_/A _16547_/Y _16557_/X vssd1 vssd1 vccd1 vccd1
+ _16558_/X sky130_fd_sc_hd__a32o_1
XANTENNA__21484__RESET_B repeater200/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15509_ _15519_/A vssd1 vssd1 vccd1 vccd1 _15509_/X sky130_fd_sc_hd__buf_1
X_19277_ _19709_/Q _19573_/Q _19565_/Q _19557_/Q _19280_/S0 _20122_/Q vssd1 vssd1
+ vccd1 vccd1 _19277_/X sky130_fd_sc_hd__mux4_2
XANTENNA__18780__S _18902_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16489_ _16490_/B vssd1 vssd1 vccd1 vccd1 _18249_/S sky130_fd_sc_hd__inv_2
XFILLER_148_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18228_ _20852_/Q input32/X _18236_/S vssd1 vssd1 vccd1 vccd1 _18228_/X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_57_HCLK_A clkbuf_4_14_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18159_ _18848_/A0 _17991_/Y _18666_/S vssd1 vssd1 vccd1 vccd1 _18159_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21170_ _21184_/CLK _21170_/D repeater216/X vssd1 vssd1 vccd1 vccd1 _21170_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_171_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20121_ _21452_/CLK _20121_/D repeater247/X vssd1 vssd1 vccd1 vccd1 _20121_/Q sky130_fd_sc_hd__dfrtp_2
X_09932_ _11489_/C vssd1 vssd1 vccd1 vccd1 _10908_/A sky130_fd_sc_hd__buf_1
XFILLER_98_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20052_ _20066_/CLK _20052_/D repeater281/X vssd1 vssd1 vccd1 vccd1 _20052_/Q sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_48_HCLK clkbuf_opt_4_HCLK/A vssd1 vssd1 vccd1 vccd1 _21162_/CLK sky130_fd_sc_hd__clkbuf_16
X_09863_ _09853_/X _09859_/Y _09859_/B _09862_/Y vssd1 vssd1 vccd1 vccd1 _21444_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_97_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09794_ _21458_/Q _18976_/S _18964_/X vssd1 vssd1 vccd1 vccd1 _09795_/A sky130_fd_sc_hd__a21oi_2
XFILLER_245_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrepeater152 _18902_/S vssd1 vssd1 vccd1 vccd1 _18896_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_27_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater163 _18910_/S vssd1 vssd1 vccd1 vccd1 _18907_/S sky130_fd_sc_hd__clkbuf_16
XANTENNA__18955__S _18962_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19275__S1 _21004_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrepeater174 _18885_/S vssd1 vssd1 vccd1 vccd1 _18879_/S sky130_fd_sc_hd__buf_8
XPHY_4306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater185 repeater186/X vssd1 vssd1 vccd1 vccd1 repeater185/X sky130_fd_sc_hd__buf_8
XPHY_4317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater196 repeater198/X vssd1 vssd1 vccd1 vccd1 repeater196/X sky130_fd_sc_hd__buf_8
X_20954_ _20981_/CLK _20954_/D repeater186/X vssd1 vssd1 vccd1 vccd1 _20954_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_4339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20885_ _21444_/CLK _20885_/D repeater246/X vssd1 vssd1 vccd1 vccd1 _20885_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__14413__B2 _20028_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12975__A1 _20700_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18690__S _18897_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21437_ _21438_/CLK _21437_/D repeater239/X vssd1 vssd1 vccd1 vccd1 _21437_/Q sky130_fd_sc_hd__dfrtp_1
X_12170_ _12328_/A _20357_/Q _12119_/X _20356_/Q vssd1 vssd1 vccd1 vccd1 _12170_/X
+ sky130_fd_sc_hd__a22o_1
X_21368_ _21368_/CLK _21368_/D repeater257/X vssd1 vssd1 vccd1 vccd1 _21368_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11121_ _11076_/X _11112_/X _11100_/X _11120_/X vssd1 vssd1 vccd1 vccd1 _21225_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_107_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20319_ _20322_/CLK _20319_/D repeater262/X vssd1 vssd1 vccd1 vccd1 _20319_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_174_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21299_ _21302_/CLK _21299_/D repeater209/X vssd1 vssd1 vccd1 vccd1 _21299_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_107_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11052_ _11112_/A _11113_/A _11052_/C _11052_/D vssd1 vssd1 vccd1 vccd1 _11108_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_89_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10003_ _21416_/Q vssd1 vssd1 vccd1 vccd1 _10003_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19026__S _19026_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15860_ _19599_/Q _15856_/X _15793_/X _15857_/X vssd1 vssd1 vccd1 vccd1 _19599_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__20036__RESET_B repeater220/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input21_A HADDR[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14811_ _20118_/Q _14311_/X _14794_/A _14810_/X vssd1 vssd1 vccd1 vccd1 _20118_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_218_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18865__S _18930_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15791_ _16012_/A vssd1 vssd1 vccd1 vccd1 _15791_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_190_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19266__S1 _21006_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17530_ _20120_/Q _17446_/X _17527_/X _17528_/X _17529_/Y vssd1 vssd1 vccd1 vccd1
+ _17530_/X sky130_fd_sc_hd__o221a_1
XFILLER_233_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14742_ _14744_/A _14561_/A _15799_/A vssd1 vssd1 vccd1 vccd1 _14742_/X sky130_fd_sc_hd__o21a_1
X_11954_ _19109_/X _11128_/X _11142_/X vssd1 vssd1 vccd1 vccd1 _11955_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__17989__B _17989_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10905_ _21249_/Q _09919_/B _11021_/B vssd1 vssd1 vccd1 vccd1 _21249_/D sky130_fd_sc_hd__a21o_1
XFILLER_244_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17461_ _17453_/Y _17136_/A _17454_/Y _17376_/X _17460_/X vssd1 vssd1 vccd1 vccd1
+ _17461_/X sky130_fd_sc_hd__o221a_2
XFILLER_32_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14673_ _14673_/A vssd1 vssd1 vccd1 vccd1 _14673_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14404__A1 _14403_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11885_ _11885_/A _11885_/B vssd1 vssd1 vccd1 vccd1 _11886_/A sky130_fd_sc_hd__nand2_1
XFILLER_33_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output108_A _17805_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19200_ _17769_/Y _17770_/Y _17771_/Y _17772_/Y _20130_/Q _20131_/Q vssd1 vssd1 vccd1
+ vccd1 _19200_/X sky130_fd_sc_hd__mux4_2
XFILLER_44_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16412_ _19329_/Q _16406_/X _16204_/X _16408_/X vssd1 vssd1 vccd1 vccd1 _19329_/D
+ sky130_fd_sc_hd__a22o_1
X_13624_ _20384_/Q _13619_/X _13479_/X _13620_/X vssd1 vssd1 vccd1 vccd1 _20384_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_177_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10836_ _10836_/A vssd1 vssd1 vccd1 vccd1 _10836_/Y sky130_fd_sc_hd__inv_2
XFILLER_220_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17392_ _17386_/Y _17387_/X _11508_/Y _17378_/X _17391_/X vssd1 vssd1 vccd1 vccd1
+ _17392_/X sky130_fd_sc_hd__o221a_1
XFILLER_186_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19131_ _19127_/X _19128_/X _19129_/X _19130_/X _21018_/Q _21019_/Q vssd1 vssd1 vccd1
+ vccd1 _19131_/X sky130_fd_sc_hd__mux4_2
X_16343_ _19366_/Q _16334_/X _16342_/X _16336_/X vssd1 vssd1 vccd1 vccd1 _19366_/D
+ sky130_fd_sc_hd__a22o_1
X_13555_ input55/X vssd1 vssd1 vccd1 vccd1 _13555_/X sky130_fd_sc_hd__buf_4
XANTENNA_repeater160_A _18841_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10767_ _10767_/A _10767_/B vssd1 vssd1 vccd1 vccd1 _10815_/A sky130_fd_sc_hd__or2_1
X_12506_ _12506_/A _12506_/B vssd1 vssd1 vccd1 vccd1 _12506_/X sky130_fd_sc_hd__or2_1
XFILLER_201_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19062_ _21189_/Q _21131_/Q _19910_/Q vssd1 vssd1 vccd1 vccd1 _19062_/X sky130_fd_sc_hd__mux2_1
XANTENNA__19972__RESET_B repeater184/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16274_ _19398_/Q _16269_/X _16127_/X _16270_/X vssd1 vssd1 vccd1 vccd1 _19398_/D
+ sky130_fd_sc_hd__a22o_1
X_13486_ _20451_/Q _13481_/X _13485_/X _13483_/X vssd1 vssd1 vccd1 vccd1 _20451_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_73_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10698_ _21323_/Q _10697_/Y _10712_/A _10653_/B vssd1 vssd1 vccd1 vccd1 _21323_/D
+ sky130_fd_sc_hd__o211a_1
X_15225_ _20479_/Q vssd1 vssd1 vccd1 vccd1 _17896_/A sky130_fd_sc_hd__inv_2
X_18013_ _18149_/X _17954_/X _18162_/X _17955_/X vssd1 vssd1 vccd1 vccd1 _18014_/D
+ sky130_fd_sc_hd__a22o_2
XFILLER_139_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12437_ _20945_/Q _20944_/Q _12437_/C vssd1 vssd1 vccd1 vccd1 _12437_/X sky130_fd_sc_hd__and3_1
X_15156_ _15154_/Y _20045_/Q _20449_/Q _15074_/A _15155_/X vssd1 vssd1 vccd1 vccd1
+ _15157_/D sky130_fd_sc_hd__o221a_1
XANTENNA__18854__A0 _17079_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12368_ _12036_/X _12317_/B _12364_/X _12366_/Y vssd1 vssd1 vccd1 vccd1 _20964_/D
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__15668__B1 _15585_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20806__RESET_B repeater235/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14107_ _14102_/Y _20290_/Q _20539_/Q _14103_/X _14106_/X vssd1 vssd1 vccd1 vccd1
+ _14120_/A sky130_fd_sc_hd__o221a_1
X_11319_ _19882_/Q vssd1 vssd1 vccd1 vccd1 _12515_/A sky130_fd_sc_hd__buf_1
XANTENNA__11558__A input64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19964_ _20413_/CLK _19964_/D repeater184/X vssd1 vssd1 vccd1 vccd1 _19964_/Q sky130_fd_sc_hd__dfrtp_1
X_15087_ _15087_/A _15165_/A vssd1 vssd1 vccd1 vccd1 _15088_/B sky130_fd_sc_hd__or2_2
X_12299_ _20933_/Q _12297_/Y _12298_/Y _20529_/Q vssd1 vssd1 vccd1 vccd1 _12299_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_234_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13143__A1 _20614_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14038_ _14031_/A _14031_/B _20291_/Q _13976_/D _13980_/X vssd1 vssd1 vccd1 vccd1
+ _20291_/D sky130_fd_sc_hd__o221a_1
X_18915_ _18914_/X _21408_/Q _20869_/Q vssd1 vssd1 vccd1 vccd1 _18915_/X sky130_fd_sc_hd__mux2_1
X_19895_ _21191_/CLK _19895_/D repeater224/X vssd1 vssd1 vccd1 vccd1 _19895_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_68_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18846_ _18845_/X _14397_/Y _18897_/S vssd1 vssd1 vccd1 vccd1 _18846_/X sky130_fd_sc_hd__mux2_1
XFILLER_227_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10901__B1 _10900_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18777_ _18845_/A0 _13813_/Y _18896_/S vssd1 vssd1 vccd1 vccd1 _18777_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18775__S _18775_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15989_ _19541_/Q _15986_/X _15969_/X _15988_/X vssd1 vssd1 vccd1 vccd1 _19541_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19257__S1 _20131_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17728_ _17720_/Y _17301_/X _17723_/X _17727_/X vssd1 vssd1 vccd1 vccd1 _17728_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_236_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19925__CLK _21342_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17659_ _17889_/A vssd1 vssd1 vccd1 vccd1 _17839_/A sky130_fd_sc_hd__buf_1
XFILLER_90_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20670_ _21294_/CLK _20670_/D repeater211/X vssd1 vssd1 vccd1 vccd1 _20670_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_211_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10417__C1 _10375_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19329_ _19834_/CLK _19329_/D vssd1 vssd1 vccd1 vccd1 _19329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13013__A _13013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19193__S0 _19280_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18845__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21222_ _21222_/CLK _21222_/D repeater235/X vssd1 vssd1 vccd1 vccd1 _21222_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_144_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21153_ _21429_/CLK _21153_/D repeater231/X vssd1 vssd1 vccd1 vccd1 _21153_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_144_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20104_ _20107_/CLK _20104_/D repeater259/X vssd1 vssd1 vccd1 vccd1 _20104_/Q sky130_fd_sc_hd__dfrtp_1
X_09915_ _09895_/Y _09897_/Y _21257_/Q _17024_/A _09914_/X vssd1 vssd1 vccd1 vccd1
+ _09915_/X sky130_fd_sc_hd__o221a_1
X_21084_ _21087_/CLK _21084_/D repeater228/X vssd1 vssd1 vccd1 vccd1 _21084_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_120_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18073__A1 _18408_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09846_ _09876_/A _09878_/A _09846_/C vssd1 vssd1 vccd1 vccd1 _09871_/A sky130_fd_sc_hd__or3_4
XFILLER_100_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20035_ _21421_/CLK _20035_/D repeater239/X vssd1 vssd1 vccd1 vccd1 _20035_/Q sky130_fd_sc_hd__dfrtp_1
X_09777_ _09777_/A _09777_/B vssd1 vssd1 vccd1 vccd1 _09777_/X sky130_fd_sc_hd__or2_1
XANTENNA__19248__S1 _20131_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18685__S _18841_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20937_ _20937_/CLK _20937_/D repeater277/X vssd1 vssd1 vccd1 vccd1 _20937_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_4169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__21335__RESET_B repeater203/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17584__B1 _18761_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_241_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11931__A _21007_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11670_ _21090_/Q vssd1 vssd1 vccd1 vccd1 _11670_/Y sky130_fd_sc_hd__inv_2
XPHY_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20868_ _21452_/CLK _20868_/D repeater247/X vssd1 vssd1 vccd1 vccd1 _20868_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10621_ _21335_/Q _10618_/Y _21324_/Q _10619_/Y _10620_/X vssd1 vssd1 vccd1 vccd1
+ _10622_/D sky130_fd_sc_hd__o221a_1
XPHY_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13070__B1 _12920_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20799_ _21407_/CLK _20799_/D repeater255/X vssd1 vssd1 vccd1 vccd1 _20799_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13340_ _13352_/A vssd1 vssd1 vccd1 vccd1 _13340_/X sky130_fd_sc_hd__buf_1
XFILLER_183_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10552_ _10702_/A _10701_/C _10552_/C _10552_/D vssd1 vssd1 vccd1 vccd1 _10650_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_155_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15898__B1 _15788_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13271_ _20560_/Q _13264_/X _13270_/X _13268_/X vssd1 vssd1 vccd1 vccd1 _20560_/D
+ sky130_fd_sc_hd__a22o_1
X_10483_ _10759_/A _20671_/Q _21280_/Q _10479_/Y _10482_/X vssd1 vssd1 vccd1 vccd1
+ _10496_/B sky130_fd_sc_hd__o221a_1
XANTENNA_clkbuf_leaf_40_HCLK_A clkbuf_4_11_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20970__RESET_B repeater187/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15010_ _20085_/Q _15009_/Y _15006_/B _14978_/X vssd1 vssd1 vccd1 vccd1 _20085_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__19184__S0 _19280_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12222_ _20510_/Q vssd1 vssd1 vccd1 vccd1 _12222_/Y sky130_fd_sc_hd__inv_2
XANTENNA_input69_A HWDATA[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12153_ _20353_/Q vssd1 vssd1 vccd1 vccd1 _12153_/Y sky130_fd_sc_hd__inv_2
XFILLER_162_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20217__RESET_B repeater202/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11104_ _11104_/A vssd1 vssd1 vccd1 vccd1 _11105_/B sky130_fd_sc_hd__inv_2
XFILLER_96_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12084_ _20368_/Q vssd1 vssd1 vccd1 vccd1 _17539_/A sky130_fd_sc_hd__inv_2
X_16961_ _16966_/B _16960_/X _16939_/X vssd1 vssd1 vccd1 vccd1 _16961_/X sky130_fd_sc_hd__o21a_1
XFILLER_96_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18700_ _18699_/X _17707_/Y _18910_/S vssd1 vssd1 vccd1 vccd1 _18700_/X sky130_fd_sc_hd__mux2_1
X_15912_ _15912_/A vssd1 vssd1 vccd1 vccd1 _15912_/X sky130_fd_sc_hd__buf_1
X_11035_ _19963_/Q _19962_/Q _16930_/A vssd1 vssd1 vccd1 vccd1 _16937_/A sky130_fd_sc_hd__or3_4
XFILLER_77_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11687__A1 _21085_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19680_ _19812_/CLK _19680_/D vssd1 vssd1 vccd1 vccd1 _19680_/Q sky130_fd_sc_hd__dfxtp_1
X_16892_ _16892_/A vssd1 vssd1 vccd1 vccd1 _16892_/Y sky130_fd_sc_hd__inv_2
XFILLER_209_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18631_ _18845_/A0 _13768_/Y _18896_/S vssd1 vssd1 vccd1 vccd1 _18631_/X sky130_fd_sc_hd__mux2_1
XFILLER_237_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15843_ _19609_/Q _15841_/X _09832_/X _15842_/X vssd1 vssd1 vccd1 vccd1 _19609_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_76_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18595__S _18874_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14625__A1 _20193_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19239__S1 _20131_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18562_ _18561_/X _14575_/A _18748_/S vssd1 vssd1 vccd1 vccd1 _18562_/X sky130_fd_sc_hd__mux2_2
X_12986_ _13020_/A vssd1 vssd1 vccd1 vccd1 _13013_/A sky130_fd_sc_hd__clkbuf_2
X_15774_ _15774_/A vssd1 vssd1 vccd1 vccd1 _15774_/X sky130_fd_sc_hd__buf_1
XFILLER_218_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20925__CLK _20930_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17513_ _19626_/Q vssd1 vssd1 vccd1 vccd1 _17513_/Y sky130_fd_sc_hd__inv_2
X_14725_ _20147_/Q _14723_/X _13707_/X _14724_/X vssd1 vssd1 vccd1 vccd1 _20147_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_233_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18493_ _17079_/Y _12067_/Y _18908_/S vssd1 vssd1 vccd1 vccd1 _18493_/X sky130_fd_sc_hd__mux2_1
X_11937_ _21009_/Q vssd1 vssd1 vccd1 vccd1 _11940_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_32_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12937__A _12961_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14389__B1 _21467_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_233_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17444_ _20142_/Q vssd1 vssd1 vccd1 vccd1 _17444_/Y sky130_fd_sc_hd__inv_2
X_14656_ _14656_/A vssd1 vssd1 vccd1 vccd1 _19124_/S sky130_fd_sc_hd__inv_2
X_11868_ _11863_/X _11864_/X _10964_/X vssd1 vssd1 vccd1 vccd1 _11868_/X sky130_fd_sc_hd__o21a_1
XANTENNA__21005__RESET_B repeater235/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_221_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13607_ _13633_/A vssd1 vssd1 vccd1 vccd1 _13626_/A sky130_fd_sc_hd__clkbuf_2
X_10819_ _21290_/Q _10818_/Y _10812_/X _10767_/B vssd1 vssd1 vccd1 vccd1 _21290_/D
+ sky130_fd_sc_hd__o211a_1
X_17375_ _21082_/Q vssd1 vssd1 vccd1 vccd1 _17375_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17327__B1 _18847_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14587_ _14587_/A _14587_/B vssd1 vssd1 vccd1 vccd1 _14613_/A sky130_fd_sc_hd__or2_1
X_11799_ _21218_/Q vssd1 vssd1 vccd1 vccd1 _11817_/A sky130_fd_sc_hd__inv_2
XFILLER_229_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19114_ _16594_/Y _10985_/Y _19118_/S vssd1 vssd1 vccd1 vccd1 _19114_/X sky130_fd_sc_hd__mux2_2
XFILLER_201_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16326_ _16334_/A vssd1 vssd1 vccd1 vccd1 _16326_/X sky130_fd_sc_hd__buf_1
X_13538_ input62/X vssd1 vssd1 vccd1 vccd1 _13538_/X sky130_fd_sc_hd__buf_4
X_19045_ _16804_/X _20824_/Q _19046_/S vssd1 vssd1 vccd1 vccd1 _19931_/D sky130_fd_sc_hd__mux2_1
X_13469_ _20459_/Q _13466_/X _13280_/X _13467_/X vssd1 vssd1 vccd1 vccd1 _20459_/D
+ sky130_fd_sc_hd__a22o_1
X_16257_ _19409_/Q _16255_/X _16120_/X _16256_/X vssd1 vssd1 vccd1 vccd1 _19409_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_173_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19175__S0 _19280_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15208_ _15208_/A vssd1 vssd1 vccd1 vccd1 _15208_/Y sky130_fd_sc_hd__inv_2
X_16188_ _16188_/A vssd1 vssd1 vccd1 vccd1 _16188_/X sky130_fd_sc_hd__buf_1
X_15139_ _15137_/Y _20069_/Q _15138_/Y _20055_/Q vssd1 vssd1 vccd1 vccd1 _15139_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_114_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19947_ _20841_/CLK _19947_/D repeater251/X vssd1 vssd1 vccd1 vccd1 _19947_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_141_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09700_ input38/X vssd1 vssd1 vccd1 vccd1 _15354_/A sky130_fd_sc_hd__buf_2
XFILLER_229_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19878_ _21193_/CLK _21126_/Q repeater223/X vssd1 vssd1 vccd1 vccd1 _19878_/Q sky130_fd_sc_hd__dfrtp_1
X_09631_ _21482_/Q _09620_/X _09630_/X _09624_/X vssd1 vssd1 vccd1 vccd1 _21482_/D
+ sky130_fd_sc_hd__a22o_1
X_18829_ _18828_/X _19251_/X _18930_/S vssd1 vssd1 vccd1 vccd1 _18829_/X sky130_fd_sc_hd__mux2_2
XFILLER_110_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16319__A _16319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20722_ _20724_/CLK _20722_/D repeater264/X vssd1 vssd1 vccd1 vccd1 _20722_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20653_ _20657_/CLK _20653_/D repeater197/X vssd1 vssd1 vccd1 vccd1 _20653_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_149_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20799__RESET_B repeater255/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20584_ _20946_/CLK _20584_/D repeater274/X vssd1 vssd1 vccd1 vccd1 _20584_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_192_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20728__RESET_B repeater257/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19166__S0 _20123_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12563__C1 _11795_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15893__A _16237_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21205_ _21207_/CLK _21205_/D repeater256/X vssd1 vssd1 vccd1 vccd1 _21205_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_151_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21136_ _21147_/CLK _21136_/D repeater215/X vssd1 vssd1 vccd1 vccd1 _21136_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_132_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21067_ _21087_/CLK _21067_/D repeater228/X vssd1 vssd1 vccd1 vccd1 _21067_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_59_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12866__B1 _12699_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20018_ _21417_/CLK _20018_/D repeater230/X vssd1 vssd1 vccd1 vccd1 _20018_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_247_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09829_ _09829_/A vssd1 vssd1 vccd1 vccd1 _09829_/X sky130_fd_sc_hd__buf_1
XFILLER_46_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12840_ _20758_/Q _12835_/X _09628_/X _12836_/X vssd1 vssd1 vccd1 vccd1 _20758_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_227_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12771_ _12777_/A vssd1 vssd1 vccd1 vccd1 _12771_/X sky130_fd_sc_hd__buf_1
XFILLER_215_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14510_ _14510_/A vssd1 vssd1 vccd1 vccd1 _14510_/Y sky130_fd_sc_hd__inv_2
XFILLER_202_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11722_ _21067_/Q _11720_/X _11565_/X _11721_/X vssd1 vssd1 vccd1 vccd1 _21067_/D
+ sky130_fd_sc_hd__a22o_1
X_15490_ _15490_/A _16481_/A vssd1 vssd1 vccd1 vccd1 _16229_/C sky130_fd_sc_hd__or2_2
XFILLER_203_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14441_ _14465_/A _20026_/Q _21481_/Q _14461_/A _14440_/X vssd1 vssd1 vccd1 vccd1
+ _14449_/B sky130_fd_sc_hd__o221a_1
X_11653_ _13327_/A _13327_/B _13047_/C vssd1 vssd1 vccd1 vccd1 _17157_/D sky130_fd_sc_hd__or3_4
XPHY_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13043__B1 _12879_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16780__A1 _16777_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10604_ _10700_/A _20738_/Q _10654_/A _20753_/Q _10603_/X vssd1 vssd1 vccd1 vccd1
+ _10605_/D sky130_fd_sc_hd__o221a_1
XFILLER_168_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14372_ _14460_/B _14372_/B vssd1 vssd1 vccd1 vccd1 _14480_/A sky130_fd_sc_hd__or2_1
X_17160_ _20893_/Q vssd1 vssd1 vccd1 vccd1 _17160_/Y sky130_fd_sc_hd__inv_2
XPHY_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11584_ _21244_/Q _11584_/B _11584_/C vssd1 vssd1 vccd1 vccd1 _11590_/B sky130_fd_sc_hd__or3_1
XFILLER_196_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16111_ _16121_/A vssd1 vssd1 vccd1 vccd1 _16111_/X sky130_fd_sc_hd__clkbuf_2
X_13323_ _20533_/Q _13321_/X _13166_/X _13322_/X vssd1 vssd1 vccd1 vccd1 _20533_/D
+ sky130_fd_sc_hd__a22o_1
X_10535_ _21339_/Q vssd1 vssd1 vccd1 vccd1 _10574_/C sky130_fd_sc_hd__inv_2
XANTENNA__13588__A _13594_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17091_ _21309_/Q _20772_/Q vssd1 vssd1 vccd1 vccd1 _17091_/X sky130_fd_sc_hd__and2_2
XANTENNA__19620__CLK _21452_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19157__S0 _19285_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16042_ _16042_/A vssd1 vssd1 vccd1 vccd1 _16042_/X sky130_fd_sc_hd__buf_1
X_13254_ _13600_/A vssd1 vssd1 vccd1 vccd1 _13254_/X sky130_fd_sc_hd__clkbuf_2
X_10466_ _20672_/Q vssd1 vssd1 vccd1 vccd1 _10466_/Y sky130_fd_sc_hd__inv_2
XFILLER_171_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12205_ _12205_/A _12205_/B _12190_/X _12204_/X vssd1 vssd1 vccd1 vccd1 _12373_/A
+ sky130_fd_sc_hd__or4bb_4
X_13185_ _13185_/A _13185_/B _16525_/C vssd1 vssd1 vccd1 vccd1 _13185_/X sky130_fd_sc_hd__or3_1
X_10397_ _10397_/A vssd1 vssd1 vccd1 vccd1 _10397_/X sky130_fd_sc_hd__buf_2
XANTENNA__20051__RESET_B repeater281/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19801_ _19820_/CLK _19801_/D vssd1 vssd1 vccd1 vccd1 _19801_/Q sky130_fd_sc_hd__dfxtp_1
X_12136_ _20975_/Q _12131_/Y _12328_/A _20389_/Q _12135_/X vssd1 vssd1 vccd1 vccd1
+ _12144_/C sky130_fd_sc_hd__o221a_1
XFILLER_96_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17993_ _18213_/X _17928_/X _18156_/X _17960_/X vssd1 vssd1 vccd1 vccd1 _17993_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_215_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19732_ _19777_/CLK _19732_/D vssd1 vssd1 vccd1 vccd1 _19732_/Q sky130_fd_sc_hd__dfxtp_1
X_12067_ _20379_/Q vssd1 vssd1 vccd1 vccd1 _12067_/Y sky130_fd_sc_hd__inv_2
X_16944_ _19965_/Q vssd1 vssd1 vccd1 vccd1 _16944_/Y sky130_fd_sc_hd__inv_2
XFILLER_111_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11018_ _21246_/Q vssd1 vssd1 vccd1 vccd1 _17027_/A sky130_fd_sc_hd__inv_2
X_19663_ _21021_/CLK _19663_/D vssd1 vssd1 vccd1 vccd1 _19663_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16875_ _19948_/Q vssd1 vssd1 vccd1 vccd1 _16875_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_237_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18614_ _18613_/X _16785_/Y _18667_/S vssd1 vssd1 vccd1 vccd1 _18614_/X sky130_fd_sc_hd__mux2_1
X_15826_ _19617_/Q _15824_/X _09832_/X _15825_/X vssd1 vssd1 vccd1 vccd1 _19617_/D
+ sky130_fd_sc_hd__a22o_1
X_19594_ _19626_/CLK _19594_/D vssd1 vssd1 vccd1 vccd1 _19594_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_237_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18545_ _18544_/X _10610_/Y _18775_/S vssd1 vssd1 vccd1 vccd1 _18545_/X sky130_fd_sc_hd__mux2_1
X_15757_ _15768_/A vssd1 vssd1 vccd1 vccd1 _15757_/X sky130_fd_sc_hd__buf_1
XFILLER_33_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12969_ _12751_/A _12966_/X _10985_/A _18971_/X vssd1 vssd1 vccd1 vccd1 _12969_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_205_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11571__A _13171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14708_ _20158_/Q _14704_/X _12853_/A _14706_/X vssd1 vssd1 vccd1 vccd1 _20158_/D
+ sky130_fd_sc_hd__a22o_1
X_18476_ _18475_/X _13954_/Y _18903_/S vssd1 vssd1 vccd1 vccd1 _18476_/X sky130_fd_sc_hd__mux2_1
XFILLER_205_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15688_ _15696_/A vssd1 vssd1 vccd1 vccd1 _15688_/X sky130_fd_sc_hd__buf_1
XFILLER_33_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17427_ _19601_/Q _17631_/B vssd1 vssd1 vccd1 vccd1 _17427_/Y sky130_fd_sc_hd__nor2_1
X_14639_ _14639_/A vssd1 vssd1 vccd1 vccd1 _14639_/X sky130_fd_sc_hd__buf_2
XFILLER_159_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17358_ _19488_/Q vssd1 vssd1 vccd1 vccd1 _17358_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16309_ _19383_/Q _16305_/X _16293_/X _16306_/X vssd1 vssd1 vccd1 vccd1 _19383_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_173_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17289_ _21081_/Q vssd1 vssd1 vccd1 vccd1 _17289_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20139__RESET_B repeater250/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19148__S0 _19285_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19028_ _16877_/Y _20841_/Q _19058_/S vssd1 vssd1 vccd1 vccd1 _19948_/D sky130_fd_sc_hd__mux2_1
XFILLER_118_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09961__B1 _09698_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09614_ _20882_/Q _20881_/Q _20884_/Q _20883_/Q vssd1 vssd1 vccd1 vccd1 _09615_/D
+ sky130_fd_sc_hd__or4_4
XFILLER_44_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13273__B1 _13272_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_212_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20909__RESET_B repeater218/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20705_ _21349_/CLK _20705_/D repeater210/X vssd1 vssd1 vccd1 vccd1 _20705_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_197_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13025__B1 _12857_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20636_ _21486_/CLK _20636_/D repeater198/X vssd1 vssd1 vccd1 vccd1 _20636_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20562__RESET_B repeater264/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20567_ _20590_/CLK _20567_/D repeater260/X vssd1 vssd1 vccd1 vccd1 _20567_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__19139__S0 _19285_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13201__A _13217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10320_ _20709_/Q vssd1 vssd1 vccd1 vccd1 _10320_/Y sky130_fd_sc_hd__inv_2
XFILLER_118_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20498_ _20929_/CLK _20498_/D repeater265/X vssd1 vssd1 vccd1 vccd1 _20498_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_3_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10251_ _21352_/Q vssd1 vssd1 vccd1 vccd1 _10268_/A sky130_fd_sc_hd__inv_2
XANTENNA__18203__S _18644_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10182_ _10182_/A vssd1 vssd1 vccd1 vccd1 _10182_/Y sky130_fd_sc_hd__inv_2
XFILLER_120_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21119_ _21120_/CLK _21119_/D repeater231/X vssd1 vssd1 vccd1 vccd1 _21119_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12839__B1 _09626_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14990_ _14961_/D _14870_/B _14987_/Y _14989_/X vssd1 vssd1 vccd1 vccd1 _20092_/D
+ sky130_fd_sc_hd__a211oi_2
X_13941_ _20637_/Q _13865_/A _13939_/Y _20297_/Q _13940_/X vssd1 vssd1 vccd1 vccd1
+ _13947_/C sky130_fd_sc_hd__o221a_1
XFILLER_47_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__21350__RESET_B repeater252/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_219_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19034__S _19046_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_234_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16660_ _19864_/Q _15298_/B _15299_/B vssd1 vssd1 vccd1 vccd1 _16660_/X sky130_fd_sc_hd__a21bo_1
XFILLER_35_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13872_ _20299_/Q vssd1 vssd1 vccd1 vccd1 _14015_/A sky130_fd_sc_hd__inv_2
XFILLER_47_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16450__B1 _19308_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_216_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15611_ _15618_/A vssd1 vssd1 vccd1 vccd1 _15611_/X sky130_fd_sc_hd__buf_1
X_12823_ _12850_/A vssd1 vssd1 vccd1 vccd1 _12842_/A sky130_fd_sc_hd__clkbuf_2
X_16591_ _16688_/A _16590_/X _11407_/Y _16575_/Y _16513_/Y vssd1 vssd1 vccd1 vccd1
+ _19915_/D sky130_fd_sc_hd__o221ai_1
XFILLER_61_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18873__S _18901_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18330_ _18329_/X _14392_/Y _18669_/S vssd1 vssd1 vccd1 vccd1 _18330_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10617__A2 _10614_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15542_ _15673_/A _15542_/B _15778_/C vssd1 vssd1 vccd1 vccd1 _15553_/A sky130_fd_sc_hd__or3_4
XPHY_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12754_ _13048_/A _17201_/A vssd1 vssd1 vccd1 vccd1 _12887_/A sky130_fd_sc_hd__or2_1
XFILLER_131_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_230_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11705_ _11705_/A vssd1 vssd1 vccd1 vccd1 _11705_/X sky130_fd_sc_hd__buf_1
XPHY_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18261_ _18260_/X _12252_/Y _18910_/S vssd1 vssd1 vccd1 vccd1 _18261_/X sky130_fd_sc_hd__mux2_1
XPHY_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13016__B1 _12930_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12685_ _12685_/A vssd1 vssd1 vccd1 vccd1 _12707_/A sky130_fd_sc_hd__buf_2
X_15473_ _15762_/A vssd1 vssd1 vccd1 vccd1 _15473_/X sky130_fd_sc_hd__buf_1
XPHY_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17212_ _17212_/A vssd1 vssd1 vccd1 vccd1 _17573_/A sky130_fd_sc_hd__buf_1
X_14424_ _21469_/Q vssd1 vssd1 vccd1 vccd1 _14424_/Y sky130_fd_sc_hd__inv_2
X_11636_ _11636_/A _20015_/Q vssd1 vssd1 vccd1 vccd1 _11637_/A sky130_fd_sc_hd__or2_1
XFILLER_129_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18192_ _18848_/A0 _10295_/Y _18884_/S vssd1 vssd1 vccd1 vccd1 _18192_/X sky130_fd_sc_hd__mux2_1
XPHY_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17143_ _17143_/A _17162_/B vssd1 vssd1 vccd1 vccd1 _17143_/X sky130_fd_sc_hd__or2_1
XFILLER_155_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14355_ _20209_/Q vssd1 vssd1 vccd1 vccd1 _14496_/A sky130_fd_sc_hd__inv_2
X_11567_ _21130_/Q _11562_/X _11565_/X _11566_/X vssd1 vssd1 vccd1 vccd1 _21130_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20232__RESET_B repeater203/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10518_ _20697_/Q vssd1 vssd1 vccd1 vccd1 _10518_/Y sky130_fd_sc_hd__inv_2
X_13306_ _20542_/Q _13300_/X _13148_/X _13302_/X vssd1 vssd1 vccd1 vccd1 _20542_/D
+ sky130_fd_sc_hd__a22o_1
X_17074_ _19883_/Q _19884_/Q _19885_/Q vssd1 vssd1 vccd1 vccd1 _19883_/D sky130_fd_sc_hd__o21ba_1
X_14286_ _20125_/Q vssd1 vssd1 vccd1 vccd1 _15357_/B sky130_fd_sc_hd__inv_2
XFILLER_128_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11498_ _11498_/A vssd1 vssd1 vccd1 vccd1 _19111_/S sky130_fd_sc_hd__buf_1
XFILLER_170_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13237_ _20574_/Q _13233_/X _13030_/X _13234_/X vssd1 vssd1 vccd1 vccd1 _20574_/D
+ sky130_fd_sc_hd__a22o_1
X_16025_ _19524_/Q _16021_/X _15762_/X _16023_/X vssd1 vssd1 vccd1 vccd1 _19524_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_226_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10449_ _21290_/Q vssd1 vssd1 vccd1 vccd1 _10766_/A sky130_fd_sc_hd__inv_2
XANTENNA__12950__A _14258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13168_ _20602_/Q _13165_/X _13166_/X _13167_/X vssd1 vssd1 vccd1 vccd1 _20602_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11750__B1 _19308_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12119_ _12327_/A vssd1 vssd1 vccd1 vccd1 _12119_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__17481__A2 _17324_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17976_ _17976_/A _17978_/B vssd1 vssd1 vccd1 vccd1 _17976_/Y sky130_fd_sc_hd__nor2_1
XFILLER_69_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13099_ _13099_/A vssd1 vssd1 vccd1 vccd1 _13099_/X sky130_fd_sc_hd__buf_1
XFILLER_242_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19715_ _21009_/CLK _19715_/D vssd1 vssd1 vccd1 vccd1 _19715_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_81_HCLK clkbuf_4_13_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _21480_/CLK sky130_fd_sc_hd__clkbuf_16
X_16927_ _16927_/A _16927_/B vssd1 vssd1 vccd1 vccd1 _16927_/Y sky130_fd_sc_hd__nor2_1
XFILLER_84_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17233__A2 _18019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19646_ _19821_/CLK _19646_/D vssd1 vssd1 vccd1 vccd1 _19646_/Q sky130_fd_sc_hd__dfxtp_1
X_16858_ _16858_/A _16858_/B vssd1 vssd1 vccd1 vccd1 _16858_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__21020__RESET_B repeater238/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_214_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18068__B _18068_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15809_ _19625_/Q _15807_/X _09832_/X _15808_/X vssd1 vssd1 vccd1 vccd1 _19625_/D
+ sky130_fd_sc_hd__a22o_1
X_19577_ _20890_/CLK _19577_/D vssd1 vssd1 vccd1 vccd1 _19577_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__18783__S _18908_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16789_ _19928_/Q vssd1 vssd1 vccd1 vccd1 _16791_/A sky130_fd_sc_hd__inv_2
XFILLER_179_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10608__A2 _20744_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18528_ _17941_/Y _21480_/Q _18669_/S vssd1 vssd1 vccd1 vccd1 _18528_/X sky130_fd_sc_hd__mux2_1
XFILLER_206_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_222_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18459_ _18458_/X _14415_/Y _18897_/S vssd1 vssd1 vccd1 vccd1 _18459_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21470_ _21477_/CLK _21470_/D repeater204/X vssd1 vssd1 vccd1 vccd1 _21470_/Q sky130_fd_sc_hd__dfrtp_1
X_20421_ _20422_/CLK _20421_/D repeater271/X vssd1 vssd1 vccd1 vccd1 _20421_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_119_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13021__A _13041_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20352_ _20982_/CLK _20352_/D repeater279/X vssd1 vssd1 vccd1 vccd1 _20352_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12860__A _12860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20283_ _20661_/CLK _20283_/D repeater262/X vssd1 vssd1 vccd1 vccd1 _20283_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__16332__A _16332_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21179__RESET_B repeater216/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18958__S _18962_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20004__D _20004_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13246__B1 _13245_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18693__S _18849_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12100__A _20395_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12470_ _12470_/A _12488_/A vssd1 vssd1 vccd1 vccd1 _12486_/A sky130_fd_sc_hd__or2_1
XFILLER_184_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12754__B _17201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11421_ _11421_/A vssd1 vssd1 vccd1 vccd1 _11421_/X sky130_fd_sc_hd__buf_1
XFILLER_200_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20619_ _20622_/CLK _20619_/D repeater195/X vssd1 vssd1 vccd1 vccd1 _20619_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_137_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14140_ _14139_/Y _20274_/Q _20545_/Q _14084_/A vssd1 vssd1 vccd1 vccd1 _14140_/X
+ sky130_fd_sc_hd__o22a_1
X_11352_ _21173_/Q vssd1 vssd1 vccd1 vccd1 _11390_/B sky130_fd_sc_hd__inv_2
XFILLER_165_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10303_ _20708_/Q vssd1 vssd1 vccd1 vccd1 _10303_/Y sky130_fd_sc_hd__inv_2
XFILLER_180_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19029__S _19046_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14071_ _14071_/A _14228_/A vssd1 vssd1 vccd1 vccd1 _14072_/B sky130_fd_sc_hd__or2_2
X_11283_ _20914_/Q _20913_/Q _11283_/C _12505_/B vssd1 vssd1 vccd1 vccd1 _11299_/D
+ sky130_fd_sc_hd__or4_4
X_13022_ _20681_/Q _13019_/X _12849_/X _13021_/X vssd1 vssd1 vccd1 vccd1 _20681_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_140_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input51_A HWDATA[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10234_ _21369_/Q vssd1 vssd1 vccd1 vccd1 _10284_/A sky130_fd_sc_hd__inv_2
XFILLER_180_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18868__S _18928_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17830_ _17830_/A vssd1 vssd1 vccd1 vccd1 _17830_/X sky130_fd_sc_hd__buf_2
X_10165_ _10183_/A vssd1 vssd1 vccd1 vccd1 _10166_/A sky130_fd_sc_hd__buf_1
XFILLER_120_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_158_HCLK_A clkbuf_opt_1_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17761_ _19629_/Q vssd1 vssd1 vccd1 vccd1 _17761_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14973_ _15059_/B vssd1 vssd1 vccd1 vccd1 _14973_/X sky130_fd_sc_hd__buf_1
X_10096_ _10153_/A _20789_/Q _21392_/Q _10095_/Y vssd1 vssd1 vccd1 vccd1 _10096_/X
+ sky130_fd_sc_hd__o22a_1
X_19500_ _20327_/CLK _19500_/D vssd1 vssd1 vccd1 vccd1 _19500_/Q sky130_fd_sc_hd__dfxtp_1
X_16712_ _16718_/A _18937_/X vssd1 vssd1 vccd1 vccd1 _19899_/D sky130_fd_sc_hd__and2_1
XANTENNA__18412__A1 _13911_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13924_ _13923_/Y _20309_/Q _20652_/Q _13972_/B vssd1 vssd1 vccd1 vccd1 _13930_/B
+ sky130_fd_sc_hd__o22a_1
X_17692_ _19596_/Q vssd1 vssd1 vccd1 vccd1 _17692_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19431_ _20137_/CLK _19431_/D vssd1 vssd1 vccd1 vccd1 _19431_/Q sky130_fd_sc_hd__dfxtp_1
X_16643_ _16643_/A _18958_/X vssd1 vssd1 vccd1 vccd1 _19856_/D sky130_fd_sc_hd__and2_1
XFILLER_47_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13237__B1 _13030_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13855_ _20306_/Q vssd1 vssd1 vccd1 vccd1 _13882_/A sky130_fd_sc_hd__inv_2
XANTENNA_repeater190_A repeater233/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12806_ _20775_/Q _12803_/X _11739_/X _12804_/X vssd1 vssd1 vccd1 vccd1 _20775_/D
+ sky130_fd_sc_hd__a22o_1
X_19362_ _21001_/CLK _19362_/D vssd1 vssd1 vccd1 vccd1 _19362_/Q sky130_fd_sc_hd__dfxtp_1
X_16574_ _16576_/B _16573_/A _16507_/B _16573_/Y _11371_/A vssd1 vssd1 vccd1 vccd1
+ _16574_/X sky130_fd_sc_hd__o221a_1
XANTENNA__18176__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13786_ _13767_/X _13786_/B _13786_/C _13786_/D vssd1 vssd1 vccd1 vccd1 _13837_/B
+ sky130_fd_sc_hd__and4b_1
X_10998_ _21012_/Q vssd1 vssd1 vccd1 vccd1 _11008_/B sky130_fd_sc_hd__inv_2
XFILLER_222_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18313_ _18312_/X _10618_/Y _18897_/S vssd1 vssd1 vccd1 vccd1 _18313_/X sky130_fd_sc_hd__mux2_1
X_15525_ _19759_/Q _15516_/X _15524_/X _15519_/X vssd1 vssd1 vccd1 vccd1 _19759_/D
+ sky130_fd_sc_hd__a22o_1
X_19293_ _19776_/CLK _19293_/D vssd1 vssd1 vccd1 vccd1 _19293_/Q sky130_fd_sc_hd__dfxtp_1
X_12737_ _12750_/A _14686_/B vssd1 vssd1 vccd1 vccd1 _14685_/A sky130_fd_sc_hd__or2_1
XFILLER_188_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20413__RESET_B repeater185/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17923__B1 _18928_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14737__B1 _13712_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18244_ _19136_/X _20162_/Q _18249_/S vssd1 vssd1 vccd1 vccd1 _18244_/X sky130_fd_sc_hd__mux2_1
XFILLER_230_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15456_ _15663_/A vssd1 vssd1 vccd1 vccd1 _15456_/X sky130_fd_sc_hd__clkbuf_2
XPHY_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12668_ input55/X vssd1 vssd1 vccd1 vccd1 _12668_/X sky130_fd_sc_hd__clkbuf_4
XPHY_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14407_ _20233_/Q _20025_/Q _20233_/Q _20025_/Q vssd1 vssd1 vccd1 vccd1 _14407_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_11619_ _21110_/Q _11613_/A _11614_/Y _11617_/X _11618_/Y vssd1 vssd1 vccd1 vccd1
+ _21110_/D sky130_fd_sc_hd__a32o_1
X_18175_ _18174_/X _17014_/Y _18875_/S vssd1 vssd1 vccd1 vccd1 _18175_/X sky130_fd_sc_hd__mux2_1
X_15387_ _19819_/Q _15376_/X _15386_/X _15380_/X vssd1 vssd1 vccd1 vccd1 _19819_/D
+ sky130_fd_sc_hd__a22o_1
X_12599_ _20873_/Q _12594_/X _18225_/X _12595_/X vssd1 vssd1 vccd1 vccd1 _20873_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17126_ _19325_/Q vssd1 vssd1 vccd1 vccd1 _17126_/Y sky130_fd_sc_hd__inv_2
X_14338_ _20227_/Q vssd1 vssd1 vccd1 vccd1 _14461_/A sky130_fd_sc_hd__inv_2
XFILLER_183_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17057_ _20036_/Q vssd1 vssd1 vccd1 vccd1 _17057_/Y sky130_fd_sc_hd__inv_2
X_14269_ _20247_/Q _14267_/X _13707_/X _14268_/X vssd1 vssd1 vccd1 vccd1 _20247_/D
+ sky130_fd_sc_hd__a22o_1
X_16008_ _16008_/A vssd1 vssd1 vccd1 vccd1 _16008_/X sky130_fd_sc_hd__buf_1
XANTENNA__18778__S _18897_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21272__RESET_B repeater245/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16662__B1 _18962_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17959_ _20415_/Q vssd1 vssd1 vccd1 vccd1 _17959_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_17_HCLK_A clkbuf_4_3_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20970_ _20971_/CLK _20970_/D repeater187/X vssd1 vssd1 vccd1 vccd1 _20970_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_226_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19629_ _21040_/CLK _19629_/D vssd1 vssd1 vccd1 vccd1 _19629_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_5_HCLK_A clkbuf_opt_2_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12855__A _12855_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14728__B1 _13714_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_opt_6_HCLK clkbuf_opt_7_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_opt_6_HCLK/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_31_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21453_ _21453_/CLK _21453_/D repeater247/X vssd1 vssd1 vccd1 vccd1 _21453_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__13400__B1 _13277_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20404_ _20422_/CLK _20404_/D repeater188/X vssd1 vssd1 vccd1 vccd1 _20404_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_174_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21384_ _21390_/CLK _21384_/D repeater252/X vssd1 vssd1 vccd1 vccd1 _21384_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_134_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20335_ _20809_/CLK _20335_/D repeater188/X vssd1 vssd1 vccd1 vccd1 _20335_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_190_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20539__CLK _20592_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_227_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20266_ _20286_/CLK _20266_/D repeater264/X vssd1 vssd1 vccd1 vccd1 _20266_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18688__S _18880_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20197_ _20626_/CLK _20197_/D repeater193/X vssd1 vssd1 vccd1 vccd1 _20197_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_163_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11970_ _11973_/A _11966_/X _13717_/B _18974_/X vssd1 vssd1 vccd1 vccd1 _11978_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_72_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20924__RESET_B repeater267/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10921_ _21206_/Q _11810_/A _10920_/Y _21033_/Q vssd1 vssd1 vccd1 vccd1 _10931_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_84_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10852_ _18279_/X _10847_/X _21273_/Q _10849_/X vssd1 vssd1 vccd1 vccd1 _21273_/D
+ sky130_fd_sc_hd__o22a_1
X_13640_ _13652_/A vssd1 vssd1 vccd1 vccd1 _13640_/X sky130_fd_sc_hd__buf_1
XFILLER_72_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10783_ _10783_/A _10783_/B vssd1 vssd1 vccd1 vccd1 _10784_/A sky130_fd_sc_hd__or2_1
XFILLER_12_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13571_ _20413_/Q _13566_/X _13489_/X _13567_/X vssd1 vssd1 vccd1 vccd1 _20413_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16237__A _16237_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15310_ _15310_/A vssd1 vssd1 vccd1 vccd1 _16632_/A sky130_fd_sc_hd__inv_2
XFILLER_200_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12522_ _20915_/Q _12520_/X _12502_/A _12521_/X vssd1 vssd1 vccd1 vccd1 _20915_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_200_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14719__B1 _14258_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16290_ _19393_/Q _16287_/X _16288_/X _16289_/X vssd1 vssd1 vccd1 vccd1 _19393_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15241_ _20495_/Q _15088_/A _15237_/Y _20046_/Q _15240_/X vssd1 vssd1 vccd1 vccd1
+ _15250_/B sky130_fd_sc_hd__o221a_1
X_12453_ _12453_/A vssd1 vssd1 vccd1 vccd1 _12453_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_184_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11404_ _11420_/A vssd1 vssd1 vccd1 vccd1 _11404_/X sky130_fd_sc_hd__buf_1
X_15172_ _15084_/A _15084_/B _15179_/A _15169_/Y vssd1 vssd1 vccd1 vccd1 _20070_/D
+ sky130_fd_sc_hd__a211oi_2
X_12384_ _20955_/Q _12383_/Y _12373_/X _12310_/B vssd1 vssd1 vccd1 vccd1 _20955_/D
+ sky130_fd_sc_hd__o211a_1
X_11335_ _11363_/A _21178_/Q _11362_/C vssd1 vssd1 vccd1 vccd1 _11346_/C sky130_fd_sc_hd__or3_1
X_14123_ _20543_/Q _20272_/Q _14122_/Y _14082_/A vssd1 vssd1 vccd1 vccd1 _14123_/X
+ sky130_fd_sc_hd__o22a_1
X_19980_ _20428_/CLK _19980_/D repeater270/X vssd1 vssd1 vccd1 vccd1 _19980_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_126_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18931_ _16739_/X _21193_/Q _18931_/S vssd1 vssd1 vccd1 vccd1 _18931_/X sky130_fd_sc_hd__mux2_1
XFILLER_153_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11266_ _20908_/Q _20907_/Q _20906_/Q _20905_/Q vssd1 vssd1 vccd1 vccd1 _11294_/A
+ sky130_fd_sc_hd__or4_4
X_14054_ _20274_/Q vssd1 vssd1 vccd1 vccd1 _14084_/A sky130_fd_sc_hd__inv_2
XANTENNA__18598__S _18644_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13005_ _13012_/A vssd1 vssd1 vccd1 vccd1 _13005_/X sky130_fd_sc_hd__buf_1
XFILLER_79_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10217_ _21381_/Q _10216_/Y _10203_/B _10140_/X vssd1 vssd1 vccd1 vccd1 _21381_/D
+ sky130_fd_sc_hd__o211a_1
X_18862_ _18861_/X _17275_/Y _18927_/S vssd1 vssd1 vccd1 vccd1 _18862_/X sky130_fd_sc_hd__mux2_1
XANTENNA__18094__C1 _18093_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater203_A repeater204/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11197_ _21214_/Q _11191_/X _10898_/X _11193_/X vssd1 vssd1 vccd1 vccd1 _21214_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_121_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17813_ _20819_/Q _18666_/S vssd1 vssd1 vccd1 vccd1 _17813_/Y sky130_fd_sc_hd__nand2_1
XFILLER_39_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10148_ _10220_/A _10148_/B vssd1 vssd1 vccd1 vccd1 _10149_/B sky130_fd_sc_hd__or2_2
X_18793_ _18792_/X _09752_/Y _18928_/S vssd1 vssd1 vccd1 vccd1 _18793_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17744_ _19397_/Q vssd1 vssd1 vccd1 vccd1 _17744_/Y sky130_fd_sc_hd__inv_2
X_14956_ _14883_/A _14883_/B _14884_/Y _15025_/C vssd1 vssd1 vccd1 vccd1 _20106_/D
+ sky130_fd_sc_hd__a211oi_2
X_10079_ _21407_/Q vssd1 vssd1 vccd1 vccd1 _10079_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13907_ _20634_/Q vssd1 vssd1 vccd1 vccd1 _13907_/Y sky130_fd_sc_hd__inv_2
XFILLER_223_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17675_ _19388_/Q vssd1 vssd1 vccd1 vccd1 _17675_/Y sky130_fd_sc_hd__inv_2
X_14887_ _20584_/Q _20095_/Q _14886_/Y _14961_/C vssd1 vssd1 vccd1 vccd1 _14901_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_236_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19414_ _19784_/CLK _19414_/D vssd1 vssd1 vccd1 vccd1 _19414_/Q sky130_fd_sc_hd__dfxtp_1
X_16626_ _21070_/Q vssd1 vssd1 vccd1 vccd1 _16628_/A sky130_fd_sc_hd__inv_2
X_13838_ _14597_/A vssd1 vssd1 vccd1 vccd1 _14639_/A sky130_fd_sc_hd__buf_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19345_ _19626_/CLK _19345_/D vssd1 vssd1 vccd1 vccd1 _19345_/Q sky130_fd_sc_hd__dfxtp_1
X_16557_ _16566_/A _21148_/Q _16554_/Y _16556_/Y vssd1 vssd1 vccd1 vccd1 _16557_/X
+ sky130_fd_sc_hd__a31o_1
X_13769_ _20206_/Q vssd1 vssd1 vccd1 vccd1 _14595_/A sky130_fd_sc_hd__inv_2
XANTENNA__13630__B1 _13489_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15508_ _15516_/A vssd1 vssd1 vccd1 vccd1 _15519_/A sky130_fd_sc_hd__inv_2
XFILLER_149_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19276_ _19272_/X _19273_/X _19274_/X _19275_/X _21005_/Q _21006_/Q vssd1 vssd1 vccd1
+ vccd1 _19276_/X sky130_fd_sc_hd__mux4_2
XFILLER_31_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19704__CLK _19706_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16488_ _16488_/A vssd1 vssd1 vccd1 vccd1 _18928_/S sky130_fd_sc_hd__clkinv_16
XFILLER_248_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18227_ _20851_/Q input31/X _18236_/S vssd1 vssd1 vccd1 vccd1 _18227_/X sky130_fd_sc_hd__mux2_1
XFILLER_248_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15439_ _19795_/Q _15434_/X _15386_/X _15436_/X vssd1 vssd1 vccd1 vccd1 _19795_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_163_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18158_ _18157_/X _21299_/Q _18617_/S vssd1 vssd1 vccd1 vccd1 _18158_/X sky130_fd_sc_hd__mux2_1
XANTENNA__21453__RESET_B repeater247/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18081__B _18083_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17109_ _21213_/Q vssd1 vssd1 vccd1 vccd1 _18109_/A sky130_fd_sc_hd__inv_2
XFILLER_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18089_ _18619_/X _17954_/A _18658_/X _17572_/B vssd1 vssd1 vccd1 vccd1 _18090_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_172_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20120_ _20172_/CLK _20120_/D repeater248/X vssd1 vssd1 vccd1 vccd1 _20120_/Q sky130_fd_sc_hd__dfrtp_1
X_09931_ _16342_/A vssd1 vssd1 vccd1 vccd1 _09931_/X sky130_fd_sc_hd__buf_1
XFILLER_132_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13697__B1 _13584_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20051_ _20066_/CLK _20051_/D repeater281/X vssd1 vssd1 vccd1 vccd1 _20051_/Q sky130_fd_sc_hd__dfrtp_4
X_09862_ _09853_/X _09857_/A _15314_/A vssd1 vssd1 vccd1 vccd1 _09862_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__18301__S _18666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09793_ _09804_/A _09803_/A _09793_/C _21457_/Q vssd1 vssd1 vccd1 vccd1 _16620_/C
+ sky130_fd_sc_hd__or4_4
XFILLER_133_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_141_HCLK_A clkbuf_4_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater153 _18898_/S vssd1 vssd1 vccd1 vccd1 _18748_/S sky130_fd_sc_hd__buf_8
XFILLER_39_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrepeater164 _18835_/S vssd1 vssd1 vccd1 vccd1 _18787_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_27_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater175 _18644_/S vssd1 vssd1 vccd1 vccd1 _18885_/S sky130_fd_sc_hd__buf_8
XPHY_4307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater186 repeater187/X vssd1 vssd1 vccd1 vccd1 repeater186/X sky130_fd_sc_hd__buf_8
XFILLER_66_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20953_ _20957_/CLK _20953_/D repeater187/X vssd1 vssd1 vccd1 vccd1 _20953_/Q sky130_fd_sc_hd__dfrtp_4
Xrepeater197 repeater198/X vssd1 vssd1 vccd1 vccd1 repeater197/X sky130_fd_sc_hd__clkbuf_8
XPHY_4329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20884_ _21444_/CLK _20884_/D repeater243/X vssd1 vssd1 vccd1 vccd1 _20884_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_3639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13621__B1 _13560_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18560__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21436_ _21438_/CLK _21436_/D repeater239/X vssd1 vssd1 vccd1 vccd1 _21436_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__13924__A1 _13923_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18312__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21194__RESET_B repeater220/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21367_ _21367_/CLK _21367_/D repeater254/X vssd1 vssd1 vccd1 vccd1 _21367_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21123__RESET_B repeater190/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11120_ _21225_/Q _09744_/X _11112_/X _11113_/X vssd1 vssd1 vccd1 vccd1 _11120_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_107_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20318_ _20322_/CLK _20318_/D repeater262/X vssd1 vssd1 vccd1 vccd1 _20318_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_122_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21298_ _21302_/CLK _21298_/D repeater209/X vssd1 vssd1 vccd1 vccd1 _21298_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_107_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11051_ _11100_/A vssd1 vssd1 vccd1 vccd1 _11051_/X sky130_fd_sc_hd__buf_1
XFILLER_1_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20249_ _21421_/CLK _20249_/D repeater214/X vssd1 vssd1 vccd1 vccd1 _20249_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18211__S _18896_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10002_ _09999_/X _10000_/X _20018_/Q _10001_/Y vssd1 vssd1 vccd1 vccd1 _17034_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_77_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11664__A _21071_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14810_ _14800_/A _14800_/B _14800_/Y _14807_/X vssd1 vssd1 vccd1 vccd1 _14810_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_190_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18379__A0 _17281_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15790_ _19633_/Q _15787_/X _15788_/X _15789_/X vssd1 vssd1 vccd1 vccd1 _19633_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14040__A _20288_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_134_HCLK clkbuf_4_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _21372_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_123_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input14_A HADDR[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14741_ _19122_/X vssd1 vssd1 vccd1 vccd1 _14744_/A sky130_fd_sc_hd__inv_2
XFILLER_217_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11953_ _21006_/Q _11955_/A _11124_/Y _11952_/A vssd1 vssd1 vccd1 vccd1 _21006_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_233_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_63_HCLK_A clkbuf_4_14_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20076__RESET_B repeater259/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19042__S _19046_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_232_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17460_ _17455_/Y _17301_/A _17456_/Y _17378_/X _17459_/X vssd1 vssd1 vccd1 vccd1
+ _17460_/X sky130_fd_sc_hd__o221a_1
X_10904_ _17019_/A _11584_/C vssd1 vssd1 vccd1 vccd1 _11021_/B sky130_fd_sc_hd__and2_1
XFILLER_233_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14672_ _12740_/B _12735_/A _14674_/A _11800_/A vssd1 vssd1 vccd1 vccd1 _14673_/A
+ sky130_fd_sc_hd__o211a_1
X_11884_ _11874_/Y _10983_/A _21022_/Q _11883_/X vssd1 vssd1 vccd1 vccd1 _11885_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_45_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20005__RESET_B repeater190/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16411_ _19330_/Q _16406_/X _16202_/X _16408_/X vssd1 vssd1 vccd1 vccd1 _19330_/D
+ sky130_fd_sc_hd__a22o_1
X_13623_ _20385_/Q _13619_/X _13477_/X _13620_/X vssd1 vssd1 vccd1 vccd1 _20385_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_60_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17391_ _17388_/Y _14256_/A _17389_/Y _17390_/X vssd1 vssd1 vccd1 vccd1 _17391_/X
+ sky130_fd_sc_hd__o22a_1
X_10835_ _10758_/A _10758_/B _10827_/X _10833_/Y vssd1 vssd1 vccd1 vccd1 _21281_/D
+ sky130_fd_sc_hd__a211oi_4
XFILLER_44_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13612__B1 _13547_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18881__S _18899_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19130_ _19654_/Q _19646_/Q _19630_/Q _19814_/Q _19285_/S0 _21017_/Q vssd1 vssd1
+ vccd1 vccd1 _19130_/X sky130_fd_sc_hd__mux4_2
X_16342_ _16342_/A vssd1 vssd1 vccd1 vccd1 _16342_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_186_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13554_ _20423_/Q _13549_/X _13553_/X _13551_/X vssd1 vssd1 vccd1 vccd1 _20423_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_13_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10766_ _10766_/A _10818_/A vssd1 vssd1 vccd1 vccd1 _10767_/B sky130_fd_sc_hd__or2_1
XFILLER_158_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12505_ _12505_/A _12505_/B vssd1 vssd1 vccd1 vccd1 _12506_/B sky130_fd_sc_hd__or2_1
X_19061_ _21190_/Q _21132_/Q _19910_/Q vssd1 vssd1 vccd1 vccd1 _19061_/X sky130_fd_sc_hd__mux2_1
XFILLER_201_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15365__B1 _15343_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16273_ _19399_/Q _16269_/X _16125_/X _16270_/X vssd1 vssd1 vccd1 vccd1 _19399_/D
+ sky130_fd_sc_hd__a22o_1
X_10697_ _10697_/A vssd1 vssd1 vccd1 vccd1 _10697_/Y sky130_fd_sc_hd__inv_2
XANTENNA_repeater153_A _18898_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13485_ input47/X vssd1 vssd1 vccd1 vccd1 _13485_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_173_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18012_ _18374_/X _17951_/X _18153_/X _17952_/X vssd1 vssd1 vccd1 vccd1 _18014_/C
+ sky130_fd_sc_hd__a22o_1
X_15224_ _20468_/Q _15062_/A _15221_/Y _20051_/Q _15223_/X vssd1 vssd1 vccd1 vccd1
+ _15232_/B sky130_fd_sc_hd__o221a_1
X_12436_ _12436_/A _12436_/B vssd1 vssd1 vccd1 vccd1 _12437_/C sky130_fd_sc_hd__nor2_1
XANTENNA__18303__A0 _17079_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15155_ _20464_/Q _15090_/Y _20457_/Q _15104_/X vssd1 vssd1 vccd1 vccd1 _15155_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_5_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12367_ _20965_/Q _12366_/Y _12359_/X _12319_/B vssd1 vssd1 vccd1 vccd1 _20965_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_154_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output82_A _17883_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14106_ _17809_/A _20267_/Q _17940_/A _20276_/Q vssd1 vssd1 vccd1 vccd1 _14106_/X
+ sky130_fd_sc_hd__o22a_1
X_11318_ _16689_/A _12525_/C vssd1 vssd1 vccd1 vccd1 _11322_/B sky130_fd_sc_hd__nand2_1
XFILLER_181_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19963_ _20890_/CLK _19963_/D repeater185/X vssd1 vssd1 vccd1 vccd1 _19963_/Q sky130_fd_sc_hd__dfrtp_1
X_15086_ _15086_/A _15086_/B vssd1 vssd1 vccd1 vccd1 _15165_/A sky130_fd_sc_hd__or2_1
X_12298_ _20949_/Q vssd1 vssd1 vccd1 vccd1 _12298_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11249_ _19062_/X _11244_/X _21190_/Q _11245_/X vssd1 vssd1 vccd1 vccd1 _21190_/D
+ sky130_fd_sc_hd__a22o_1
X_14037_ _14037_/A _14037_/B _14037_/C vssd1 vssd1 vccd1 vccd1 _20292_/D sky130_fd_sc_hd__nor3_1
X_18914_ _18913_/X _21412_/Q _20870_/Q vssd1 vssd1 vccd1 vccd1 _18914_/X sky130_fd_sc_hd__mux2_1
X_19894_ _21191_/CLK _19894_/D repeater222/X vssd1 vssd1 vccd1 vccd1 _19894_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__20846__RESET_B repeater243/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18845_ _18845_/A0 _13830_/Y _18896_/S vssd1 vssd1 vccd1 vccd1 _18845_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18776_ _18775_/X _10757_/A _18880_/S vssd1 vssd1 vccd1 vccd1 _18776_/X sky130_fd_sc_hd__mux2_1
X_15988_ _15994_/A vssd1 vssd1 vccd1 vccd1 _15988_/X sky130_fd_sc_hd__buf_1
X_17727_ _17724_/Y _17290_/X _16631_/A _17292_/X _17726_/X vssd1 vssd1 vccd1 vccd1
+ _17727_/X sky130_fd_sc_hd__o221a_1
X_14939_ _20583_/Q vssd1 vssd1 vccd1 vccd1 _14939_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17658_ _18718_/X _17397_/X _18715_/X _17398_/X _17657_/X vssd1 vssd1 vccd1 vccd1
+ _17658_/X sky130_fd_sc_hd__o221a_1
XANTENNA__18076__B _18076_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16609_ _16609_/A _19913_/Q vssd1 vssd1 vccd1 vccd1 _17064_/B sky130_fd_sc_hd__or2_2
XFILLER_23_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18791__S _18926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17589_ _19643_/Q vssd1 vssd1 vccd1 vccd1 _17589_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19328_ _20137_/CLK _19328_/D vssd1 vssd1 vccd1 vccd1 _19328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_204_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18542__A0 _18541_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19259_ _17265_/Y _17266_/Y _17267_/Y _17268_/Y _20130_/Q _20131_/Q vssd1 vssd1 vccd1
+ vccd1 _19259_/X sky130_fd_sc_hd__mux4_1
XANTENNA__15356__B1 _15355_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19098__A1 _21080_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20040__SET_B repeater216/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_15_HCLK clkbuf_opt_2_HCLK/A vssd1 vssd1 vccd1 vccd1 _19811_/CLK sky130_fd_sc_hd__clkbuf_16
X_21221_ _21222_/CLK _21221_/D repeater235/X vssd1 vssd1 vccd1 vccd1 _21221_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__19193__S1 _20122_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21152_ _21424_/CLK _21152_/D repeater229/X vssd1 vssd1 vccd1 vccd1 _21152_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_132_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20103_ _20107_/CLK _20103_/D repeater259/X vssd1 vssd1 vccd1 vccd1 _20103_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_104_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09914_ _21255_/Q _17022_/A _09905_/X _09910_/X _09913_/X vssd1 vssd1 vccd1 vccd1
+ _09914_/X sky130_fd_sc_hd__o2111a_1
X_21083_ _21424_/CLK _21083_/D repeater230/X vssd1 vssd1 vccd1 vccd1 _21083_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA__16340__A _16340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_157_HCLK clkbuf_opt_1_HCLK/A vssd1 vssd1 vccd1 vccd1 _21453_/CLK sky130_fd_sc_hd__clkbuf_16
X_20034_ _21445_/CLK _20034_/D repeater244/X vssd1 vssd1 vccd1 vccd1 _20034_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_58_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09845_ _21441_/Q vssd1 vssd1 vccd1 vccd1 _09846_/C sky130_fd_sc_hd__inv_2
XANTENNA_input6_A HADDR[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09776_ _09787_/A _09781_/B _21462_/Q _09775_/Y vssd1 vssd1 vccd1 vccd1 _21462_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_160_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20936_ _20937_/CLK _20936_/D repeater277/X vssd1 vssd1 vccd1 vccd1 _20936_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10120__A2 _10119_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_214_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14398__A1 _21485_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20867_ _21444_/CLK _20867_/D repeater247/X vssd1 vssd1 vccd1 vccd1 _20867_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10620_ _10557_/A _20758_/Q _10574_/C _20767_/Q vssd1 vssd1 vccd1 vccd1 _10620_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_168_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21375__RESET_B repeater257/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20798_ _21374_/CLK _20798_/D repeater253/X vssd1 vssd1 vccd1 vccd1 _20798_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10551_ _10707_/A _10706_/A _10551_/C _10708_/A vssd1 vssd1 vccd1 vccd1 _10552_/D
+ sky130_fd_sc_hd__or4_4
XFILLER_10_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18206__S _18784_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19089__A1 _21057_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10482_ _21300_/Q _10480_/Y _10765_/A _20678_/Q vssd1 vssd1 vccd1 vccd1 _10482_/X
+ sky130_fd_sc_hd__o22a_1
X_13270_ input61/X vssd1 vssd1 vccd1 vccd1 _13270_/X sky130_fd_sc_hd__buf_2
XFILLER_211_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19184__S1 _20122_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12221_ _20505_/Q vssd1 vssd1 vccd1 vccd1 _12221_/Y sky130_fd_sc_hd__inv_2
X_21419_ _21419_/CLK _21419_/D repeater232/X vssd1 vssd1 vccd1 vccd1 _21419_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12152_ _12036_/X _20346_/Q _20956_/Q _12150_/Y _12151_/X vssd1 vssd1 vccd1 vccd1
+ _12159_/B sky130_fd_sc_hd__a221o_1
XFILLER_162_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11103_ _11103_/A vssd1 vssd1 vccd1 vccd1 _21230_/D sky130_fd_sc_hd__inv_2
XFILLER_123_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_2_2_0_HCLK_A clkbuf_2_3_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19037__S _19046_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12083_ _20374_/Q vssd1 vssd1 vccd1 vccd1 _12083_/Y sky130_fd_sc_hd__inv_2
X_16960_ _16958_/A _16958_/C _19968_/Q vssd1 vssd1 vccd1 vccd1 _16960_/X sky130_fd_sc_hd__o21a_1
XFILLER_2_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11034_ _19961_/Q _16926_/A vssd1 vssd1 vccd1 vccd1 _16930_/A sky130_fd_sc_hd__or2_2
X_15911_ _15911_/A vssd1 vssd1 vccd1 vccd1 _15911_/X sky130_fd_sc_hd__buf_1
XFILLER_49_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16891_ _19952_/Q vssd1 vssd1 vccd1 vccd1 _16891_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18876__S _18899_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18630_ _18629_/X _12270_/Y _18910_/S vssd1 vssd1 vccd1 vccd1 _18630_/X sky130_fd_sc_hd__mux2_1
XFILLER_209_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15842_ _15842_/A vssd1 vssd1 vccd1 vccd1 _15842_/X sky130_fd_sc_hd__buf_1
XANTENNA__10895__B1 _10894_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18561_ _18560_/X _14396_/Y _18897_/S vssd1 vssd1 vccd1 vccd1 _18561_/X sky130_fd_sc_hd__mux2_1
XANTENNA_output120_A _18113_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15773_ _19640_/Q _15768_/X _15772_/X _15770_/X vssd1 vssd1 vccd1 vccd1 _19640_/D
+ sky130_fd_sc_hd__a22o_1
X_12985_ _13018_/A vssd1 vssd1 vccd1 vccd1 _13020_/A sky130_fd_sc_hd__inv_2
X_17512_ _19345_/Q vssd1 vssd1 vccd1 vccd1 _17512_/Y sky130_fd_sc_hd__inv_2
X_14724_ _14724_/A vssd1 vssd1 vccd1 vccd1 _14724_/X sky130_fd_sc_hd__buf_1
X_18492_ _18491_/X _14930_/Y _18907_/S vssd1 vssd1 vccd1 vccd1 _18492_/X sky130_fd_sc_hd__mux2_1
XFILLER_73_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11936_ _21009_/Q vssd1 vssd1 vccd1 vccd1 _11936_/Y sky130_fd_sc_hd__inv_2
XFILLER_233_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17443_ _19465_/Q vssd1 vssd1 vccd1 vccd1 _17443_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14655_ _20173_/Q vssd1 vssd1 vccd1 vccd1 _14655_/Y sky130_fd_sc_hd__inv_2
XFILLER_233_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11867_ _11867_/A vssd1 vssd1 vccd1 vccd1 _21027_/D sky130_fd_sc_hd__inv_2
XFILLER_14_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13606_ _13631_/A vssd1 vssd1 vccd1 vccd1 _13633_/A sky130_fd_sc_hd__inv_2
X_17374_ _20399_/Q vssd1 vssd1 vccd1 vccd1 _17374_/Y sky130_fd_sc_hd__inv_2
X_10818_ _10818_/A vssd1 vssd1 vccd1 vccd1 _10818_/Y sky130_fd_sc_hd__inv_2
XPHY_3992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14586_ _14586_/A _14616_/A vssd1 vssd1 vccd1 vccd1 _14587_/B sky130_fd_sc_hd__or2_2
XANTENNA__18524__A0 _18523_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_38_HCLK _20004_/CLK vssd1 vssd1 vccd1 vccd1 _21183_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__17327__B2 _17326_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11798_ input70/X _11793_/X _21040_/Q _11797_/X vssd1 vssd1 vccd1 vccd1 _21040_/D
+ sky130_fd_sc_hd__o22a_1
X_19113_ _19844_/Q _16596_/X _19870_/Q vssd1 vssd1 vccd1 vccd1 _19113_/X sky130_fd_sc_hd__mux2_1
XFILLER_186_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16325_ _16325_/A _16325_/B _16325_/C vssd1 vssd1 vccd1 vccd1 _16334_/A sky130_fd_sc_hd__or3_4
XFILLER_9_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13537_ _13566_/A vssd1 vssd1 vccd1 vccd1 _13537_/X sky130_fd_sc_hd__buf_1
XFILLER_9_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10749_ _19947_/Q _19946_/Q _16868_/A vssd1 vssd1 vccd1 vccd1 _16872_/A sky130_fd_sc_hd__or3_4
XFILLER_173_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19044_ _16807_/Y _20825_/Q _19046_/S vssd1 vssd1 vccd1 vccd1 _19932_/D sky130_fd_sc_hd__mux2_1
XFILLER_145_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16256_ _16256_/A vssd1 vssd1 vccd1 vccd1 _16256_/X sky130_fd_sc_hd__buf_1
XFILLER_185_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13468_ _20460_/Q _13466_/X _13277_/X _13467_/X vssd1 vssd1 vccd1 vccd1 _20460_/D
+ sky130_fd_sc_hd__a22o_1
X_15207_ _15065_/A _15065_/B _15205_/Y _15193_/X vssd1 vssd1 vccd1 vccd1 _20050_/D
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__19175__S1 _20122_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12419_ _12419_/A _12419_/B vssd1 vssd1 vccd1 vccd1 _12465_/A sky130_fd_sc_hd__or2_1
X_16187_ _16187_/A vssd1 vssd1 vccd1 vccd1 _16187_/X sky130_fd_sc_hd__buf_1
XFILLER_142_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13399_ _13411_/A vssd1 vssd1 vccd1 vccd1 _13399_/X sky130_fd_sc_hd__buf_1
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15138_ _20444_/Q vssd1 vssd1 vccd1 vccd1 _15138_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15069_ _15069_/A _15198_/A vssd1 vssd1 vccd1 vccd1 _15070_/B sky130_fd_sc_hd__or2_2
X_19946_ _20841_/CLK _19946_/D repeater256/X vssd1 vssd1 vccd1 vccd1 _19946_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__15510__B1 _15450_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_229_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19877_ _21193_/CLK _19877_/D repeater223/X vssd1 vssd1 vccd1 vccd1 _19877_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18786__S _18908_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09630_ input48/X vssd1 vssd1 vccd1 vccd1 _09630_/X sky130_fd_sc_hd__buf_4
X_18828_ _18827_/X _14526_/Y _18929_/S vssd1 vssd1 vccd1 vccd1 _18828_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18759_ _18758_/X _09759_/Y _18928_/S vssd1 vssd1 vccd1 vccd1 _18759_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20721_ _20724_/CLK _20721_/D repeater264/X vssd1 vssd1 vccd1 vccd1 _20721_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_23_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20652_ _20657_/CLK _20652_/D repeater196/X vssd1 vssd1 vccd1 vccd1 _20652_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17318__A1 _18844_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17318__B2 _17862_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20583_ _20946_/CLK _20583_/D repeater258/X vssd1 vssd1 vccd1 vccd1 _20583_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_165_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12863__A _12863_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19863__RESET_B repeater225/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19166__S1 _20124_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_219_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12563__B1 input37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21204_ _21255_/CLK _21204_/D repeater240/X vssd1 vssd1 vccd1 vccd1 _21204_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_145_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21135_ _21334_/CLK _21135_/D repeater221/X vssd1 vssd1 vccd1 vccd1 _21135_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA__15501__B1 _15424_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21066_ _21134_/CLK _21066_/D repeater230/X vssd1 vssd1 vccd1 vccd1 _21066_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18696__S _18906_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20017_ _21417_/CLK _20017_/D repeater230/X vssd1 vssd1 vccd1 vccd1 _20017_/Q sky130_fd_sc_hd__dfrtp_1
X_09828_ _15873_/A vssd1 vssd1 vccd1 vccd1 _09828_/X sky130_fd_sc_hd__buf_1
XFILLER_171_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09759_ _20148_/Q vssd1 vssd1 vccd1 vccd1 _09759_/Y sky130_fd_sc_hd__inv_2
XPHY_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13291__A1 _20551_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12770_ _20797_/Q _12765_/X _12670_/X _12766_/X vssd1 vssd1 vccd1 vccd1 _20797_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18754__A0 _18753_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_215_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11721_ _11721_/A vssd1 vssd1 vccd1 vccd1 _11721_/X sky130_fd_sc_hd__buf_1
XPHY_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20919_ _20949_/CLK _20919_/D repeater272/X vssd1 vssd1 vccd1 vccd1 _20919_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_215_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14440_ _14438_/Y _20212_/Q _14439_/Y _20227_/Q vssd1 vssd1 vccd1 vccd1 _14440_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11652_ _19112_/X vssd1 vssd1 vccd1 vccd1 _11652_/X sky130_fd_sc_hd__buf_1
XPHY_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10603_ _21341_/Q _10601_/Y _21333_/Q _10602_/Y vssd1 vssd1 vccd1 vccd1 _10603_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14371_ _14461_/C _14483_/A vssd1 vssd1 vccd1 vccd1 _14372_/B sky130_fd_sc_hd__or2_1
XFILLER_80_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11583_ _21125_/Q _11583_/B vssd1 vssd1 vccd1 vccd1 _21125_/D sky130_fd_sc_hd__and2_1
XPHY_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16110_ _16119_/A vssd1 vssd1 vccd1 vccd1 _16121_/A sky130_fd_sc_hd__inv_2
XFILLER_196_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13322_ _13322_/A vssd1 vssd1 vccd1 vccd1 _13322_/X sky130_fd_sc_hd__buf_1
XFILLER_127_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10534_ _10534_/A _10534_/B vssd1 vssd1 vccd1 vccd1 _10665_/A sky130_fd_sc_hd__or2_1
X_17090_ _21342_/Q _20737_/Q vssd1 vssd1 vccd1 vccd1 _17090_/X sky130_fd_sc_hd__and2_2
XPHY_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16041_ _19514_/Q _16035_/X _16006_/X _16037_/X vssd1 vssd1 vccd1 vccd1 _19514_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19157__S1 _21017_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10465_ _21295_/Q vssd1 vssd1 vccd1 vccd1 _10771_/A sky130_fd_sc_hd__inv_2
X_13253_ _20565_/Q _13248_/X _13173_/X _13249_/X vssd1 vssd1 vccd1 vccd1 _20565_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_183_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12204_ _12193_/X _12204_/B _12204_/C _12204_/D vssd1 vssd1 vccd1 vccd1 _12204_/X
+ sky130_fd_sc_hd__and4b_1
X_10396_ _21359_/Q _10394_/Y _10395_/X _10275_/B vssd1 vssd1 vccd1 vccd1 _21359_/D
+ sky130_fd_sc_hd__o211a_1
X_13184_ _11974_/X _16525_/A _13184_/S vssd1 vssd1 vccd1 vccd1 _20598_/D sky130_fd_sc_hd__mux2_1
XFILLER_123_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19800_ _19820_/CLK _19800_/D vssd1 vssd1 vccd1 vccd1 _19800_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17076__A _21135_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12135_ _12318_/A _20379_/Q _12325_/A _20386_/Q vssd1 vssd1 vccd1 vccd1 _12135_/X
+ sky130_fd_sc_hd__o22a_1
X_17992_ _20418_/Q vssd1 vssd1 vccd1 vccd1 _17992_/Y sky130_fd_sc_hd__inv_2
XFILLER_151_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16943_ _16956_/A _16943_/B vssd1 vssd1 vccd1 vccd1 _16943_/Y sky130_fd_sc_hd__nor2_1
X_19731_ _19789_/CLK _19731_/D vssd1 vssd1 vccd1 vccd1 _19731_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12066_ _20953_/Q _12061_/Y _20963_/Q _12062_/Y _12065_/X vssd1 vssd1 vccd1 vccd1
+ _12087_/A sky130_fd_sc_hd__o221a_1
XFILLER_1_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10868__B1 _09676_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11017_ _11017_/A _11017_/B vssd1 vssd1 vccd1 vccd1 _21244_/D sky130_fd_sc_hd__or2_1
XFILLER_38_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19662_ _19811_/CLK _19662_/D vssd1 vssd1 vccd1 vccd1 _19662_/Q sky130_fd_sc_hd__dfxtp_1
X_16874_ _16872_/Y _16873_/X _16848_/X vssd1 vssd1 vccd1 vccd1 _16874_/X sky130_fd_sc_hd__o21a_1
XANTENNA__14407__A2_N _20025_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15825_ _15825_/A vssd1 vssd1 vccd1 vccd1 _15825_/X sky130_fd_sc_hd__buf_1
X_18613_ _18848_/A0 _17831_/Y _18666_/S vssd1 vssd1 vccd1 vccd1 _18613_/X sky130_fd_sc_hd__mux2_1
XFILLER_237_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19593_ _20890_/CLK _19593_/D vssd1 vssd1 vccd1 vccd1 _19593_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_231_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15324__A _15330_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18544_ _18845_/A0 _10490_/Y _18896_/S vssd1 vssd1 vccd1 vccd1 _18544_/X sky130_fd_sc_hd__mux2_1
X_15756_ _15756_/A _15756_/B _16297_/C vssd1 vssd1 vccd1 vccd1 _15768_/A sky130_fd_sc_hd__or3_4
XFILLER_33_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12085__A2 _12083_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12968_ _12968_/A _16526_/A _12968_/C vssd1 vssd1 vccd1 vccd1 _12968_/X sky130_fd_sc_hd__and3_1
XFILLER_61_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14707_ _20159_/Q _14704_/X _12849_/A _14706_/X vssd1 vssd1 vccd1 vccd1 _20159_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_205_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11919_ _11176_/B _11136_/X _15609_/B _21003_/Q _11943_/A vssd1 vssd1 vccd1 vccd1
+ _11926_/B sky130_fd_sc_hd__a221o_1
X_18475_ _18848_/A0 _14139_/Y _18884_/S vssd1 vssd1 vccd1 vccd1 _18475_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15687_ _15722_/A _16311_/B _15778_/C vssd1 vssd1 vccd1 vccd1 _15696_/A sky130_fd_sc_hd__or3_4
XPHY_4490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21226__RESET_B repeater249/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12899_ _12899_/A _13261_/A vssd1 vssd1 vccd1 vccd1 _12934_/A sky130_fd_sc_hd__or2_2
XFILLER_220_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17426_ _17773_/B vssd1 vssd1 vccd1 vccd1 _17631_/B sky130_fd_sc_hd__clkbuf_2
X_14638_ _13738_/X _14637_/A _20185_/Q _14637_/Y _14599_/X vssd1 vssd1 vccd1 vccd1
+ _20185_/D sky130_fd_sc_hd__o221a_1
XFILLER_220_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17357_ _19576_/Q vssd1 vssd1 vccd1 vccd1 _17357_/Y sky130_fd_sc_hd__inv_2
X_14569_ _14569_/A _14648_/A vssd1 vssd1 vccd1 vccd1 _14570_/B sky130_fd_sc_hd__or2_2
XFILLER_147_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16308_ _19384_/Q _16305_/X _16291_/X _16306_/X vssd1 vssd1 vccd1 vccd1 _19384_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12793__B1 _09655_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17288_ _11670_/Y _17151_/X _17287_/Y _17139_/A vssd1 vssd1 vccd1 vccd1 _17288_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_109_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19027_ _16880_/X _20842_/Q _19058_/S vssd1 vssd1 vccd1 vccd1 _19949_/D sky130_fd_sc_hd__mux2_1
X_16239_ _19418_/Q _16230_/X _16006_/X _16233_/X vssd1 vssd1 vccd1 vccd1 _19418_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19148__S1 _21017_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20179__RESET_B repeater200/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20108__RESET_B repeater264/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19929_ _21238_/CLK _19929_/D repeater256/X vssd1 vssd1 vccd1 vccd1 _19929_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_205_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13019__A _13040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09613_ _20878_/Q _20877_/Q vssd1 vssd1 vccd1 vccd1 _09615_/C sky130_fd_sc_hd__or2_1
XFILLER_83_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_244_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14470__B1 _14469_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20704_ _21349_/CLK _20704_/D repeater210/X vssd1 vssd1 vccd1 vccd1 _20704_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_200_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20635_ _21486_/CLK _20635_/D repeater198/X vssd1 vssd1 vccd1 vccd1 _20635_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_149_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20566_ _20592_/CLK _20566_/D repeater260/X vssd1 vssd1 vccd1 vccd1 _20566_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_165_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19139__S1 _21017_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20497_ _20929_/CLK _20497_/D repeater265/X vssd1 vssd1 vccd1 vccd1 _20497_/Q sky130_fd_sc_hd__dfrtp_2
X_10250_ _21353_/Q vssd1 vssd1 vccd1 vccd1 _10346_/A sky130_fd_sc_hd__inv_2
XFILLER_180_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10181_ _10159_/A _10159_/B _10177_/X _10179_/Y vssd1 vssd1 vccd1 vccd1 _21398_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_79_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21118_ _21120_/CLK _21118_/D repeater233/X vssd1 vssd1 vccd1 vccd1 _21118_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_59_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21049_ _21164_/CLK _21049_/D repeater227/X vssd1 vssd1 vccd1 vccd1 _21049_/Q sky130_fd_sc_hd__dfrtp_1
X_13940_ _20638_/Q _14011_/A _20662_/Q _13894_/A vssd1 vssd1 vccd1 vccd1 _13940_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_207_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_219_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13871_ _20300_/Q vssd1 vssd1 vccd1 vccd1 _14016_/A sky130_fd_sc_hd__inv_2
XFILLER_234_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15610_ _15610_/A _16215_/B _16344_/C vssd1 vssd1 vccd1 vccd1 _15618_/A sky130_fd_sc_hd__or3_4
X_12822_ _12847_/A vssd1 vssd1 vccd1 vccd1 _12850_/A sky130_fd_sc_hd__inv_2
X_16590_ _16503_/A _16501_/X _16510_/Y vssd1 vssd1 vccd1 vccd1 _16590_/X sky130_fd_sc_hd__o21a_1
XFILLER_234_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18727__A0 _18726_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15541_ _19750_/Q _15536_/X _15526_/X _15537_/X vssd1 vssd1 vccd1 vccd1 _19750_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12753_ _12753_/A _13047_/B _13188_/C vssd1 vssd1 vccd1 vccd1 _17201_/A sky130_fd_sc_hd__or3_4
XFILLER_199_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19050__S _19058_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11704_ _11704_/A vssd1 vssd1 vccd1 vccd1 _11704_/X sky130_fd_sc_hd__buf_1
XPHY_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18260_ _18259_/X _12187_/Y _18787_/S vssd1 vssd1 vccd1 vccd1 _18260_/X sky130_fd_sc_hd__mux2_1
XPHY_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15472_ _19781_/Q _15468_/X _15469_/X _15471_/X vssd1 vssd1 vccd1 vccd1 _19781_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_230_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12684_ _20827_/Q _12679_/X _09638_/X _12680_/X vssd1 vssd1 vccd1 vccd1 _20827_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17211_ _17211_/A vssd1 vssd1 vccd1 vccd1 _17211_/X sky130_fd_sc_hd__clkbuf_2
XPHY_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14423_ _21466_/Q _14351_/A _14421_/Y _20029_/Q _14422_/X vssd1 vssd1 vccd1 vccd1
+ _14434_/A sky130_fd_sc_hd__o221a_1
XPHY_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_230_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18191_ _18190_/X _14584_/A _18748_/S vssd1 vssd1 vccd1 vccd1 _18191_/X sky130_fd_sc_hd__mux2_1
X_11635_ _14813_/C _11631_/B _11613_/A _11638_/A vssd1 vssd1 vccd1 vccd1 _21104_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_118_HCLK_A clkbuf_opt_3_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14764__B2 _20130_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17142_ _17142_/A vssd1 vssd1 vccd1 vccd1 _17162_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__12775__B1 _09626_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14354_ _20214_/Q vssd1 vssd1 vccd1 vccd1 _14499_/A sky130_fd_sc_hd__inv_2
XPHY_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11566_ _11566_/A vssd1 vssd1 vccd1 vccd1 _11566_/X sky130_fd_sc_hd__buf_1
XPHY_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13305_ _20543_/Q _13300_/X _13146_/X _13302_/X vssd1 vssd1 vccd1 vccd1 _20543_/D
+ sky130_fd_sc_hd__a22o_1
X_17073_ _17076_/C _17073_/B _19889_/Q vssd1 vssd1 vccd1 vccd1 _19885_/D sky130_fd_sc_hd__nor3_1
X_10517_ _20682_/Q vssd1 vssd1 vccd1 vccd1 _10517_/Y sky130_fd_sc_hd__inv_2
XFILLER_143_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14285_ _14276_/Y _14284_/X _14276_/Y _14284_/X vssd1 vssd1 vccd1 vccd1 _14302_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_11497_ _11497_/A vssd1 vssd1 vccd1 vccd1 _11498_/A sky130_fd_sc_hd__inv_2
XFILLER_170_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16024_ _19525_/Q _16021_/X _15758_/X _16023_/X vssd1 vssd1 vccd1 vccd1 _19525_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_6_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13236_ _20575_/Q _13233_/X _13154_/X _13234_/X vssd1 vssd1 vccd1 vccd1 _20575_/D
+ sky130_fd_sc_hd__a22o_1
X_10448_ _21279_/Q vssd1 vssd1 vccd1 vccd1 _10756_/A sky130_fd_sc_hd__inv_2
XFILLER_152_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20272__RESET_B repeater264/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13167_ _13167_/A vssd1 vssd1 vccd1 vccd1 _13167_/X sky130_fd_sc_hd__buf_1
X_10379_ _10283_/A _10283_/B _10377_/Y _10405_/B vssd1 vssd1 vccd1 vccd1 _21368_/D
+ sky130_fd_sc_hd__a211oi_4
XANTENNA__20201__RESET_B repeater193/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12118_ _20974_/Q vssd1 vssd1 vccd1 vccd1 _12327_/A sky130_fd_sc_hd__inv_2
XFILLER_97_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17975_ _17975_/A _17978_/B vssd1 vssd1 vccd1 vccd1 _17975_/Y sky130_fd_sc_hd__nor2_1
XFILLER_111_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13098_ _13098_/A vssd1 vssd1 vccd1 vccd1 _13098_/X sky130_fd_sc_hd__buf_1
Xclkbuf_3_0_0_HCLK clkbuf_3_1_0_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_1_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_242_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19714_ _21222_/CLK _19714_/D vssd1 vssd1 vccd1 vccd1 _19714_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12049_ _20973_/Q vssd1 vssd1 vccd1 vccd1 _12326_/A sky130_fd_sc_hd__inv_2
X_16926_ _16926_/A vssd1 vssd1 vccd1 vccd1 _16931_/B sky130_fd_sc_hd__inv_2
XANTENNA__10305__A2 _20732_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19645_ _20327_/CLK _19645_/D vssd1 vssd1 vccd1 vccd1 _19645_/Q sky130_fd_sc_hd__dfxtp_1
X_16857_ _16861_/B vssd1 vssd1 vccd1 vccd1 _16863_/B sky130_fd_sc_hd__inv_2
XFILLER_65_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21407__RESET_B repeater252/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15808_ _15808_/A vssd1 vssd1 vccd1 vccd1 _15808_/X sky130_fd_sc_hd__buf_1
XFILLER_81_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19576_ _20890_/CLK _19576_/D vssd1 vssd1 vccd1 vccd1 _19576_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16788_ _16791_/B _16787_/X _16779_/X vssd1 vssd1 vccd1 vccd1 _16788_/X sky130_fd_sc_hd__o21a_1
XFILLER_92_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18527_ _18526_/X _14939_/Y _18907_/S vssd1 vssd1 vccd1 vccd1 _18527_/X sky130_fd_sc_hd__mux2_1
X_15739_ _19656_/Q _15736_/X _15701_/X _15737_/X vssd1 vssd1 vccd1 vccd1 _19656_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_179_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18458_ _18845_/A0 _13789_/Y _18896_/S vssd1 vssd1 vccd1 vccd1 _18458_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18084__B _18084_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_5_0_HCLK_A clkbuf_3_5_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17409_ _19697_/Q vssd1 vssd1 vccd1 vccd1 _17409_/Y sky130_fd_sc_hd__inv_2
X_18389_ _18388_/X _14889_/Y _18907_/S vssd1 vssd1 vccd1 vccd1 _18389_/X sky130_fd_sc_hd__mux2_1
XFILLER_187_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20420_ _20957_/CLK _20420_/D repeater187/X vssd1 vssd1 vccd1 vccd1 _20420_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__09631__B1 _09630_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20351_ _20480_/CLK _20351_/D repeater183/X vssd1 vssd1 vccd1 vccd1 _20351_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_162_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18304__S _18906_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20282_ _20286_/CLK _20282_/D repeater264/X vssd1 vssd1 vccd1 vccd1 _20282_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_162_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18709__A0 _17281_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19760__CLK _19765_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11420_ _11420_/A vssd1 vssd1 vccd1 vccd1 _11420_/X sky130_fd_sc_hd__buf_1
X_20618_ _20622_/CLK _20618_/D repeater195/X vssd1 vssd1 vccd1 vccd1 _20618_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_20_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16499__A1 _16495_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20712__RESET_B repeater254/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11351_ _21172_/Q vssd1 vssd1 vccd1 vccd1 _11390_/C sky130_fd_sc_hd__buf_1
X_20549_ _20947_/CLK _20549_/D repeater266/X vssd1 vssd1 vccd1 vccd1 _20549_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__18214__S _18902_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10302_ _10286_/A _20730_/Q _21358_/Q _17901_/A _10301_/X vssd1 vssd1 vccd1 vccd1
+ _10307_/C sky130_fd_sc_hd__o221a_1
X_14070_ _14070_/A _14070_/B vssd1 vssd1 vccd1 vccd1 _14228_/A sky130_fd_sc_hd__or2_2
XFILLER_125_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11282_ _20908_/Q _11310_/C _11299_/C vssd1 vssd1 vccd1 vccd1 _11290_/C sky130_fd_sc_hd__or3_4
XFILLER_134_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13021_ _13041_/A vssd1 vssd1 vccd1 vccd1 _13021_/X sky130_fd_sc_hd__buf_1
X_10233_ _21370_/Q vssd1 vssd1 vccd1 vccd1 _10285_/A sky130_fd_sc_hd__inv_2
XFILLER_126_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_239_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input44_A HWDATA[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10164_ _10164_/A vssd1 vssd1 vccd1 vccd1 _10164_/Y sky130_fd_sc_hd__inv_2
XFILLER_126_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19045__S _19046_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17760_ _19348_/Q vssd1 vssd1 vccd1 vccd1 _17760_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14972_ _14972_/A vssd1 vssd1 vccd1 vccd1 _14972_/Y sky130_fd_sc_hd__inv_2
X_10095_ _20789_/Q vssd1 vssd1 vccd1 vccd1 _10095_/Y sky130_fd_sc_hd__inv_2
XANTENNA__09689__B1 _09688_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16711_ _16711_/A vssd1 vssd1 vccd1 vccd1 _16718_/A sky130_fd_sc_hd__clkbuf_2
X_13923_ _20652_/Q vssd1 vssd1 vccd1 vccd1 _13923_/Y sky130_fd_sc_hd__inv_2
XFILLER_235_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17691_ _19612_/Q vssd1 vssd1 vccd1 vccd1 _17691_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18884__S _18884_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16642_ _19856_/Q _15290_/B _15291_/B vssd1 vssd1 vccd1 vccd1 _16642_/X sky130_fd_sc_hd__a21bo_1
X_19430_ _20137_/CLK _19430_/D vssd1 vssd1 vccd1 vccd1 _19430_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13854_ _20307_/Q vssd1 vssd1 vccd1 vccd1 _13883_/A sky130_fd_sc_hd__inv_2
XANTENNA__19966__RESET_B repeater185/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12805_ _20776_/Q _12803_/X _11736_/X _12804_/X vssd1 vssd1 vccd1 vccd1 _20776_/D
+ sky130_fd_sc_hd__a22o_1
X_16573_ _16573_/A vssd1 vssd1 vccd1 vccd1 _16573_/Y sky130_fd_sc_hd__inv_2
XFILLER_204_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13106__B _13106_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19361_ _21222_/CLK _19361_/D vssd1 vssd1 vccd1 vccd1 _19361_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13785_ _13780_/Y _20194_/Q _20605_/Q _14572_/A _13784_/X vssd1 vssd1 vccd1 vccd1
+ _13786_/D sky130_fd_sc_hd__o221a_1
XFILLER_27_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10997_ _15375_/A _10996_/X _15375_/A _10996_/X vssd1 vssd1 vccd1 vccd1 _11012_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_31_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18312_ _18845_/A0 _10513_/Y _18896_/S vssd1 vssd1 vccd1 vccd1 _18312_/X sky130_fd_sc_hd__mux2_1
X_15524_ _15793_/A vssd1 vssd1 vccd1 vccd1 _15524_/X sky130_fd_sc_hd__buf_1
XFILLER_16_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19292_ _19776_/CLK _19292_/D vssd1 vssd1 vccd1 vccd1 _19292_/Q sky130_fd_sc_hd__dfxtp_1
X_12736_ _12740_/B vssd1 vssd1 vccd1 vccd1 _14686_/B sky130_fd_sc_hd__inv_2
XFILLER_30_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09600__A _20888_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18243_ _19131_/X _20161_/Q _18249_/S vssd1 vssd1 vccd1 vccd1 _18243_/X sky130_fd_sc_hd__mux2_1
XFILLER_176_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15455_ _19788_/Q _15449_/X _15454_/X _15452_/X vssd1 vssd1 vccd1 vccd1 _19788_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12667_ _20837_/Q _12662_/X _12666_/X _12664_/X vssd1 vssd1 vccd1 vccd1 _20837_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14406_ _21471_/Q vssd1 vssd1 vccd1 vccd1 _14406_/Y sky130_fd_sc_hd__inv_2
XPHY_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11618_ _11636_/A _21110_/Q vssd1 vssd1 vccd1 vccd1 _11618_/Y sky130_fd_sc_hd__nor2_1
X_18174_ _17281_/X _18100_/Y _18874_/S vssd1 vssd1 vccd1 vccd1 _18174_/X sky130_fd_sc_hd__mux2_1
XFILLER_156_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19220__S0 _20130_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12212__A2 _20502_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15386_ _15663_/A vssd1 vssd1 vccd1 vccd1 _15386_/X sky130_fd_sc_hd__buf_1
XFILLER_128_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12598_ _20874_/Q _12594_/X _18226_/X _12595_/X vssd1 vssd1 vccd1 vccd1 _20874_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17125_ _19349_/Q vssd1 vssd1 vccd1 vccd1 _17125_/Y sky130_fd_sc_hd__inv_2
XPHY_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14337_ _20228_/Q vssd1 vssd1 vccd1 vccd1 _14461_/C sky130_fd_sc_hd__inv_2
XFILLER_7_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11549_ _11549_/A vssd1 vssd1 vccd1 vccd1 _17387_/A sky130_fd_sc_hd__buf_1
XFILLER_144_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12961__A _12961_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17056_ _19845_/Q _19846_/Q _19847_/Q vssd1 vssd1 vccd1 vccd1 _19845_/D sky130_fd_sc_hd__o21ba_1
XFILLER_132_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14268_ _14268_/A vssd1 vssd1 vccd1 vccd1 _14268_/X sky130_fd_sc_hd__buf_1
XFILLER_144_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16007_ _19530_/Q _16000_/X _16006_/X _16002_/X vssd1 vssd1 vccd1 vccd1 _19530_/D
+ sky130_fd_sc_hd__a22o_1
X_13219_ input47/X vssd1 vssd1 vccd1 vccd1 _13219_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_143_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14199_ _20278_/Q _14198_/Y _14183_/X _14089_/B vssd1 vssd1 vccd1 vccd1 _20278_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_140_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17958_ _20829_/Q vssd1 vssd1 vccd1 vccd1 _17958_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16909_ _16909_/A vssd1 vssd1 vccd1 vccd1 _16914_/B sky130_fd_sc_hd__inv_2
XFILLER_238_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18794__S _18929_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17889_ _17889_/A vssd1 vssd1 vccd1 vccd1 _18020_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_26_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19628_ _21040_/CLK _19628_/D vssd1 vssd1 vccd1 vccd1 _19628_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_226_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13779__A2 _14566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19559_ _19706_/CLK _19559_/D vssd1 vssd1 vccd1 vccd1 _19559_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15925__B1 _15893_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21452_ _21452_/CLK _21452_/D repeater247/X vssd1 vssd1 vccd1 vccd1 _21452_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_119_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19211__S0 _20132_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_101_HCLK_A clkbuf_4_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20194__RESET_B repeater193/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20403_ _20809_/CLK _20403_/D repeater188/X vssd1 vssd1 vccd1 vccd1 _20403_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_147_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_164_HCLK_A clkbuf_opt_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21383_ _21390_/CLK _21383_/D repeater214/X vssd1 vssd1 vccd1 vccd1 _21383_/Q sky130_fd_sc_hd__dfrtp_1
X_20334_ _20809_/CLK _20334_/D repeater188/X vssd1 vssd1 vccd1 vccd1 _20334_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_190_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13164__B1 _13163_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_227_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20265_ _20286_/CLK _20265_/D repeater265/X vssd1 vssd1 vccd1 vccd1 _20265_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_163_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12911__B1 _12663_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20196_ _20626_/CLK _20196_/D repeater193/X vssd1 vssd1 vccd1 vccd1 _20196_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_142_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21329__RESET_B repeater204/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17174__A _20497_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19278__S0 _19280_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13207__A _13217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10920_ _21206_/Q vssd1 vssd1 vccd1 vccd1 _10920_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10851_ _18280_/X _10847_/X _21274_/Q _10849_/X vssd1 vssd1 vccd1 vccd1 _21274_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_32_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18209__S _18787_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20964__RESET_B repeater186/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13570_ _20414_/Q _13566_/X _13487_/X _13567_/X vssd1 vssd1 vccd1 vccd1 _20414_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_241_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10782_ _10782_/A _10790_/A vssd1 vssd1 vccd1 vccd1 _10783_/B sky130_fd_sc_hd__or2_2
XFILLER_201_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12521_ _12521_/A vssd1 vssd1 vccd1 vccd1 _12521_/X sky130_fd_sc_hd__buf_1
XFILLER_13_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15240_ _15238_/Y _20072_/Q _15239_/Y _20062_/Q vssd1 vssd1 vccd1 vccd1 _15240_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12452_ _20939_/Q _12451_/Y _12448_/X _12429_/B vssd1 vssd1 vccd1 vccd1 _20939_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__19202__S0 _19275_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_71_HCLK clkbuf_opt_6_HCLK/X vssd1 vssd1 vccd1 vccd1 _19907_/CLK sky130_fd_sc_hd__clkbuf_16
X_11403_ _11403_/A vssd1 vssd1 vccd1 vccd1 _11420_/A sky130_fd_sc_hd__inv_2
XFILLER_184_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15171_ _15193_/A vssd1 vssd1 vccd1 vccd1 _15179_/A sky130_fd_sc_hd__buf_2
X_12383_ _12383_/A vssd1 vssd1 vccd1 vccd1 _12383_/Y sky130_fd_sc_hd__inv_2
XFILLER_126_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11953__A1 _21006_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14122_ _20543_/Q vssd1 vssd1 vccd1 vccd1 _14122_/Y sky130_fd_sc_hd__inv_2
X_11334_ _21173_/Q _21172_/Q _11350_/A vssd1 vssd1 vccd1 vccd1 _11362_/C sky130_fd_sc_hd__or3_1
XFILLER_114_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_23_HCLK_A clkbuf_4_9_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18879__S _18879_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13155__B1 _13154_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18930_ _18929_/X _19276_/X _18930_/S vssd1 vssd1 vccd1 vccd1 _18930_/X sky130_fd_sc_hd__mux2_2
X_14053_ _20275_/Q vssd1 vssd1 vccd1 vccd1 _14085_/A sky130_fd_sc_hd__inv_2
XFILLER_125_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_86_HCLK_A clkbuf_4_12_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11265_ _20904_/Q _20903_/Q _20902_/Q _20901_/Q vssd1 vssd1 vccd1 vccd1 _11299_/C
+ sky130_fd_sc_hd__or4_4
XFILLER_141_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13004_ _20690_/Q _12995_/X _13003_/X _12997_/X vssd1 vssd1 vccd1 vccd1 _20690_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_122_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10216_ _10216_/A vssd1 vssd1 vccd1 vccd1 _10216_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14301__A1_N _20122_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18861_ _17277_/Y _17276_/Y _18926_/S vssd1 vssd1 vccd1 vccd1 _18861_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11196_ _21215_/Q _11191_/X _10896_/X _11193_/X vssd1 vssd1 vccd1 vccd1 _21215_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_121_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17812_ _17812_/A _17812_/B vssd1 vssd1 vccd1 vccd1 _17812_/Y sky130_fd_sc_hd__nor2_1
XFILLER_121_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10147_ _10147_/A _10227_/C _10147_/C vssd1 vssd1 vccd1 vccd1 _21406_/D sky130_fd_sc_hd__nor3_1
XANTENNA__19269__S0 _20130_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18792_ _18791_/X _17444_/Y _18927_/S vssd1 vssd1 vccd1 vccd1 _18792_/X sky130_fd_sc_hd__mux2_1
XFILLER_153_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14955_ _14989_/A vssd1 vssd1 vccd1 vccd1 _15025_/C sky130_fd_sc_hd__clkbuf_2
X_17743_ _19429_/Q vssd1 vssd1 vccd1 vccd1 _17743_/Y sky130_fd_sc_hd__inv_2
X_10078_ _10078_/A vssd1 vssd1 vccd1 vccd1 _10147_/A sky130_fd_sc_hd__inv_2
XFILLER_48_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13906_ _13903_/Y _20302_/Q _20645_/Q _13876_/C _13905_/X vssd1 vssd1 vccd1 vccd1
+ _13914_/B sky130_fd_sc_hd__o221a_1
XFILLER_236_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14886_ _20584_/Q vssd1 vssd1 vccd1 vccd1 _14886_/Y sky130_fd_sc_hd__inv_2
X_17674_ _19524_/Q vssd1 vssd1 vccd1 vccd1 _17674_/Y sky130_fd_sc_hd__inv_2
X_19413_ _21001_/CLK _19413_/D vssd1 vssd1 vccd1 vccd1 _19413_/Q sky130_fd_sc_hd__dfxtp_1
X_16625_ _11327_/X _16507_/B _19998_/Q _16624_/Y vssd1 vssd1 vccd1 vccd1 _19998_/D
+ sky130_fd_sc_hd__a31o_1
X_13837_ _13837_/A _13837_/B _13837_/C _13837_/D vssd1 vssd1 vccd1 vccd1 _14597_/A
+ sky130_fd_sc_hd__and4_1
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16556_ _16556_/A _16556_/B vssd1 vssd1 vccd1 vccd1 _16556_/Y sky130_fd_sc_hd__nor2_1
X_19344_ _20137_/CLK _19344_/D vssd1 vssd1 vccd1 vccd1 _19344_/Q sky130_fd_sc_hd__dfxtp_1
X_13768_ _20629_/Q vssd1 vssd1 vccd1 vccd1 _13768_/Y sky130_fd_sc_hd__inv_2
XFILLER_204_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12719_ _20809_/Q vssd1 vssd1 vccd1 vccd1 _16915_/A sky130_fd_sc_hd__clkbuf_2
X_15507_ _15516_/A vssd1 vssd1 vccd1 vccd1 _15507_/X sky130_fd_sc_hd__buf_1
X_19275_ _17105_/Y _17106_/Y _17107_/Y _17108_/Y _19275_/S0 _21004_/Q vssd1 vssd1
+ vccd1 vccd1 _19275_/X sky130_fd_sc_hd__mux4_2
X_16487_ _16487_/A vssd1 vssd1 vccd1 vccd1 _18927_/S sky130_fd_sc_hd__inv_4
X_13699_ _13706_/A vssd1 vssd1 vccd1 vccd1 _13699_/X sky130_fd_sc_hd__buf_1
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18226_ _20850_/Q input30/X _18236_/S vssd1 vssd1 vccd1 vccd1 _18226_/X sky130_fd_sc_hd__mux2_1
X_15438_ _19796_/Q _15434_/X _15383_/X _15436_/X vssd1 vssd1 vccd1 vccd1 _19796_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_129_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13394__B1 _13265_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15369_ _19824_/Q _15366_/X _15350_/X _15367_/X vssd1 vssd1 vccd1 vccd1 _19824_/D
+ sky130_fd_sc_hd__a22o_1
X_18157_ _18005_/Y _20760_/Q _18775_/S vssd1 vssd1 vccd1 vccd1 _18157_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17108_ _19398_/Q vssd1 vssd1 vccd1 vccd1 _17108_/Y sky130_fd_sc_hd__inv_2
X_18088_ _18662_/X _17951_/A _18664_/X _17952_/A vssd1 vssd1 vccd1 vccd1 _18090_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_172_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17039_ _21410_/Q vssd1 vssd1 vccd1 vccd1 _17039_/Y sky130_fd_sc_hd__inv_2
X_09930_ input38/X vssd1 vssd1 vccd1 vccd1 _16342_/A sky130_fd_sc_hd__buf_2
XFILLER_172_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13697__A1 _20341_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20050_ _20066_/CLK _20050_/D repeater281/X vssd1 vssd1 vccd1 vccd1 _20050_/Q sky130_fd_sc_hd__dfrtp_2
X_09861_ _10842_/A _09861_/B vssd1 vssd1 vccd1 vccd1 _15314_/A sky130_fd_sc_hd__or2_4
XFILLER_86_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09792_ _09792_/A vssd1 vssd1 vccd1 vccd1 _09804_/A sky130_fd_sc_hd__buf_1
XFILLER_97_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater154 _18617_/S vssd1 vssd1 vccd1 vccd1 _18898_/S sky130_fd_sc_hd__buf_8
XFILLER_238_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater165 _18874_/S vssd1 vssd1 vccd1 vccd1 _18835_/S sky130_fd_sc_hd__buf_8
XFILLER_213_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13027__A _13041_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater176 _18644_/S vssd1 vssd1 vccd1 vccd1 _18849_/S sky130_fd_sc_hd__clkbuf_8
XPHY_4308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater187 repeater271/X vssd1 vssd1 vccd1 vccd1 repeater187/X sky130_fd_sc_hd__buf_8
X_20952_ _20957_/CLK _20952_/D repeater271/X vssd1 vssd1 vccd1 vccd1 _20952_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater198 repeater199/X vssd1 vssd1 vccd1 vccd1 repeater198/X sky130_fd_sc_hd__buf_8
XFILLER_199_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20883_ _21444_/CLK _20883_/D repeater243/X vssd1 vssd1 vccd1 vccd1 _20883_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_53_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16338__A _16338_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20375__RESET_B repeater186/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_94_HCLK clkbuf_4_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20947_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_42_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21435_ _21438_/CLK _21435_/D repeater239/X vssd1 vssd1 vccd1 vccd1 _21435_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17169__A _17169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16323__B1 _16014_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21366_ _21366_/CLK _21366_/D repeater254/X vssd1 vssd1 vccd1 vccd1 _21366_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18699__S _18909_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13137__B1 _12932_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_0_HCLK clkbuf_opt_0_HCLK/A vssd1 vssd1 vccd1 vccd1 _19777_/CLK sky130_fd_sc_hd__clkbuf_16
X_20317_ _20322_/CLK _20317_/D repeater262/X vssd1 vssd1 vccd1 vccd1 _20317_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_89_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21297_ _21357_/CLK _21297_/D repeater209/X vssd1 vssd1 vccd1 vccd1 _21297_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_150_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11050_ _11050_/A _14309_/A vssd1 vssd1 vccd1 vccd1 _11100_/A sky130_fd_sc_hd__or2_2
XFILLER_89_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20248_ _21147_/CLK _20248_/D repeater215/X vssd1 vssd1 vccd1 vccd1 _20248_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__21163__RESET_B repeater226/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10001_ _09999_/X _20017_/Q _20018_/Q vssd1 vssd1 vccd1 vccd1 _10001_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_49_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20179_ _21485_/CLK _20179_/D repeater200/X vssd1 vssd1 vccd1 vccd1 _20179_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_191_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14740_ _13600_/X _11076_/X _14740_/S vssd1 vssd1 vccd1 vccd1 _20138_/D sky130_fd_sc_hd__mux2_1
XFILLER_218_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11952_ _11952_/A vssd1 vssd1 vccd1 vccd1 _11955_/A sky130_fd_sc_hd__inv_2
XFILLER_45_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17587__C1 _17586_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_217_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17989__D _17989_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10903_ _21123_/Q _21122_/Q _21124_/Q _21121_/Q _21125_/Q vssd1 vssd1 vccd1 vccd1
+ _11584_/C sky130_fd_sc_hd__a41o_1
X_14671_ _14659_/A _14663_/Y _14659_/A _14663_/Y vssd1 vssd1 vccd1 vccd1 _20172_/D
+ sky130_fd_sc_hd__o2bb2a_1
X_11883_ _11883_/A vssd1 vssd1 vccd1 vccd1 _11883_/X sky130_fd_sc_hd__buf_1
XFILLER_233_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11680__A _12544_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16410_ _19331_/Q _16406_/X _16200_/X _16408_/X vssd1 vssd1 vccd1 vccd1 _19331_/D
+ sky130_fd_sc_hd__a22o_1
X_13622_ _20386_/Q _13619_/X _13475_/X _13620_/X vssd1 vssd1 vccd1 vccd1 _20386_/D
+ sky130_fd_sc_hd__a22o_1
X_17390_ _17390_/A vssd1 vssd1 vccd1 vccd1 _17390_/X sky130_fd_sc_hd__clkbuf_2
X_10834_ _21282_/Q _10833_/Y _10830_/X _10760_/B vssd1 vssd1 vccd1 vccd1 _21282_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09816__B1 input74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16341_ _19367_/Q _16334_/X _16340_/X _16336_/X vssd1 vssd1 vccd1 vccd1 _19367_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_198_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13553_ input56/X vssd1 vssd1 vccd1 vccd1 _13553_/X sky130_fd_sc_hd__buf_4
XFILLER_13_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10765_ _10765_/A _10765_/B vssd1 vssd1 vccd1 vccd1 _10818_/A sky130_fd_sc_hd__or2_1
XFILLER_158_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20045__RESET_B repeater276/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12504_ _12504_/A _12504_/B vssd1 vssd1 vccd1 vccd1 _16689_/C sky130_fd_sc_hd__or2_1
X_19060_ _21191_/Q _21133_/Q _19910_/Q vssd1 vssd1 vccd1 vccd1 _19060_/X sky130_fd_sc_hd__mux2_1
X_16272_ _19400_/Q _16269_/X _16123_/X _16270_/X vssd1 vssd1 vccd1 vccd1 _19400_/D
+ sky130_fd_sc_hd__a22o_1
X_13484_ _20452_/Q _13481_/X _13482_/X _13483_/X vssd1 vssd1 vccd1 vccd1 _20452_/D
+ sky130_fd_sc_hd__a22o_1
X_10696_ _10653_/A _10653_/B _10685_/X _10693_/Y vssd1 vssd1 vccd1 vccd1 _21324_/D
+ sky130_fd_sc_hd__a211oi_2
X_15223_ _15222_/Y _20060_/Q _20472_/Q _15066_/A vssd1 vssd1 vccd1 vccd1 _15223_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__13376__B1 _13163_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18011_ _18158_/X _17907_/X _18269_/X _17908_/X vssd1 vssd1 vccd1 vccd1 _18014_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17079__A _17174_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12435_ _20947_/Q _12434_/Y _12407_/C _12434_/A _12411_/X vssd1 vssd1 vccd1 vccd1
+ _20947_/D sky130_fd_sc_hd__o221a_1
XFILLER_138_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_repeater146_A _19026_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15154_ _20434_/Q vssd1 vssd1 vccd1 vccd1 _15154_/Y sky130_fd_sc_hd__inv_2
X_12366_ _12366_/A vssd1 vssd1 vccd1 vccd1 _12366_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13128__B1 _13006_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14105_ _20547_/Q vssd1 vssd1 vccd1 vccd1 _17940_/A sky130_fd_sc_hd__inv_2
X_11317_ _11545_/B _11322_/A _11317_/C _11316_/X vssd1 vssd1 vccd1 vccd1 _12525_/C
+ sky130_fd_sc_hd__or4b_4
XFILLER_154_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15085_ _15085_/A _15169_/A vssd1 vssd1 vccd1 vccd1 _15086_/B sky130_fd_sc_hd__or2_2
X_19962_ _20408_/CLK _19962_/D repeater185/X vssd1 vssd1 vccd1 vccd1 _19962_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18402__S _18874_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12297_ _20513_/Q vssd1 vssd1 vccd1 vccd1 _12297_/Y sky130_fd_sc_hd__inv_2
XFILLER_141_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14036_ _14031_/A _14031_/B _14031_/C vssd1 vssd1 vccd1 vccd1 _14037_/B sky130_fd_sc_hd__o21a_1
X_18913_ _20109_/Q _21112_/Q _20871_/Q vssd1 vssd1 vccd1 vccd1 _18913_/X sky130_fd_sc_hd__mux2_1
X_11248_ _19061_/X _11244_/X _21191_/Q _11245_/X vssd1 vssd1 vccd1 vccd1 _21191_/D
+ sky130_fd_sc_hd__a22o_1
X_19893_ _21141_/CLK _19893_/D repeater192/X vssd1 vssd1 vccd1 vccd1 _19893_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_68_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18844_ _18843_/X _10755_/A _18898_/S vssd1 vssd1 vccd1 vccd1 _18844_/X sky130_fd_sc_hd__mux2_2
X_11179_ _16342_/A vssd1 vssd1 vccd1 vccd1 _11179_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_227_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18775_ _18774_/X _10578_/Y _18775_/S vssd1 vssd1 vccd1 vccd1 _18775_/X sky130_fd_sc_hd__mux2_1
XFILLER_227_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15987_ _15993_/A vssd1 vssd1 vccd1 vccd1 _15994_/A sky130_fd_sc_hd__inv_2
X_17726_ _16551_/Y _17550_/A _17725_/Y _17295_/X vssd1 vssd1 vccd1 vccd1 _17726_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_36_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14938_ _20568_/Q vssd1 vssd1 vccd1 vccd1 _14938_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20815__RESET_B repeater212/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17657_ _18739_/X _17216_/A _18710_/X _17223_/A vssd1 vssd1 vccd1 vccd1 _17657_/X
+ sky130_fd_sc_hd__o22a_2
X_14869_ _14962_/A _14991_/A vssd1 vssd1 vccd1 vccd1 _14870_/B sky130_fd_sc_hd__or2_1
XANTENNA__12686__A _12707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16608_ _16607_/Y _16605_/X _16566_/X vssd1 vssd1 vccd1 vccd1 _19990_/D sky130_fd_sc_hd__o21ai_1
XFILLER_223_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17588_ _19499_/Q vssd1 vssd1 vccd1 vccd1 _17588_/Y sky130_fd_sc_hd__inv_2
XFILLER_195_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19327_ _21234_/CLK _19327_/D vssd1 vssd1 vccd1 vccd1 _19327_/Q sky130_fd_sc_hd__dfxtp_1
X_16539_ _16539_/A vssd1 vssd1 vccd1 vccd1 _16539_/X sky130_fd_sc_hd__buf_1
XFILLER_176_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19258_ _17261_/Y _17262_/Y _17263_/Y _17264_/Y _20130_/Q _20131_/Q vssd1 vssd1 vccd1
+ vccd1 _19258_/X sky130_fd_sc_hd__mux4_2
XFILLER_148_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13367__B1 _13151_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18209_ _18208_/X _12161_/Y _18787_/S vssd1 vssd1 vccd1 vccd1 _18209_/X sky130_fd_sc_hd__mux2_2
X_19189_ _19731_/Q _19371_/Q _19787_/Q _19771_/Q _19280_/S0 _20122_/Q vssd1 vssd1
+ vccd1 vccd1 _19189_/X sky130_fd_sc_hd__mux4_1
XANTENNA__14406__A _21471_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21220_ _21222_/CLK _21220_/D repeater235/X vssd1 vssd1 vccd1 vccd1 _21220_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__13119__B1 _12993_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21151_ _21151_/CLK _21151_/D repeater223/X vssd1 vssd1 vccd1 vccd1 _21151_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18312__S _18896_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20102_ _20107_/CLK _20102_/D repeater259/X vssd1 vssd1 vccd1 vccd1 _20102_/Q sky130_fd_sc_hd__dfrtp_1
X_09913_ _21256_/Q _17023_/A _21256_/Q _17023_/A vssd1 vssd1 vccd1 vccd1 _09913_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_21082_ _21424_/CLK _21082_/D repeater230/X vssd1 vssd1 vccd1 vccd1 _21082_/Q sky130_fd_sc_hd__dfstp_2
X_20033_ _21445_/CLK _20033_/D repeater244/X vssd1 vssd1 vccd1 vccd1 _20033_/Q sky130_fd_sc_hd__dfrtp_1
X_09844_ _21439_/Q vssd1 vssd1 vccd1 vccd1 _09878_/A sky130_fd_sc_hd__inv_2
XFILLER_113_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09775_ _09775_/A _09777_/A _09781_/B vssd1 vssd1 vccd1 vccd1 _09775_/Y sky130_fd_sc_hd__nor3_1
XFILLER_227_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20935_ _20943_/CLK _20935_/D repeater277/X vssd1 vssd1 vccd1 vccd1 _20935_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_4149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20866_ _21040_/CLK _20866_/D repeater247/X vssd1 vssd1 vccd1 vccd1 _20866_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__16792__B1 _16779_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20797_ _21374_/CLK _20797_/D repeater255/X vssd1 vssd1 vccd1 vccd1 _20797_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15700__A input60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10550_ _21320_/Q vssd1 vssd1 vccd1 vccd1 _10708_/A sky130_fd_sc_hd__inv_2
XFILLER_183_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10481_ _21289_/Q vssd1 vssd1 vccd1 vccd1 _10765_/A sky130_fd_sc_hd__inv_2
XFILLER_5_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12220_ _20925_/Q vssd1 vssd1 vccd1 vccd1 _12473_/A sky130_fd_sc_hd__inv_2
X_21418_ _21419_/CLK _21418_/D repeater232/X vssd1 vssd1 vccd1 vccd1 _21418_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_204_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__21344__RESET_B repeater255/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12151_ _12307_/A _20335_/Q _12109_/X _20336_/Q vssd1 vssd1 vccd1 vccd1 _12151_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_136_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21349_ _21349_/CLK _21349_/D repeater210/X vssd1 vssd1 vccd1 vccd1 _21349_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18222__S _18236_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11102_ _11096_/B _11099_/Y _11100_/X _11101_/X _11055_/A vssd1 vssd1 vccd1 vccd1
+ _11103_/A sky130_fd_sc_hd__o32a_1
XFILLER_118_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12082_ _20967_/Q vssd1 vssd1 vccd1 vccd1 _12320_/A sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_101_HCLK clkbuf_4_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20107_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_89_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11033_ _19960_/Q _16922_/A vssd1 vssd1 vccd1 vccd1 _16926_/A sky130_fd_sc_hd__or2_1
X_15910_ _19578_/Q _15904_/X _15873_/X _15906_/X vssd1 vssd1 vccd1 vccd1 _19578_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_104_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16890_ _16892_/A _16889_/X _16971_/A vssd1 vssd1 vccd1 vccd1 _16890_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_1_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15841_ _15841_/A vssd1 vssd1 vccd1 vccd1 _15841_/X sky130_fd_sc_hd__buf_1
XFILLER_76_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19053__S _19058_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18560_ _18845_/A0 _13782_/Y _18896_/S vssd1 vssd1 vccd1 vccd1 _18560_/X sky130_fd_sc_hd__mux2_1
X_15772_ _15772_/A vssd1 vssd1 vccd1 vccd1 _15772_/X sky130_fd_sc_hd__buf_1
X_12984_ input62/X vssd1 vssd1 vccd1 vccd1 _12984_/X sky130_fd_sc_hd__buf_2
X_17511_ _19321_/Q vssd1 vssd1 vccd1 vccd1 _17511_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20297__RESET_B repeater262/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14723_ _14723_/A vssd1 vssd1 vccd1 vccd1 _14723_/X sky130_fd_sc_hd__buf_1
X_11935_ _11928_/Y _19116_/S _11934_/Y vssd1 vssd1 vccd1 vccd1 _11944_/A sky130_fd_sc_hd__o21ai_1
XANTENNA_output113_A _17091_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18892__S _18898_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18491_ _18490_/X _15133_/Y _18784_/S vssd1 vssd1 vccd1 vccd1 _18491_/X sky130_fd_sc_hd__mux2_2
XANTENNA__20226__RESET_B repeater202/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14389__A2 _20027_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17442_ _19457_/Q vssd1 vssd1 vccd1 vccd1 _17442_/Y sky130_fd_sc_hd__inv_2
X_14654_ _20172_/Q vssd1 vssd1 vccd1 vccd1 _14659_/A sky130_fd_sc_hd__buf_1
XFILLER_233_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11866_ _11860_/B _11865_/X _11803_/X _11852_/X _11804_/D vssd1 vssd1 vccd1 vccd1
+ _11867_/A sky130_fd_sc_hd__o32a_1
XFILLER_177_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13605_ _13625_/A vssd1 vssd1 vccd1 vccd1 _13605_/X sky130_fd_sc_hd__buf_1
XANTENNA__13597__B1 _13449_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10817_ _10767_/A _10767_/B _10809_/X _10815_/Y vssd1 vssd1 vccd1 vccd1 _21291_/D
+ sky130_fd_sc_hd__a211oi_2
XPHY_3982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14585_ _14585_/A _14585_/B vssd1 vssd1 vccd1 vccd1 _14616_/A sky130_fd_sc_hd__or2_1
X_17373_ _20813_/Q vssd1 vssd1 vccd1 vccd1 _17373_/Y sky130_fd_sc_hd__inv_2
XPHY_3993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17327__A2 _17324_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11797_ _12620_/A vssd1 vssd1 vccd1 vccd1 _11797_/X sky130_fd_sc_hd__buf_1
XANTENNA_repeater263_A repeater264/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19112_ _17046_/B _21071_/Q _19112_/S vssd1 vssd1 vccd1 vccd1 _19112_/X sky130_fd_sc_hd__mux2_1
X_13536_ _13572_/A vssd1 vssd1 vccd1 vccd1 _13566_/A sky130_fd_sc_hd__clkbuf_2
X_16324_ _19374_/Q _16319_/X _16016_/X _16320_/X vssd1 vssd1 vccd1 vccd1 _19374_/D
+ sky130_fd_sc_hd__a22o_1
X_10748_ _19945_/Q _19944_/Q _10748_/C _16853_/B vssd1 vssd1 vccd1 vccd1 _16868_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_185_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19043_ _16811_/X _20826_/Q _19046_/S vssd1 vssd1 vccd1 vccd1 _19933_/D sky130_fd_sc_hd__mux2_1
X_16255_ _16255_/A vssd1 vssd1 vccd1 vccd1 _16255_/X sky130_fd_sc_hd__buf_1
X_13467_ _13483_/A vssd1 vssd1 vccd1 vccd1 _13467_/X sky130_fd_sc_hd__buf_1
X_10679_ _10679_/A vssd1 vssd1 vccd1 vccd1 _10679_/Y sky130_fd_sc_hd__inv_2
XFILLER_145_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15206_ _20051_/Q _15205_/Y _15177_/A _15067_/B vssd1 vssd1 vccd1 vccd1 _20051_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_127_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12418_ _12469_/B _12418_/B vssd1 vssd1 vccd1 vccd1 _12419_/B sky130_fd_sc_hd__or2_2
X_16186_ _19442_/Q _16180_/X _16139_/X _16182_/X vssd1 vssd1 vccd1 vccd1 _19442_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_154_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13398_ _13410_/A vssd1 vssd1 vccd1 vccd1 _13398_/X sky130_fd_sc_hd__buf_1
XANTENNA__12572__A1 _13188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12572__B2 _18242_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15137_ _20458_/Q vssd1 vssd1 vccd1 vccd1 _15137_/Y sky130_fd_sc_hd__inv_2
XFILLER_245_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12349_ _12364_/A vssd1 vssd1 vccd1 vccd1 _12350_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__18132__S _18669_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21014__RESET_B repeater238/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15068_ _15068_/A _15068_/B _15202_/A vssd1 vssd1 vccd1 vccd1 _15198_/A sky130_fd_sc_hd__or3_1
X_19945_ _21372_/CLK _19945_/D repeater251/X vssd1 vssd1 vccd1 vccd1 _19945_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_68_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14019_ _14017_/A _14017_/B _14017_/Y _14004_/X vssd1 vssd1 vccd1 vccd1 _20301_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_110_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19876_ _21421_/CLK _19876_/D repeater214/X vssd1 vssd1 vccd1 vccd1 _19876_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__19374__CLK _19706_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18827_ _18826_/X _09740_/Y _18928_/S vssd1 vssd1 vccd1 vccd1 _18827_/X sky130_fd_sc_hd__mux2_1
XFILLER_209_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18758_ _18757_/X _17531_/Y _18927_/S vssd1 vssd1 vccd1 vccd1 _18758_/X sky130_fd_sc_hd__mux2_1
XFILLER_243_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17709_ _20817_/Q vssd1 vssd1 vccd1 vccd1 _17709_/Y sky130_fd_sc_hd__inv_2
X_18689_ _18845_/A0 _13824_/Y _18896_/S vssd1 vssd1 vccd1 vccd1 _18689_/X sky130_fd_sc_hd__mux2_1
XANTENNA__17566__A2 _17639_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20720_ _20724_/CLK _20720_/D repeater264/X vssd1 vssd1 vccd1 vccd1 _20720_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_63_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20651_ _20657_/CLK _20651_/D repeater197/X vssd1 vssd1 vccd1 vccd1 _20651_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__16616__A _16616_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18307__S _18644_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17318__A2 _17861_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20582_ _20946_/CLK _20582_/D repeater274/X vssd1 vssd1 vccd1 vccd1 _20582_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_139_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13040__A _13040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_124_HCLK clkbuf_4_4_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20957_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_219_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21203_ _21255_/CLK _21203_/D repeater240/X vssd1 vssd1 vccd1 vccd1 _21203_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_155_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21134_ _21134_/CLK _21134_/D repeater192/X vssd1 vssd1 vccd1 vccd1 _21134_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_105_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13512__B1 _13511_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21065_ _21087_/CLK _21065_/D repeater228/X vssd1 vssd1 vccd1 vccd1 _21065_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_171_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20016_ _21424_/CLK _20016_/D repeater230/X vssd1 vssd1 vccd1 vccd1 _20016_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__20737__RESET_B repeater211/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09827_ _09827_/A vssd1 vssd1 vccd1 vccd1 _09827_/X sky130_fd_sc_hd__buf_1
XFILLER_47_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09758_ _21228_/Q vssd1 vssd1 vccd1 vccd1 _11053_/A sky130_fd_sc_hd__inv_2
XFILLER_234_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20390__RESET_B repeater278/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09689_ _21466_/Q _09673_/X _09688_/X _09678_/X vssd1 vssd1 vccd1 vccd1 _21466_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17557__A2 _17639_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18754__A1 _20502_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11720_ _11720_/A vssd1 vssd1 vccd1 vccd1 _11720_/X sky130_fd_sc_hd__buf_1
XPHY_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20918_ _20949_/CLK _20918_/D repeater269/X vssd1 vssd1 vccd1 vccd1 _20918_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17962__C1 _17961_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13579__B1 _13426_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11651_ _21408_/Q _11617_/A _21422_/Q _21096_/Q _11642_/X vssd1 vssd1 vccd1 vccd1
+ _21096_/D sky130_fd_sc_hd__a32o_1
XPHY_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20849_ _20857_/CLK _20849_/D repeater244/X vssd1 vssd1 vccd1 vccd1 _20849_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18217__S _18242_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10602_ _20761_/Q vssd1 vssd1 vccd1 vccd1 _10602_/Y sky130_fd_sc_hd__inv_2
XPHY_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14370_ _14461_/A _14370_/B vssd1 vssd1 vccd1 vccd1 _14483_/A sky130_fd_sc_hd__or2_1
XPHY_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11582_ _11590_/A vssd1 vssd1 vccd1 vccd1 _11583_/B sky130_fd_sc_hd__buf_1
XPHY_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13321_ _13321_/A vssd1 vssd1 vccd1 vccd1 _13321_/X sky130_fd_sc_hd__buf_1
X_10533_ _21337_/Q vssd1 vssd1 vccd1 vccd1 _10534_/B sky130_fd_sc_hd__inv_2
XFILLER_7_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16040_ _19515_/Q _16035_/X _15975_/X _16037_/X vssd1 vssd1 vccd1 vccd1 _19515_/D
+ sky130_fd_sc_hd__a22o_1
X_13252_ _20566_/Q _13248_/X _13171_/X _13249_/X vssd1 vssd1 vccd1 vccd1 _20566_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_input74_A RsRx_S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10464_ _21277_/Q _10459_/Y _10772_/A _20685_/Q _10463_/X vssd1 vssd1 vccd1 vccd1
+ _10471_/C sky130_fd_sc_hd__o221a_1
XFILLER_170_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12203_ _12331_/A _20360_/Q _20956_/Q _12150_/Y _12202_/X vssd1 vssd1 vccd1 vccd1
+ _12204_/D sky130_fd_sc_hd__o221a_1
XANTENNA__19048__S _19058_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13183_ _18975_/S _13178_/X _18972_/X _13521_/A _13182_/X vssd1 vssd1 vccd1 vccd1
+ _13184_/S sky130_fd_sc_hd__a2111o_2
X_10395_ _10395_/A vssd1 vssd1 vccd1 vccd1 _10395_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_123_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12134_ _20972_/Q vssd1 vssd1 vccd1 vccd1 _12325_/A sky130_fd_sc_hd__inv_2
X_17991_ _20832_/Q vssd1 vssd1 vccd1 vccd1 _17991_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18887__S _18899_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13503__B1 _13311_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19730_ _19789_/CLK _19730_/D vssd1 vssd1 vccd1 vccd1 _19730_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12065_ _12310_/A _20370_/Q _12064_/Y _20395_/Q vssd1 vssd1 vccd1 vccd1 _12065_/X
+ sky130_fd_sc_hd__o22a_1
X_16942_ _19964_/Q _16937_/A _16941_/Y _16937_/Y vssd1 vssd1 vccd1 vccd1 _16943_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_77_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18442__A0 _17079_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11016_ _09919_/B _11584_/C _21244_/Q vssd1 vssd1 vccd1 vccd1 _11017_/B sky130_fd_sc_hd__o21a_1
X_19661_ _19821_/CLK _19661_/D vssd1 vssd1 vccd1 vccd1 _19661_/Q sky130_fd_sc_hd__dfxtp_1
X_16873_ _19946_/Q _16868_/A _19947_/Q vssd1 vssd1 vccd1 vccd1 _16873_/X sky130_fd_sc_hd__o21a_1
XFILLER_93_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18612_ _18611_/X _16921_/Y _18680_/S vssd1 vssd1 vccd1 vccd1 _18612_/X sky130_fd_sc_hd__mux2_2
XANTENNA__20407__RESET_B repeater184/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15824_ _15824_/A vssd1 vssd1 vccd1 vccd1 _15824_/X sky130_fd_sc_hd__buf_1
X_19592_ _20890_/CLK _19592_/D vssd1 vssd1 vccd1 vccd1 _19592_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18543_ _17830_/X _09756_/Y _18928_/S vssd1 vssd1 vccd1 vccd1 _18543_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15755_ _19646_/Q _15750_/X _15706_/X _15751_/X vssd1 vssd1 vccd1 vccd1 _19646_/D
+ sky130_fd_sc_hd__a22o_1
X_12967_ _20806_/Q _20805_/Q _20807_/Q _12966_/X vssd1 vssd1 vccd1 vccd1 _12968_/C
+ sky130_fd_sc_hd__a31o_1
XANTENNA__18745__A1 _20742_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20060__RESET_B repeater281/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14706_ _14724_/A vssd1 vssd1 vccd1 vccd1 _14706_/X sky130_fd_sc_hd__buf_1
X_11918_ _19117_/X vssd1 vssd1 vccd1 vccd1 _11943_/A sky130_fd_sc_hd__inv_2
X_18474_ _18473_/X _14577_/A _18898_/S vssd1 vssd1 vccd1 vccd1 _18474_/X sky130_fd_sc_hd__mux2_2
XFILLER_178_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15686_ _19678_/Q _15681_/X _15592_/X _15682_/X vssd1 vssd1 vccd1 vccd1 _19678_/D
+ sky130_fd_sc_hd__a22o_1
X_12898_ _12898_/A _12898_/B vssd1 vssd1 vccd1 vccd1 _13261_/A sky130_fd_sc_hd__or2_4
XPHY_4480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17425_ _17425_/A vssd1 vssd1 vccd1 vccd1 _17425_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_220_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14637_ _14637_/A vssd1 vssd1 vccd1 vccd1 _14637_/Y sky130_fd_sc_hd__inv_2
X_11849_ _11845_/B _11816_/Y _11848_/X _11817_/X _11848_/A vssd1 vssd1 vccd1 vccd1
+ _21031_/D sky130_fd_sc_hd__a32o_1
XANTENNA__18127__S _18850_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14568_ _14568_/A _14568_/B vssd1 vssd1 vccd1 vccd1 _14648_/A sky130_fd_sc_hd__or2_1
XFILLER_147_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17356_ _19592_/Q vssd1 vssd1 vccd1 vccd1 _17356_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_147_HCLK clkbuf_opt_1_HCLK/A vssd1 vssd1 vccd1 vccd1 _20136_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_174_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16307_ _19385_/Q _16305_/X _16288_/X _16306_/X vssd1 vssd1 vccd1 vccd1 _19385_/D
+ sky130_fd_sc_hd__a22o_1
X_13519_ _20433_/Q _13514_/X _13454_/X _13515_/X vssd1 vssd1 vccd1 vccd1 _20433_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_119_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14499_ _14499_/A _14513_/A vssd1 vssd1 vccd1 vccd1 _14500_/B sky130_fd_sc_hd__or2_1
XANTENNA__10484__A _20692_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17287_ _21057_/Q vssd1 vssd1 vccd1 vccd1 _17287_/Y sky130_fd_sc_hd__inv_2
XFILLER_158_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19026_ _16884_/Y _20397_/Q _19026_/S vssd1 vssd1 vccd1 vccd1 _19950_/D sky130_fd_sc_hd__mux2_1
X_16238_ _19419_/Q _16230_/X _16237_/X _16233_/X vssd1 vssd1 vccd1 vccd1 _19419_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_173_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16169_ _19453_/Q _16166_/X _16131_/X _16168_/X vssd1 vssd1 vccd1 vccd1 _19453_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_114_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18681__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18797__S _18927_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15495__B1 _15450_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19928_ _21207_/CLK _19928_/D repeater256/X vssd1 vssd1 vccd1 vccd1 _19928_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_130_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20830__RESET_B repeater251/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19859_ _21164_/CLK _19859_/D repeater226/X vssd1 vssd1 vccd1 vccd1 _19859_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_110_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09612_ _20886_/Q _20885_/Q _20876_/Q vssd1 vssd1 vccd1 vccd1 _12716_/B sky130_fd_sc_hd__or3_4
XANTENNA__20148__RESET_B repeater250/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13035__A _13041_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10087__A2 _10086_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20703_ _21349_/CLK _20703_/D repeater210/X vssd1 vssd1 vccd1 vccd1 _20703_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_169_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20255__SET_B repeater217/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20634_ _21486_/CLK _20634_/D repeater198/X vssd1 vssd1 vccd1 vccd1 _20634_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_149_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20565_ _20592_/CLK _20565_/D repeater260/X vssd1 vssd1 vccd1 vccd1 _20565_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_166_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20496_ _20496_/CLK _20496_/D repeater273/X vssd1 vssd1 vccd1 vccd1 _20496_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_152_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17177__A _17177_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10180_ _21399_/Q _10179_/Y _10170_/X _10161_/B vssd1 vssd1 vccd1 vccd1 _21399_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_132_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21117_ _21120_/CLK _21117_/D repeater233/X vssd1 vssd1 vccd1 vccd1 _21117_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_132_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18500__S _18666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21048_ _21087_/CLK _21048_/D repeater227/X vssd1 vssd1 vccd1 vccd1 _21048_/Q sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_28_HCLK clkbuf_4_9_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _21424_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_59_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13870_ _14014_/A _14013_/A _14012_/A _14009_/A vssd1 vssd1 vccd1 vccd1 _13877_/C
+ sky130_fd_sc_hd__or4_4
X_12821_ _12841_/A vssd1 vssd1 vccd1 vccd1 _12821_/X sky130_fd_sc_hd__buf_1
XFILLER_234_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15540_ _19751_/Q _15536_/X _15524_/X _15537_/X vssd1 vssd1 vccd1 vccd1 _19751_/D
+ sky130_fd_sc_hd__a22o_1
X_12752_ _20805_/Q _12751_/Y _12748_/X vssd1 vssd1 vccd1 vccd1 _20805_/D sky130_fd_sc_hd__o21a_1
XPHY_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11703_ _21076_/Q _11697_/X _11560_/X _11699_/X vssd1 vssd1 vccd1 vccd1 _21076_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15471_ _15481_/A vssd1 vssd1 vccd1 vccd1 _15471_/X sky130_fd_sc_hd__buf_1
XFILLER_202_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12683_ _20828_/Q _12679_/X _09636_/X _12680_/X vssd1 vssd1 vccd1 vccd1 _20828_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_199_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15410__B1 _15355_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14422_ _21467_/Q _14498_/A _21480_/Q _14461_/B vssd1 vssd1 vccd1 vccd1 _14422_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17210_ _17889_/A vssd1 vssd1 vccd1 vccd1 _17211_/A sky130_fd_sc_hd__buf_1
XPHY_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11634_ _11632_/A _11632_/B _11617_/X _11632_/Y vssd1 vssd1 vccd1 vccd1 _21105_/D
+ sky130_fd_sc_hd__a211oi_2
XPHY_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18190_ _18189_/X _14385_/Y _18669_/S vssd1 vssd1 vccd1 vccd1 _18190_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14353_ _20215_/Q vssd1 vssd1 vccd1 vccd1 _14500_/A sky130_fd_sc_hd__inv_2
X_17141_ _17141_/A vssd1 vssd1 vccd1 vccd1 _17142_/A sky130_fd_sc_hd__buf_1
XPHY_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11565_ _13166_/A vssd1 vssd1 vccd1 vccd1 _11565_/X sky130_fd_sc_hd__clkbuf_2
XPHY_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13304_ _20544_/Q _13300_/X _13144_/X _13302_/X vssd1 vssd1 vccd1 vccd1 _20544_/D
+ sky130_fd_sc_hd__a22o_1
X_17072_ _17076_/C _17072_/B _19889_/Q vssd1 vssd1 vccd1 vccd1 _19884_/D sky130_fd_sc_hd__and3_1
XFILLER_183_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10516_ _21278_/Q vssd1 vssd1 vccd1 vccd1 _10755_/A sky130_fd_sc_hd__inv_2
XFILLER_183_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14284_ _20123_/Q _14280_/X _16451_/A _15919_/A _14783_/B vssd1 vssd1 vccd1 vccd1
+ _14284_/X sky130_fd_sc_hd__a32o_1
X_11496_ _11511_/B vssd1 vssd1 vccd1 vccd1 _11497_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__12008__B _19908_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13235_ _20576_/Q _13233_/X _13151_/X _13234_/X vssd1 vssd1 vccd1 vccd1 _20576_/D
+ sky130_fd_sc_hd__a22o_1
X_16023_ _16029_/A vssd1 vssd1 vccd1 vccd1 _16023_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_109_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10447_ _20668_/Q vssd1 vssd1 vccd1 vccd1 _10447_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13166_ _13166_/A vssd1 vssd1 vccd1 vccd1 _13166_/X sky130_fd_sc_hd__clkbuf_4
X_10378_ _21369_/Q _10377_/Y _10373_/X _10285_/B vssd1 vssd1 vccd1 vccd1 _21369_/D
+ sky130_fd_sc_hd__o211a_1
X_12117_ _12314_/A _20375_/Q _20964_/Q _17895_/A _12116_/X vssd1 vssd1 vccd1 vccd1
+ _12145_/C sky130_fd_sc_hd__o221a_1
XFILLER_112_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18410__S _18748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13097_ _20638_/Q _13092_/X _12872_/X _13093_/X vssd1 vssd1 vccd1 vccd1 _20638_/D
+ sky130_fd_sc_hd__a22o_1
X_17974_ _17974_/A vssd1 vssd1 vccd1 vccd1 _17978_/B sky130_fd_sc_hd__buf_4
X_19713_ _19776_/CLK _19713_/D vssd1 vssd1 vccd1 vccd1 _19713_/Q sky130_fd_sc_hd__dfxtp_1
X_12048_ _20387_/Q vssd1 vssd1 vccd1 vccd1 _12048_/Y sky130_fd_sc_hd__inv_2
X_16925_ _19960_/Q vssd1 vssd1 vccd1 vccd1 _16927_/A sky130_fd_sc_hd__inv_2
XFILLER_238_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20241__RESET_B repeater248/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19644_ _20327_/CLK _19644_/D vssd1 vssd1 vccd1 vccd1 _19644_/Q sky130_fd_sc_hd__dfxtp_1
X_16856_ _19943_/Q _16856_/B vssd1 vssd1 vccd1 vccd1 _16861_/B sky130_fd_sc_hd__or2_1
XFILLER_226_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15807_ _15807_/A vssd1 vssd1 vccd1 vccd1 _15807_/X sky130_fd_sc_hd__buf_1
X_19575_ _19961_/CLK _19575_/D vssd1 vssd1 vccd1 vccd1 _19575_/Q sky130_fd_sc_hd__dfxtp_1
X_16787_ _19926_/Q _16777_/A _19927_/Q vssd1 vssd1 vccd1 vccd1 _16787_/X sky130_fd_sc_hd__o21a_1
X_13999_ _13999_/A vssd1 vssd1 vccd1 vccd1 _13999_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18526_ _18525_/X _15096_/Y _18906_/S vssd1 vssd1 vccd1 vccd1 _18526_/X sky130_fd_sc_hd__mux2_1
XFILLER_234_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15738_ _19657_/Q _15736_/X _15697_/X _15737_/X vssd1 vssd1 vccd1 vccd1 _19657_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_222_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21447__RESET_B repeater248/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18457_ _17830_/X _09727_/Y _18928_/S vssd1 vssd1 vccd1 vccd1 _18457_/X sky130_fd_sc_hd__mux2_1
X_15669_ _19688_/Q _15666_/X _15588_/X _15667_/X vssd1 vssd1 vccd1 vccd1 _19688_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12694__A _12708_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_221_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17408_ _19641_/Q vssd1 vssd1 vccd1 vccd1 _17408_/Y sky130_fd_sc_hd__inv_2
X_18388_ _18387_/X _15123_/Y _18906_/S vssd1 vssd1 vccd1 vccd1 _18388_/X sky130_fd_sc_hd__mux2_2
XFILLER_187_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17339_ _19384_/Q vssd1 vssd1 vccd1 vccd1 _17339_/Y sky130_fd_sc_hd__inv_2
X_20350_ _20480_/CLK _20350_/D repeater183/X vssd1 vssd1 vccd1 vccd1 _20350_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_147_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19009_ _16956_/Y _20414_/Q _19019_/S vssd1 vssd1 vccd1 vccd1 _19967_/D sky130_fd_sc_hd__mux2_1
XANTENNA__13715__B1 _13714_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20281_ _20293_/CLK _20281_/D repeater263/X vssd1 vssd1 vccd1 vccd1 _20281_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_127_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18654__A0 _17079_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20329__RESET_B repeater190/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18320__S _18909_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18406__A0 _17079_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_124_HCLK_A clkbuf_4_4_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__21117__RESET_B repeater233/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_212_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19134__A1 _19375_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20617_ _20622_/CLK _20617_/D repeater194/X vssd1 vssd1 vccd1 vccd1 _20617_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_177_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11350_ _11350_/A _11366_/C vssd1 vssd1 vccd1 vccd1 _11390_/D sky130_fd_sc_hd__or2_1
XFILLER_20_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20548_ _20947_/CLK _20548_/D repeater266/X vssd1 vssd1 vccd1 vccd1 _20548_/Q sky130_fd_sc_hd__dfrtp_4
X_10301_ _21373_/Q _18083_/A _10283_/A _20727_/Q vssd1 vssd1 vccd1 vccd1 _10301_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_180_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11281_ _20907_/Q vssd1 vssd1 vccd1 vccd1 _11310_/C sky130_fd_sc_hd__buf_1
XFILLER_152_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20479_ _20480_/CLK _20479_/D repeater183/X vssd1 vssd1 vccd1 vccd1 _20479_/Q sky130_fd_sc_hd__dfrtp_1
X_13020_ _13020_/A vssd1 vssd1 vccd1 vccd1 _13041_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_4_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10232_ _21371_/Q vssd1 vssd1 vccd1 vccd1 _10286_/A sky130_fd_sc_hd__inv_2
XFILLER_105_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10163_ _10163_/A _10172_/A vssd1 vssd1 vccd1 vccd1 _10164_/A sky130_fd_sc_hd__or2_2
XANTENNA__18230__S _18236_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input37_A HTRANS[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14971_ _14880_/A _14880_/B _14970_/X _14968_/Y vssd1 vssd1 vccd1 vccd1 _20102_/D
+ sky130_fd_sc_hd__a211oi_2
X_10094_ _20783_/Q vssd1 vssd1 vccd1 vccd1 _10094_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18948__A1 _21088_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16710_ _19899_/Q _14239_/B _14240_/B vssd1 vssd1 vccd1 vccd1 _16710_/X sky130_fd_sc_hd__a21bo_1
X_13922_ _13922_/A _13922_/B _13922_/C _13921_/X vssd1 vssd1 vccd1 vccd1 _13922_/X
+ sky130_fd_sc_hd__or4b_1
X_17690_ _19628_/Q vssd1 vssd1 vccd1 vccd1 _17690_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16641_ _16643_/A _18959_/X vssd1 vssd1 vccd1 vccd1 _19855_/D sky130_fd_sc_hd__and2_1
XFILLER_90_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13853_ _20308_/Q vssd1 vssd1 vccd1 vccd1 _13884_/A sky130_fd_sc_hd__inv_2
XFILLER_62_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19061__S _19910_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_216_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19360_ _19521_/CLK _19360_/D vssd1 vssd1 vccd1 vccd1 _19360_/Q sky130_fd_sc_hd__dfxtp_1
X_12804_ _12804_/A vssd1 vssd1 vccd1 vccd1 _12804_/X sky130_fd_sc_hd__buf_1
X_16572_ _20002_/Q _19999_/Q _19998_/Q _16621_/A vssd1 vssd1 vccd1 vccd1 _16573_/A
+ sky130_fd_sc_hd__or4_4
XANTENNA_clkbuf_leaf_46_HCLK_A _20004_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13784_ _13782_/Y _20186_/Q _17978_/A _20196_/Q vssd1 vssd1 vccd1 vccd1 _13784_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_43_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10996_ _10988_/X _10992_/X _10993_/Y _10994_/X _11896_/B vssd1 vssd1 vccd1 vccd1
+ _10996_/X sky130_fd_sc_hd__a32o_1
XFILLER_204_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18311_ _18310_/X _14588_/A _18748_/S vssd1 vssd1 vccd1 vccd1 _18311_/X sky130_fd_sc_hd__mux2_1
XFILLER_35_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15523_ _15523_/A vssd1 vssd1 vccd1 vccd1 _15793_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_15_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19291_ _20075_/CLK hold9/X vssd1 vssd1 vccd1 vccd1 _19291_/Q sky130_fd_sc_hd__dfxtp_1
X_12735_ _12735_/A vssd1 vssd1 vccd1 vccd1 _16526_/A sky130_fd_sc_hd__inv_2
XFILLER_203_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_repeater176_A _18644_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18242_ _20866_/Q input16/X _18242_/S vssd1 vssd1 vccd1 vccd1 _18242_/X sky130_fd_sc_hd__mux2_1
XPHY_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15454_ _15661_/A vssd1 vssd1 vccd1 vccd1 _15454_/X sky130_fd_sc_hd__clkbuf_2
X_12666_ input56/X vssd1 vssd1 vccd1 vccd1 _12666_/X sky130_fd_sc_hd__buf_2
XFILLER_31_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19125__A1 _14313_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14405_ _14402_/Y _20222_/Q _21476_/Q _14460_/C _14404_/X vssd1 vssd1 vccd1 vccd1
+ _14420_/A sky130_fd_sc_hd__o221a_1
XFILLER_169_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11617_ _11617_/A vssd1 vssd1 vccd1 vccd1 _11617_/X sky130_fd_sc_hd__clkbuf_2
XPHY_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18173_ _18172_/X _16878_/Y _18886_/S vssd1 vssd1 vccd1 vccd1 _18173_/X sky130_fd_sc_hd__mux2_1
XPHY_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12597_ _20875_/Q _12594_/X _18227_/X _12595_/X vssd1 vssd1 vccd1 vccd1 _20875_/D
+ sky130_fd_sc_hd__a22o_1
X_15385_ _15385_/A vssd1 vssd1 vccd1 vccd1 _15663_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__16714__A _16718_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19220__S1 _20131_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18405__S _18907_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17124_ _19614_/Q vssd1 vssd1 vccd1 vccd1 _17124_/Y sky130_fd_sc_hd__inv_2
XPHY_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11548_ _21135_/Q _11547_/X _19119_/X vssd1 vssd1 vccd1 vccd1 _21135_/D sky130_fd_sc_hd__mux2_1
X_14336_ _14336_/A vssd1 vssd1 vccd1 vccd1 _14460_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_237_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17055_ _17058_/C _17055_/B _19851_/Q vssd1 vssd1 vccd1 vccd1 _19847_/D sky130_fd_sc_hd__nor3_1
XFILLER_171_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14267_ _14267_/A vssd1 vssd1 vccd1 vccd1 _14267_/X sky130_fd_sc_hd__buf_1
X_11479_ _19102_/X _11474_/X _21156_/Q _11475_/X vssd1 vssd1 vccd1 vccd1 _21156_/D
+ sky130_fd_sc_hd__a22o_1
X_16006_ _16332_/A vssd1 vssd1 vccd1 vccd1 _16006_/X sky130_fd_sc_hd__buf_2
X_13218_ _20584_/Q _13215_/X _13216_/X _13217_/X vssd1 vssd1 vccd1 vccd1 _20584_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_171_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14198_ _14198_/A vssd1 vssd1 vccd1 vccd1 _14198_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13149_ _20611_/Q _13139_/X _13148_/X _13142_/X vssd1 vssd1 vccd1 vccd1 _20611_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18140__S _18897_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17957_ _17957_/A _17957_/B _17957_/C _17957_/D vssd1 vssd1 vccd1 vccd1 _17957_/X
+ sky130_fd_sc_hd__or4_4
XFILLER_66_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18939__A1 _21137_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16908_ _19956_/Q vssd1 vssd1 vccd1 vccd1 _16910_/A sky130_fd_sc_hd__inv_2
XANTENNA__12684__B1 _09638_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17888_ _18422_/X _17200_/X _18415_/X _17224_/X _17887_/X vssd1 vssd1 vccd1 vccd1
+ _17888_/X sky130_fd_sc_hd__o221a_1
X_19627_ _21040_/CLK _19627_/D vssd1 vssd1 vccd1 vccd1 _19627_/Q sky130_fd_sc_hd__dfxtp_1
X_16839_ _19939_/Q vssd1 vssd1 vccd1 vccd1 _16839_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19558_ _19706_/CLK _19558_/D vssd1 vssd1 vccd1 vccd1 _19558_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__21281__RESET_B repeater211/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18509_ _18508_/X _14395_/Y _18897_/S vssd1 vssd1 vccd1 vccd1 _18509_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19489_ _21449_/CLK _19489_/D vssd1 vssd1 vccd1 vccd1 _19489_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19116__A1 _11916_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21451_ _21452_/CLK _21451_/D repeater247/X vssd1 vssd1 vccd1 vccd1 _21451_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__19211__S1 _20133_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18315__S _18906_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20402_ _20809_/CLK _20402_/D repeater188/X vssd1 vssd1 vccd1 vccd1 _20402_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_31_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21382_ _21390_/CLK _21382_/D repeater214/X vssd1 vssd1 vccd1 vccd1 _21382_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_147_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20333_ _20809_/CLK _20333_/D repeater270/X vssd1 vssd1 vccd1 vccd1 _20333_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_190_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13164__A1 _20603_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20264_ _21366_/CLK _20264_/D repeater265/X vssd1 vssd1 vccd1 vccd1 _20264_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_115_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17455__A _21059_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20195_ _20626_/CLK _20195_/D repeater193/X vssd1 vssd1 vccd1 vccd1 _20195_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_248_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17174__B _17174_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19278__S1 _20122_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15861__B1 _15795_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12675__B1 _12673_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__21369__RESET_B repeater254/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17902__B _17944_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10850_ _18281_/X _10847_/X _21275_/Q _10849_/X vssd1 vssd1 vccd1 vccd1 _21275_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_71_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09701__A _15354_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10781_ _10781_/A _10781_/B vssd1 vssd1 vccd1 vccd1 _10790_/A sky130_fd_sc_hd__or2_1
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12520_ _12520_/A vssd1 vssd1 vccd1 vccd1 _12520_/X sky130_fd_sc_hd__buf_1
XANTENNA__13223__A input45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_234_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19107__A1 _14313_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12451_ _12451_/A vssd1 vssd1 vccd1 vccd1 _12451_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18225__S _18236_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19202__S1 _21004_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11402_ _16507_/A _11402_/B vssd1 vssd1 vccd1 vccd1 _11403_/A sky130_fd_sc_hd__or2_2
XFILLER_172_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15170_ _20071_/Q _15169_/Y _15166_/X _15086_/B vssd1 vssd1 vccd1 vccd1 _20071_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_138_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12382_ _12310_/A _12310_/B _12350_/A _12380_/Y vssd1 vssd1 vccd1 vccd1 _20956_/D
+ sky130_fd_sc_hd__a211oi_2
X_14121_ _20532_/Q vssd1 vssd1 vccd1 vccd1 _14121_/Y sky130_fd_sc_hd__inv_2
X_11333_ _21175_/Q _21174_/Q _11367_/B vssd1 vssd1 vccd1 vccd1 _11350_/A sky130_fd_sc_hd__or3_1
XFILLER_165_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13155__A1 _20609_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14052_ _20276_/Q vssd1 vssd1 vccd1 vccd1 _14086_/A sky130_fd_sc_hd__inv_2
XFILLER_113_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11264_ _20914_/Q vssd1 vssd1 vccd1 vccd1 _11541_/A sky130_fd_sc_hd__buf_1
XFILLER_140_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13003_ input54/X vssd1 vssd1 vccd1 vccd1 _13003_/X sky130_fd_sc_hd__buf_2
XFILLER_137_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19056__S _19058_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10215_ _10203_/A _10203_/B _10213_/Y _10177_/X vssd1 vssd1 vccd1 vccd1 _21382_/D
+ sky130_fd_sc_hd__a211oi_2
X_18860_ _18859_/X _21247_/Q _20869_/Q vssd1 vssd1 vccd1 vccd1 _18860_/X sky130_fd_sc_hd__mux2_1
X_11195_ _21216_/Q _11191_/X _10894_/X _11193_/X vssd1 vssd1 vccd1 vccd1 _21216_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_239_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17811_ _17811_/A _17812_/B vssd1 vssd1 vccd1 vccd1 _17811_/Y sky130_fd_sc_hd__nor2_1
XFILLER_79_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10146_ _10077_/C _10168_/B _10077_/A vssd1 vssd1 vccd1 vccd1 _10147_/C sky130_fd_sc_hd__o21a_1
X_18791_ _17447_/Y _17446_/X _18926_/S vssd1 vssd1 vccd1 vccd1 _18791_/X sky130_fd_sc_hd__mux2_1
XANTENNA__18895__S _18901_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19269__S1 _20131_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17742_ _19365_/Q vssd1 vssd1 vccd1 vccd1 _17742_/Y sky130_fd_sc_hd__inv_2
X_14954_ _14954_/A vssd1 vssd1 vccd1 vccd1 _14989_/A sky130_fd_sc_hd__buf_1
X_10077_ _10077_/A _10220_/A _10077_/C vssd1 vssd1 vccd1 vccd1 _10078_/A sky130_fd_sc_hd__or3_1
XFILLER_94_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_235_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20928__CLK _20930_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13905_ _13904_/Y _20322_/Q _20665_/Q _13899_/Y vssd1 vssd1 vccd1 vccd1 _13905_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_235_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17812__B _17812_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17673_ _19412_/Q vssd1 vssd1 vccd1 vccd1 _17673_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14885_ _20107_/Q vssd1 vssd1 vccd1 vccd1 _14885_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14407__B2 _20025_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21039__RESET_B repeater242/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19412_ _21001_/CLK _19412_/D vssd1 vssd1 vccd1 vccd1 _19412_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_235_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16624_ _16624_/A vssd1 vssd1 vccd1 vccd1 _16624_/Y sky130_fd_sc_hd__inv_2
XFILLER_47_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13836_ _13836_/A _13836_/B _13836_/C _13836_/D vssd1 vssd1 vccd1 vccd1 _13837_/D
+ sky130_fd_sc_hd__and4_1
XANTENNA_clkbuf_leaf_170_HCLK_A clkbuf_opt_2_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19343_ _19961_/CLK _19343_/D vssd1 vssd1 vccd1 vccd1 _19343_/Q sky130_fd_sc_hd__dfxtp_1
X_16555_ _19996_/Q vssd1 vssd1 vccd1 vccd1 _16556_/B sky130_fd_sc_hd__inv_2
X_13767_ _20601_/Q _14568_/A _13763_/Y _20178_/Q _13766_/X vssd1 vssd1 vccd1 vccd1
+ _13767_/X sky130_fd_sc_hd__a221o_1
XFILLER_50_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10979_ _20999_/Q _11190_/A _11153_/A vssd1 vssd1 vccd1 vccd1 _15505_/C sky130_fd_sc_hd__or3_4
XFILLER_90_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13091__B1 _13032_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15506_ _15528_/A _15542_/B _15722_/C vssd1 vssd1 vccd1 vccd1 _15516_/A sky130_fd_sc_hd__or3_4
XFILLER_231_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10444__A2 _20695_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12718_ _11179_/X _20810_/Q _12718_/S vssd1 vssd1 vccd1 vccd1 _20810_/D sky130_fd_sc_hd__mux2_1
X_19274_ _17101_/Y _17102_/Y _17103_/Y _17104_/Y _19275_/S0 _21004_/Q vssd1 vssd1
+ vccd1 vccd1 _19274_/X sky130_fd_sc_hd__mux4_2
X_16486_ _17684_/A vssd1 vssd1 vccd1 vccd1 _18929_/S sky130_fd_sc_hd__clkinv_8
X_13698_ _20340_/Q _13693_/X _13586_/X _13694_/X vssd1 vssd1 vccd1 vccd1 _20340_/D
+ sky130_fd_sc_hd__a22o_1
X_18225_ _20849_/Q input29/X _18236_/S vssd1 vssd1 vccd1 vccd1 _18225_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13918__B1 _13917_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15437_ _19797_/Q _15434_/X _15378_/X _15436_/X vssd1 vssd1 vccd1 vccd1 _19797_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_248_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12649_ _12685_/A vssd1 vssd1 vccd1 vccd1 _12679_/A sky130_fd_sc_hd__buf_1
XANTENNA__18135__S _18667_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20674__RESET_B repeater208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18156_ _18155_/X _10774_/A _18617_/S vssd1 vssd1 vccd1 vccd1 _18156_/X sky130_fd_sc_hd__mux2_1
X_15368_ _19825_/Q _15366_/X _15346_/X _15367_/X vssd1 vssd1 vccd1 vccd1 _19825_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_7_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17107_ _19292_/Q vssd1 vssd1 vccd1 vccd1 _17107_/Y sky130_fd_sc_hd__inv_2
X_14319_ _14292_/X _14315_/Y _14318_/X vssd1 vssd1 vccd1 vccd1 _14319_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_116_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18087_ _18617_/X _17907_/A _18627_/X _17908_/A vssd1 vssd1 vccd1 vccd1 _18090_/B
+ sky130_fd_sc_hd__a22o_1
X_15299_ _19865_/Q _15299_/B vssd1 vssd1 vccd1 vccd1 _15302_/A sky130_fd_sc_hd__or2_2
XFILLER_172_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17038_ _17038_/A _17038_/B vssd1 vssd1 vccd1 vccd1 _20022_/D sky130_fd_sc_hd__nor2_1
XFILLER_113_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21245__SET_B repeater238/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19905__D _19905_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09860_ _20034_/Q vssd1 vssd1 vccd1 vccd1 _10842_/A sky130_fd_sc_hd__inv_2
XANTENNA__19750__CLK _21009_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09791_ _16619_/B _09789_/Y _16619_/A _09788_/X vssd1 vssd1 vccd1 vccd1 _21458_/D
+ sky130_fd_sc_hd__o22ai_1
X_18989_ _21264_/Q _21116_/Q _18992_/S vssd1 vssd1 vccd1 vccd1 _18989_/X sky130_fd_sc_hd__mux2_1
XFILLER_227_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12657__B1 _12656_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21462__RESET_B repeater245/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater155 _18875_/S vssd1 vssd1 vccd1 vccd1 _18680_/S sky130_fd_sc_hd__buf_8
Xrepeater166 _18906_/S vssd1 vssd1 vccd1 vccd1 _18784_/S sky130_fd_sc_hd__buf_6
XFILLER_238_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20951_ _20951_/CLK _20951_/D repeater272/X vssd1 vssd1 vccd1 vccd1 _20951_/Q sky130_fd_sc_hd__dfrtp_1
Xrepeater177 _18666_/S vssd1 vssd1 vccd1 vccd1 _18644_/S sky130_fd_sc_hd__buf_6
XPHY_4309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater188 repeater270/X vssd1 vssd1 vccd1 vccd1 repeater188/X sky130_fd_sc_hd__buf_6
Xrepeater199 repeater209/X vssd1 vssd1 vccd1 vccd1 repeater199/X sky130_fd_sc_hd__clkbuf_8
XFILLER_27_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15523__A _15523_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20882_ _21444_/CLK _20882_/D repeater244/X vssd1 vssd1 vccd1 vccd1 _20882_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13082__B1 _12849_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_92_HCLK_A clkbuf_4_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19196__S0 _20123_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18848__A0 _18848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21434_ _21438_/CLK _21434_/D repeater236/X vssd1 vssd1 vccd1 vccd1 _21434_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17169__B _17169_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16323__A1 _19375_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21365_ _21366_/CLK _21365_/D repeater254/X vssd1 vssd1 vccd1 vccd1 _21365_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_174_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20316_ _20316_/CLK _20316_/D repeater262/X vssd1 vssd1 vccd1 vccd1 _20316_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_123_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21296_ _21302_/CLK _21296_/D repeater208/X vssd1 vssd1 vccd1 vccd1 _21296_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_89_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17185__A _20700_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20247_ _21421_/CLK _20247_/D repeater214/X vssd1 vssd1 vccd1 vccd1 _20247_/Q sky130_fd_sc_hd__dfrtp_1
X_10000_ _20017_/Q vssd1 vssd1 vccd1 vccd1 _10000_/X sky130_fd_sc_hd__buf_1
X_20178_ _21485_/CLK _20178_/D repeater200/X vssd1 vssd1 vccd1 vccd1 _20178_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_76_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09989_ _20022_/Q _09988_/B _09988_/Y vssd1 vssd1 vccd1 vccd1 _17038_/A sky130_fd_sc_hd__o21ai_1
XFILLER_237_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11951_ _11951_/A _11951_/B vssd1 vssd1 vccd1 vccd1 _11952_/A sky130_fd_sc_hd__or2_1
XFILLER_44_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10902_ _11584_/B vssd1 vssd1 vccd1 vccd1 _17019_/A sky130_fd_sc_hd__inv_2
X_14670_ _14657_/X _14534_/X _14663_/B _14669_/X vssd1 vssd1 vccd1 vccd1 _20173_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_83_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11882_ _11878_/Y _10983_/A _11881_/Y vssd1 vssd1 vccd1 vccd1 _11885_/A sky130_fd_sc_hd__o21ai_1
XFILLER_233_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10833_ _10833_/A vssd1 vssd1 vccd1 vccd1 _10833_/Y sky130_fd_sc_hd__inv_2
X_13621_ _20387_/Q _13619_/X _13560_/X _13620_/X vssd1 vssd1 vccd1 vccd1 _20387_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_83_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_241_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16340_ _16340_/A vssd1 vssd1 vccd1 vccd1 _16340_/X sky130_fd_sc_hd__clkbuf_2
X_10764_ _10764_/A _10821_/A vssd1 vssd1 vccd1 vccd1 _10765_/B sky130_fd_sc_hd__or2_2
X_13552_ _20424_/Q _13549_/X _13550_/X _13551_/X vssd1 vssd1 vccd1 vccd1 _20424_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_198_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16011__B1 _16009_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12503_ _19882_/Q _12503_/B vssd1 vssd1 vccd1 vccd1 _16569_/A sky130_fd_sc_hd__or2_1
X_13483_ _13483_/A vssd1 vssd1 vccd1 vccd1 _13483_/X sky130_fd_sc_hd__buf_1
X_16271_ _19401_/Q _16269_/X _16120_/X _16270_/X vssd1 vssd1 vccd1 vccd1 _19401_/D
+ sky130_fd_sc_hd__a22o_1
X_10695_ _21325_/Q _10693_/Y _10712_/A _10655_/B vssd1 vssd1 vccd1 vccd1 _21325_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_13_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12792__A _12804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19187__S0 _19280_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18010_ _18352_/X _17947_/X _18295_/X _17948_/X vssd1 vssd1 vccd1 vccd1 _18014_/A
+ sky130_fd_sc_hd__o22ai_2
XANTENNA__13376__A1 _20502_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15222_ _20481_/Q vssd1 vssd1 vccd1 vccd1 _15222_/Y sky130_fd_sc_hd__inv_2
X_12434_ _12434_/A vssd1 vssd1 vccd1 vccd1 _12434_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18839__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15153_ _15111_/Y _20050_/Q _15151_/Y _20060_/Q _15152_/X vssd1 vssd1 vccd1 vccd1
+ _15157_/C sky130_fd_sc_hd__o221a_1
X_12365_ _12089_/X _12319_/B _12364_/X _12362_/Y vssd1 vssd1 vccd1 vccd1 _20966_/D
+ sky130_fd_sc_hd__a211oi_2
X_11316_ _12506_/A _11316_/B vssd1 vssd1 vccd1 vccd1 _11316_/X sky130_fd_sc_hd__or2_2
XFILLER_153_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20014__RESET_B repeater233/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14104_ _20538_/Q vssd1 vssd1 vccd1 vccd1 _17809_/A sky130_fd_sc_hd__inv_2
XFILLER_181_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15084_ _15084_/A _15084_/B vssd1 vssd1 vccd1 vccd1 _15169_/A sky130_fd_sc_hd__or2_1
X_19961_ _19961_/CLK _19961_/D repeater185/X vssd1 vssd1 vccd1 vccd1 _19961_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_153_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17807__B _17807_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12296_ _20525_/Q vssd1 vssd1 vccd1 vccd1 _12296_/Y sky130_fd_sc_hd__inv_2
X_14035_ _13865_/B _14034_/A _20293_/Q _14037_/A _13980_/X vssd1 vssd1 vccd1 vccd1
+ _20293_/D sky130_fd_sc_hd__o221a_1
X_18912_ _17159_/Y _20035_/Q _18912_/S vssd1 vssd1 vccd1 vccd1 _18912_/X sky130_fd_sc_hd__mux2_1
X_11247_ _19060_/X _11244_/X _21192_/Q _11245_/X vssd1 vssd1 vccd1 vccd1 _21192_/D
+ sky130_fd_sc_hd__a22o_1
X_19892_ _21141_/CLK _19892_/D repeater192/X vssd1 vssd1 vccd1 vccd1 _19892_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_141_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18843_ _18842_/X _10611_/Y _18891_/S vssd1 vssd1 vccd1 vccd1 _18843_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09606__A _13110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11178_ _11176_/A _11176_/B _11176_/Y vssd1 vssd1 vccd1 vccd1 _21219_/D sky130_fd_sc_hd__a21oi_1
XFILLER_122_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10129_ _20788_/Q vssd1 vssd1 vccd1 vccd1 _10129_/Y sky130_fd_sc_hd__inv_2
X_18774_ _18845_/A0 _10479_/Y _18896_/S vssd1 vssd1 vccd1 vccd1 _18774_/X sky130_fd_sc_hd__mux2_1
X_15986_ _15993_/A vssd1 vssd1 vccd1 vccd1 _15986_/X sky130_fd_sc_hd__buf_1
XFILLER_94_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17725_ _21192_/Q vssd1 vssd1 vccd1 vccd1 _17725_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17542__B _17542_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14937_ _20590_/Q vssd1 vssd1 vccd1 vccd1 _14937_/Y sky130_fd_sc_hd__inv_2
XFILLER_94_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15343__A _15421_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17656_ _18732_/X _17472_/X _18731_/X _17474_/X vssd1 vssd1 vccd1 vccd1 _17656_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_36_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14868_ _14962_/B _14868_/B vssd1 vssd1 vccd1 vccd1 _14991_/A sky130_fd_sc_hd__or2_1
XFILLER_235_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16607_ _19990_/Q vssd1 vssd1 vccd1 vccd1 _16607_/Y sky130_fd_sc_hd__inv_2
X_13819_ _20608_/Q vssd1 vssd1 vccd1 vccd1 _13819_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13064__B1 _13001_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17587_ _17548_/X _17559_/X _17560_/X _17568_/X _17586_/X vssd1 vssd1 vccd1 vccd1
+ _17587_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_189_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14799_ _14795_/Y _14797_/A _20118_/Q _14796_/A vssd1 vssd1 vccd1 vccd1 _14800_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_16_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19326_ _20137_/CLK _19326_/D vssd1 vssd1 vccd1 vccd1 _19326_/Q sky130_fd_sc_hd__dfxtp_1
X_16538_ _19995_/Q vssd1 vssd1 vccd1 vccd1 _16539_/A sky130_fd_sc_hd__inv_2
XFILLER_177_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20855__RESET_B repeater243/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12811__A0 _12809_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19257_ _17257_/Y _17258_/Y _17259_/Y _17260_/Y _20130_/Q _20131_/Q vssd1 vssd1 vccd1
+ vccd1 _19257_/X sky130_fd_sc_hd__mux4_1
X_16469_ _19299_/Q _16466_/X _16277_/X _16468_/X vssd1 vssd1 vccd1 vccd1 _19299_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19178__S0 _19280_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18208_ _17079_/Y _12051_/Y _18908_/S vssd1 vssd1 vccd1 vccd1 _18208_/X sky130_fd_sc_hd__mux2_1
XFILLER_163_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19188_ _19547_/Q _19539_/Q _19531_/Q _19515_/Q _19280_/S0 _20122_/Q vssd1 vssd1
+ vccd1 vccd1 _19188_/X sky130_fd_sc_hd__mux4_2
X_18139_ _18845_/A0 _13755_/Y _18896_/S vssd1 vssd1 vccd1 vccd1 _18139_/X sky130_fd_sc_hd__mux2_1
XFILLER_163_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21150_ _21151_/CLK _21150_/D repeater224/X vssd1 vssd1 vccd1 vccd1 _21150_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_172_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20101_ _20101_/CLK _20101_/D repeater259/X vssd1 vssd1 vccd1 vccd1 _20101_/Q sky130_fd_sc_hd__dfrtp_1
X_09912_ _09912_/A _09912_/B vssd1 vssd1 vccd1 vccd1 _17023_/A sky130_fd_sc_hd__or2_1
X_21081_ _21087_/CLK _21081_/D repeater228/X vssd1 vssd1 vccd1 vccd1 _21081_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_113_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20032_ _21481_/CLK _20032_/D repeater205/X vssd1 vssd1 vccd1 vccd1 _20032_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_101_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09843_ _21440_/Q vssd1 vssd1 vccd1 vccd1 _09876_/A sky130_fd_sc_hd__inv_2
XANTENNA__17805__B2 _17797_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_219_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09774_ _21460_/Q vssd1 vssd1 vccd1 vccd1 _09777_/A sky130_fd_sc_hd__inv_2
XFILLER_39_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_61_HCLK clkbuf_4_14_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _21477_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_227_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20934_ _20943_/CLK _20934_/D repeater275/X vssd1 vssd1 vccd1 vccd1 _20934_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_54_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20865_ _21444_/CLK _20865_/D repeater247/X vssd1 vssd1 vccd1 vccd1 _20865_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_42_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12802__B1 _11733_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20796_ _21407_/CLK _20796_/D repeater252/X vssd1 vssd1 vccd1 vccd1 _20796_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19169__S0 _19280_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10480_ _20689_/Q vssd1 vssd1 vccd1 vccd1 _10480_/Y sky130_fd_sc_hd__inv_2
XFILLER_183_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21417_ _21417_/CLK _21417_/D repeater232/X vssd1 vssd1 vccd1 vccd1 _21417_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_185_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18503__S _18775_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09982__B1 _09702_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12150_ _20338_/Q vssd1 vssd1 vccd1 vccd1 _12150_/Y sky130_fd_sc_hd__inv_2
X_21348_ _21349_/CLK _21348_/D repeater210/X vssd1 vssd1 vccd1 vccd1 _21348_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_150_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11101_ _11101_/A vssd1 vssd1 vccd1 vccd1 _11101_/X sky130_fd_sc_hd__buf_1
XFILLER_151_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12081_ _12313_/A vssd1 vssd1 vccd1 vccd1 _12081_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__12869__B1 _12544_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21279_ _21306_/CLK _21279_/D repeater207/X vssd1 vssd1 vccd1 vccd1 _21279_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__21384__RESET_B repeater252/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11032_ _19959_/Q _19958_/Q _16913_/A vssd1 vssd1 vccd1 vccd1 _16922_/A sky130_fd_sc_hd__or3_1
XANTENNA__21129__CLK _21134_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15840_ _19610_/Q _15834_/X _09828_/X _15836_/X vssd1 vssd1 vccd1 vccd1 _19610_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_77_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15283__A1 _20482_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15771_ _19641_/Q _15768_/X _15769_/X _15770_/X vssd1 vssd1 vccd1 vccd1 _19641_/D
+ sky130_fd_sc_hd__a22o_1
X_12983_ _13012_/A vssd1 vssd1 vccd1 vccd1 _12983_/X sky130_fd_sc_hd__buf_1
XFILLER_45_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17510_ _19450_/Q vssd1 vssd1 vccd1 vccd1 _17510_/Y sky130_fd_sc_hd__inv_2
X_14722_ _20148_/Q _14717_/X _13704_/X _14718_/X vssd1 vssd1 vccd1 vccd1 _20148_/D
+ sky130_fd_sc_hd__a22o_1
X_18490_ _17079_/Y _15266_/Y _18908_/S vssd1 vssd1 vccd1 vccd1 _18490_/X sky130_fd_sc_hd__mux2_1
XFILLER_91_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11934_ _11947_/A _11947_/B vssd1 vssd1 vccd1 vccd1 _11934_/Y sky130_fd_sc_hd__nand2_1
XFILLER_17_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17441_ _19441_/Q vssd1 vssd1 vccd1 vccd1 _17441_/Y sky130_fd_sc_hd__inv_2
X_14653_ _20176_/Q _14469_/X _14624_/A _14651_/A vssd1 vssd1 vccd1 vccd1 _20176_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_33_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11865_ _11863_/X _11864_/X _10964_/X _11804_/D vssd1 vssd1 vccd1 vccd1 _11865_/X
+ sky130_fd_sc_hd__o31a_1
XANTENNA_output106_A _17665_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16783__B2 _16777_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13604_ _13631_/A vssd1 vssd1 vccd1 vccd1 _13625_/A sky130_fd_sc_hd__clkbuf_2
XPHY_3972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17372_ _17449_/A _20111_/Q vssd1 vssd1 vccd1 vccd1 _17372_/X sky130_fd_sc_hd__and2_1
X_10816_ _21292_/Q _10815_/Y _10812_/X _10769_/B vssd1 vssd1 vccd1 vccd1 _21292_/D
+ sky130_fd_sc_hd__o211a_1
X_14584_ _14584_/A _14619_/A vssd1 vssd1 vccd1 vccd1 _14585_/B sky130_fd_sc_hd__or2_2
X_11796_ _12638_/A vssd1 vssd1 vccd1 vccd1 _12620_/A sky130_fd_sc_hd__buf_1
XPHY_3983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19111_ _17064_/B _20251_/Q _19111_/S vssd1 vssd1 vccd1 vccd1 _19111_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16323_ _19375_/Q _16319_/X _16014_/X _16320_/X vssd1 vssd1 vccd1 vccd1 _19375_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__20266__RESET_B repeater264/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13535_ _13657_/A _13535_/B vssd1 vssd1 vccd1 vccd1 _13572_/A sky130_fd_sc_hd__or2_2
XFILLER_41_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10747_ _16813_/B _10747_/B vssd1 vssd1 vccd1 vccd1 _16853_/B sky130_fd_sc_hd__or2_1
XANTENNA_repeater256_A repeater257/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19042_ _16816_/X _20827_/Q _19046_/S vssd1 vssd1 vccd1 vccd1 _19934_/D sky130_fd_sc_hd__mux2_1
X_16254_ _19410_/Q _16248_/X _16117_/X _16250_/X vssd1 vssd1 vccd1 vccd1 _19410_/D
+ sky130_fd_sc_hd__a22o_1
X_10678_ _10663_/A _10663_/B _10677_/X _10675_/Y vssd1 vssd1 vccd1 vccd1 _21334_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_145_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13466_ _13481_/A vssd1 vssd1 vccd1 vccd1 _13466_/X sky130_fd_sc_hd__buf_1
XFILLER_145_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15205_ _15205_/A vssd1 vssd1 vccd1 vccd1 _15205_/Y sky130_fd_sc_hd__inv_2
X_12417_ _12496_/C _12417_/B _12417_/C vssd1 vssd1 vccd1 vccd1 _20948_/D sky130_fd_sc_hd__nor3_1
XFILLER_138_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16185_ _19443_/Q _16180_/X _16137_/X _16182_/X vssd1 vssd1 vccd1 vccd1 _19443_/D
+ sky130_fd_sc_hd__a22o_1
X_13397_ _20493_/Q _13390_/X _13274_/X _13393_/X vssd1 vssd1 vccd1 vccd1 _20493_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18413__S _18850_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09973__B1 _09670_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12572__A2 _12566_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15136_ _20433_/Q vssd1 vssd1 vccd1 vccd1 _15136_/Y sky130_fd_sc_hd__inv_2
XFILLER_154_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12348_ _20975_/Q _12347_/Y _12344_/X _12329_/B vssd1 vssd1 vccd1 vccd1 _20975_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_245_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15067_ _15093_/A _15067_/B vssd1 vssd1 vccd1 vccd1 _15202_/A sky130_fd_sc_hd__or2_2
XFILLER_4_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12279_ _20929_/Q vssd1 vssd1 vccd1 vccd1 _12398_/C sky130_fd_sc_hd__inv_2
X_19944_ _20841_/CLK _19944_/D repeater251/X vssd1 vssd1 vccd1 vccd1 _19944_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_101_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14018_ _20302_/Q _14017_/Y _13988_/A _13879_/B vssd1 vssd1 vccd1 vccd1 _20302_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_141_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_84_HCLK clkbuf_4_12_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _21357_/CLK sky130_fd_sc_hd__clkbuf_16
X_19875_ _21151_/CLK _19875_/D repeater226/X vssd1 vssd1 vccd1 vccd1 _19875_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_96_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__21054__RESET_B repeater225/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11532__B1 _10889_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17799__B1 _18380_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17553__A _17553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18826_ _18825_/X _17366_/Y _18927_/S vssd1 vssd1 vccd1 vccd1 _18826_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18757_ _17533_/Y _17532_/Y _18926_/S vssd1 vssd1 vccd1 vccd1 _18757_/X sky130_fd_sc_hd__mux2_1
X_15969_ _16231_/A vssd1 vssd1 vccd1 vccd1 _15969_/X sky130_fd_sc_hd__buf_1
XANTENNA__13285__B1 _13284_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19669__CLK _19813_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_224_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17708_ _20744_/Q vssd1 vssd1 vccd1 vccd1 _17708_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18688_ _18687_/X _10760_/A _18880_/S vssd1 vssd1 vccd1 vccd1 _18688_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17639_ _17639_/A vssd1 vssd1 vccd1 vccd1 _17639_/X sky130_fd_sc_hd__buf_1
XANTENNA__13037__B1 _12954_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20650_ _20657_/CLK _20650_/D repeater196/X vssd1 vssd1 vccd1 vccd1 _20650_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_23_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19309_ _20142_/CLK _19309_/D vssd1 vssd1 vccd1 vccd1 _19309_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20581_ _20946_/CLK _20581_/D repeater258/X vssd1 vssd1 vccd1 vccd1 _20581_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__14417__A _21486_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17723__B1 _17722_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18323__S _18680_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21202_ _21255_/CLK _21202_/D repeater240/X vssd1 vssd1 vccd1 vccd1 _21202_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_155_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21133_ _21191_/CLK _21133_/D repeater192/X vssd1 vssd1 vccd1 vccd1 _21133_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__14152__A _20552_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21064_ _21134_/CLK _21064_/D repeater230/X vssd1 vssd1 vccd1 vccd1 _21064_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_48_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20015_ _21417_/CLK _20015_/D repeater231/X vssd1 vssd1 vccd1 vccd1 _20015_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_86_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17463__A _21139_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09826_ _21449_/Q vssd1 vssd1 vccd1 vccd1 _15876_/A sky130_fd_sc_hd__buf_1
XFILLER_246_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17182__B _17187_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09757_ _21236_/Q vssd1 vssd1 vccd1 vccd1 _11061_/A sky130_fd_sc_hd__inv_2
XFILLER_73_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09688_ _10894_/A vssd1 vssd1 vccd1 vccd1 _09688_/X sky130_fd_sc_hd__clkbuf_4
XPHY_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20706__RESET_B repeater210/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20917_ _21196_/CLK _20917_/D repeater218/X vssd1 vssd1 vccd1 vccd1 _20917_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13028__B1 _12860_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11650_ _18983_/X _11640_/A _21097_/Q _11646_/X vssd1 vssd1 vccd1 vccd1 _21097_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_230_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20848_ _20857_/CLK _20848_/D repeater244/X vssd1 vssd1 vccd1 vccd1 _20848_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_42_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10601_ _20769_/Q vssd1 vssd1 vccd1 vccd1 _10601_/Y sky130_fd_sc_hd__inv_2
XPHY_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11581_ _21126_/Q _11577_/Y _19357_/Q _11577_/A _16740_/A vssd1 vssd1 vccd1 vccd1
+ _21126_/D sky130_fd_sc_hd__o221a_1
XFILLER_167_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20779_ _21147_/CLK _20779_/D repeater215/X vssd1 vssd1 vccd1 vccd1 _20779_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17714__B1 _17713_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10532_ _21338_/Q vssd1 vssd1 vccd1 vccd1 _10534_/A sky130_fd_sc_hd__inv_2
XFILLER_155_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13320_ _20534_/Q _13315_/X _13163_/X _13316_/X vssd1 vssd1 vccd1 vccd1 _20534_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10463_ _21305_/Q _10461_/Y _10781_/A _20694_/Q vssd1 vssd1 vccd1 vccd1 _10463_/X
+ sky130_fd_sc_hd__o22a_1
X_13251_ _20567_/Q _13248_/X _13169_/X _13249_/X vssd1 vssd1 vccd1 vccd1 _20567_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18233__S _18236_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09955__B1 _09682_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12202_ _20950_/Q _12201_/Y _12304_/A _20332_/Q vssd1 vssd1 vccd1 vccd1 _12202_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_170_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13182_ _13182_/A _13182_/B _13182_/C vssd1 vssd1 vccd1 vccd1 _13182_/X sky130_fd_sc_hd__and3_1
XANTENNA_input67_A HWDATA[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10394_ _10394_/A vssd1 vssd1 vccd1 vccd1 _10394_/Y sky130_fd_sc_hd__inv_2
XFILLER_135_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11686__A _12550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12133_ _20965_/Q vssd1 vssd1 vccd1 vccd1 _12318_/A sky130_fd_sc_hd__inv_2
X_17990_ _20655_/Q vssd1 vssd1 vccd1 vccd1 _17990_/Y sky130_fd_sc_hd__inv_2
XFILLER_123_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12064_ _20981_/Q vssd1 vssd1 vccd1 vccd1 _12064_/Y sky130_fd_sc_hd__inv_2
X_16941_ _19964_/Q vssd1 vssd1 vccd1 vccd1 _16941_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19064__S _19910_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11015_ _11590_/A vssd1 vssd1 vccd1 vccd1 _11017_/A sky130_fd_sc_hd__inv_2
XFILLER_1_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19660_ _20172_/CLK _19660_/D vssd1 vssd1 vccd1 vccd1 _19660_/Q sky130_fd_sc_hd__dfxtp_1
X_16872_ _16872_/A vssd1 vssd1 vccd1 vccd1 _16872_/Y sky130_fd_sc_hd__inv_2
XFILLER_226_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18611_ _17281_/X _17832_/Y _18835_/S vssd1 vssd1 vccd1 vccd1 _18611_/X sky130_fd_sc_hd__mux2_1
XFILLER_93_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15823_ _19618_/Q _15817_/X _09828_/X _15819_/X vssd1 vssd1 vccd1 vccd1 _19618_/D
+ sky130_fd_sc_hd__a22o_1
X_19591_ _20890_/CLK _19591_/D vssd1 vssd1 vccd1 vccd1 _19591_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18542_ _18541_/X _20582_/Q _18907_/S vssd1 vssd1 vccd1 vccd1 _18542_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15754_ _19647_/Q _15750_/X _15703_/X _15751_/X vssd1 vssd1 vccd1 vccd1 _19647_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_234_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12966_ _14686_/B vssd1 vssd1 vccd1 vccd1 _12966_/X sky130_fd_sc_hd__buf_1
XFILLER_73_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14705_ _14705_/A vssd1 vssd1 vccd1 vccd1 _14724_/A sky130_fd_sc_hd__inv_2
X_18473_ _18472_/X _14431_/Y _18897_/S vssd1 vssd1 vccd1 vccd1 _18473_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11917_ _19117_/X vssd1 vssd1 vccd1 vccd1 _11917_/X sky130_fd_sc_hd__buf_1
X_15685_ _19679_/Q _15681_/X _15590_/X _15682_/X vssd1 vssd1 vccd1 vccd1 _19679_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12897_ _12891_/X _20735_/Q _12897_/S vssd1 vssd1 vccd1 vccd1 _20735_/D sky130_fd_sc_hd__mux2_1
XANTENNA__18408__S _18907_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17424_ _19585_/Q vssd1 vssd1 vccd1 vccd1 _17425_/A sky130_fd_sc_hd__inv_2
XPHY_4492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14636_ _14636_/A _14636_/B _14636_/C vssd1 vssd1 vccd1 vccd1 _20186_/D sky130_fd_sc_hd__nor3_1
X_11848_ _11848_/A _11848_/B vssd1 vssd1 vccd1 vccd1 _11848_/X sky130_fd_sc_hd__or2_1
XFILLER_220_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17355_ _19608_/Q vssd1 vssd1 vccd1 vccd1 _17355_/Y sky130_fd_sc_hd__inv_2
XFILLER_220_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14567_ _14567_/A _14651_/A vssd1 vssd1 vccd1 vccd1 _14568_/B sky130_fd_sc_hd__or2_1
X_11779_ _15310_/A _16597_/A _11413_/B vssd1 vssd1 vccd1 vccd1 _11780_/S sky130_fd_sc_hd__o21ai_1
X_16306_ _16306_/A vssd1 vssd1 vccd1 vccd1 _16306_/X sky130_fd_sc_hd__buf_1
X_13518_ _20434_/Q _13514_/X _13452_/X _13515_/X vssd1 vssd1 vccd1 vccd1 _20434_/D
+ sky130_fd_sc_hd__a22o_1
X_17286_ _17286_/A vssd1 vssd1 vccd1 vccd1 _17286_/X sky130_fd_sc_hd__buf_1
XFILLER_146_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14498_ _14498_/A _14515_/A vssd1 vssd1 vccd1 vccd1 _14513_/A sky130_fd_sc_hd__or2_1
XFILLER_158_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19025_ _16890_/Y _20398_/Q _19026_/S vssd1 vssd1 vccd1 vccd1 _19951_/D sky130_fd_sc_hd__mux2_1
X_16237_ _16237_/A vssd1 vssd1 vccd1 vccd1 _16237_/X sky130_fd_sc_hd__buf_2
XFILLER_146_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13449_ _13710_/A vssd1 vssd1 vccd1 vccd1 _13449_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__18143__S _18669_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16452__A _16459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16168_ _16174_/A vssd1 vssd1 vccd1 vccd1 _16168_/X sky130_fd_sc_hd__buf_1
XFILLER_115_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15119_ _20461_/Q vssd1 vssd1 vccd1 vccd1 _15119_/Y sky130_fd_sc_hd__inv_2
XFILLER_114_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16099_ _19483_/Q _16094_/X _15871_/X _16096_/X vssd1 vssd1 vccd1 vccd1 _19483_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_114_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19927_ _20841_/CLK _19927_/D repeater256/X vssd1 vssd1 vccd1 vccd1 _19927_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_228_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19858_ _21162_/CLK _19858_/D repeater227/X vssd1 vssd1 vccd1 vccd1 _19858_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_110_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09611_ _11489_/C _11200_/A vssd1 vssd1 vccd1 vccd1 _11182_/A sky130_fd_sc_hd__or2_1
X_18809_ _18808_/X _10629_/Y _18879_/S vssd1 vssd1 vccd1 vccd1 _18809_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13258__A0 _13254_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19789_ _19789_/CLK _19789_/D vssd1 vssd1 vccd1 vccd1 _19789_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20870__RESET_B repeater238/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20188__RESET_B repeater200/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18318__S _18667_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20117__RESET_B repeater247/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20702_ _21125_/CLK _20702_/D repeater190/X vssd1 vssd1 vccd1 vccd1 _20702_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_212_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20633_ _21481_/CLK _20633_/D repeater206/X vssd1 vssd1 vccd1 vccd1 _20633_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20564_ _20724_/CLK _20564_/D repeater264/X vssd1 vssd1 vccd1 vccd1 _20564_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20495_ _20495_/CLK _20495_/D repeater273/X vssd1 vssd1 vccd1 vccd1 _20495_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__12890__A input38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_147_HCLK_A clkbuf_opt_1_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11744__B1 _11743_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21116_ _21120_/CLK _21116_/D repeater233/X vssd1 vssd1 vccd1 vccd1 _21116_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_59_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13497__B1 _13424_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21047_ _21164_/CLK _21047_/D repeater226/X vssd1 vssd1 vccd1 vccd1 _21047_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__20958__RESET_B repeater186/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15706__A _16016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09809_ _16619_/A _16620_/B _09795_/A vssd1 vssd1 vccd1 vccd1 _09809_/X sky130_fd_sc_hd__o21a_1
XFILLER_75_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12820_ _12847_/A vssd1 vssd1 vccd1 vccd1 _12841_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_216_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12751_ _12751_/A _12751_/B vssd1 vssd1 vccd1 vccd1 _12751_/Y sky130_fd_sc_hd__nor2_1
XPHY_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18228__S _18236_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17935__B1 _18540_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11702_ _21077_/Q _11697_/X _11686_/X _11699_/X vssd1 vssd1 vccd1 vccd1 _21077_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15470_ _15479_/A vssd1 vssd1 vccd1 vccd1 _15481_/A sky130_fd_sc_hd__inv_2
XPHY_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12682_ _20829_/Q _12679_/X _09633_/X _12680_/X vssd1 vssd1 vccd1 vccd1 _20829_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14421_ _20237_/Q vssd1 vssd1 vccd1 vccd1 _14421_/Y sky130_fd_sc_hd__inv_2
XPHY_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11633_ _21106_/Q _11632_/Y _11623_/B _11628_/A vssd1 vssd1 vccd1 vccd1 _21106_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13421__B1 _13418_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17140_ _17169_/C _17140_/B _17838_/A vssd1 vssd1 vccd1 vccd1 _17141_/A sky130_fd_sc_hd__or3_4
X_14352_ _20216_/Q vssd1 vssd1 vccd1 vccd1 _14501_/A sky130_fd_sc_hd__inv_2
XPHY_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11564_ _16335_/A vssd1 vssd1 vccd1 vccd1 _13166_/A sky130_fd_sc_hd__buf_4
XPHY_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18360__A0 _18848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13303_ _20545_/Q _13300_/X _13140_/X _13302_/X vssd1 vssd1 vccd1 vccd1 _20545_/D
+ sky130_fd_sc_hd__a22o_1
X_17071_ _19889_/D vssd1 vssd1 vccd1 vccd1 _17076_/C sky130_fd_sc_hd__inv_2
XANTENNA__19059__S _19910_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10515_ _10760_/A _20672_/Q _10769_/A _20682_/Q _10514_/X vssd1 vssd1 vccd1 vccd1
+ _10522_/C sky130_fd_sc_hd__o221a_1
X_11495_ _17549_/A _14256_/B vssd1 vssd1 vccd1 vccd1 _11511_/B sky130_fd_sc_hd__or2_1
X_14283_ _20123_/Q _14283_/B vssd1 vssd1 vccd1 vccd1 _14783_/B sky130_fd_sc_hd__nand2_1
XFILLER_155_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16022_ _16028_/A vssd1 vssd1 vccd1 vccd1 _16029_/A sky130_fd_sc_hd__inv_2
X_10446_ _10446_/A _10446_/B _10446_/C _10446_/D vssd1 vssd1 vccd1 vccd1 _10523_/A
+ sky130_fd_sc_hd__and4_1
X_13234_ _13249_/A vssd1 vssd1 vccd1 vccd1 _13234_/X sky130_fd_sc_hd__buf_1
XANTENNA__18898__S _18898_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13165_ _13165_/A vssd1 vssd1 vccd1 vccd1 _13165_/X sky130_fd_sc_hd__buf_1
X_10377_ _10377_/A vssd1 vssd1 vccd1 vccd1 _10377_/Y sky130_fd_sc_hd__inv_2
XANTENNA_repeater219_A repeater220/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_69_HCLK_A clkbuf_opt_7_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12116_ _12324_/A _20385_/Q _20967_/Q _17937_/A vssd1 vssd1 vccd1 vccd1 _12116_/X
+ sky130_fd_sc_hd__o22a_1
X_17973_ _17925_/X _17973_/B _17973_/C vssd1 vssd1 vccd1 vccd1 _17973_/Y sky130_fd_sc_hd__nand3b_4
XFILLER_69_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13096_ _20639_/Q _13092_/X _12957_/X _13093_/X vssd1 vssd1 vccd1 vccd1 _20639_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_112_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16924_ _16927_/B _16923_/X _16915_/X vssd1 vssd1 vccd1 vccd1 _16924_/X sky130_fd_sc_hd__o21a_1
X_12047_ _20980_/Q _12042_/Y _12331_/A _20392_/Q _12046_/X vssd1 vssd1 vccd1 vccd1
+ _12060_/B sky130_fd_sc_hd__o221a_1
X_19712_ _19776_/CLK _19712_/D vssd1 vssd1 vccd1 vccd1 _19712_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__20699__RESET_B repeater210/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_238_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16855_ _19943_/Q vssd1 vssd1 vccd1 vccd1 _16858_/A sky130_fd_sc_hd__inv_2
X_19643_ _20327_/CLK _19643_/D vssd1 vssd1 vccd1 vccd1 _19643_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15806_ _19626_/Q _15800_/X _09828_/X _15802_/X vssd1 vssd1 vccd1 vccd1 _19626_/D
+ sky130_fd_sc_hd__a22o_1
X_19574_ _20890_/CLK _19574_/D vssd1 vssd1 vccd1 vccd1 _19574_/Q sky130_fd_sc_hd__dfxtp_1
X_16786_ _16786_/A vssd1 vssd1 vccd1 vccd1 _16791_/B sky130_fd_sc_hd__inv_2
XANTENNA__18179__A0 _18848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13998_ _13972_/B _13885_/B _13996_/Y _13991_/X vssd1 vssd1 vccd1 vccd1 _20309_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_241_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_114_HCLK clkbuf_opt_3_HCLK/A vssd1 vssd1 vccd1 vccd1 _20476_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_234_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18525_ _17079_/Y _15239_/Y _18908_/S vssd1 vssd1 vccd1 vccd1 _18525_/X sky130_fd_sc_hd__mux2_1
XANTENNA__20281__RESET_B repeater263/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15737_ _15737_/A vssd1 vssd1 vccd1 vccd1 _15737_/X sky130_fd_sc_hd__buf_1
XFILLER_45_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12949_ _15377_/A vssd1 vssd1 vccd1 vccd1 _14258_/A sky130_fd_sc_hd__buf_2
XANTENNA__18138__S _18910_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_234_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20210__RESET_B repeater203/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18456_ _18455_/X _21358_/Q _18850_/S vssd1 vssd1 vccd1 vccd1 _18456_/X sky130_fd_sc_hd__mux2_1
XFILLER_178_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15668_ _19689_/Q _15666_/X _15585_/X _15667_/X vssd1 vssd1 vccd1 vccd1 _19689_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_221_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17407_ _19497_/Q vssd1 vssd1 vccd1 vccd1 _17407_/Y sky130_fd_sc_hd__inv_2
X_14619_ _14619_/A vssd1 vssd1 vccd1 vccd1 _14619_/Y sky130_fd_sc_hd__inv_2
XFILLER_194_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18387_ _17079_/Y _15265_/Y _18908_/S vssd1 vssd1 vccd1 vccd1 _18387_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13412__B1 _13216_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15599_ _19725_/Q _15596_/X _15469_/X _15598_/X vssd1 vssd1 vccd1 vccd1 _19725_/D
+ sky130_fd_sc_hd__a22o_1
X_17338_ _19520_/Q vssd1 vssd1 vccd1 vccd1 _17338_/Y sky130_fd_sc_hd__inv_2
XFILLER_147_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19908__D _19908_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17269_ _19326_/Q vssd1 vssd1 vccd1 vccd1 _17269_/Y sky130_fd_sc_hd__inv_2
XFILLER_146_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19008_ _16961_/X _20415_/Q _19019_/S vssd1 vssd1 vccd1 vccd1 _19968_/D sky130_fd_sc_hd__mux2_1
X_20280_ _20286_/CLK _20280_/D repeater262/X vssd1 vssd1 vccd1 vccd1 _20280_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_134_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20834__CLK _20930_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18601__S _18903_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_216_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15526__A _15592_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14430__A _21480_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20369__RESET_B repeater187/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13046__A _13046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_2_0_HCLK clkbuf_4_3_0_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_opt_2_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_231_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17917__B1 _18460_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18590__A0 _18589_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_196_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13403__B1 _13284_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20616_ _20622_/CLK _20616_/D repeater195/X vssd1 vssd1 vccd1 vccd1 _20616_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__18342__A0 _17079_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20547_ _20947_/CLK _20547_/D repeater266/X vssd1 vssd1 vccd1 vccd1 _20547_/Q sky130_fd_sc_hd__dfrtp_2
X_10300_ _20732_/Q vssd1 vssd1 vccd1 vccd1 _18083_/A sky130_fd_sc_hd__inv_2
X_11280_ _11280_/A _11299_/A vssd1 vssd1 vccd1 vccd1 _11284_/B sky130_fd_sc_hd__nand2_1
XFILLER_180_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20478_ _20480_/CLK _20478_/D repeater183/X vssd1 vssd1 vccd1 vccd1 _20478_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_10_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10231_ _21372_/Q vssd1 vssd1 vccd1 vccd1 _10287_/A sky130_fd_sc_hd__inv_2
XFILLER_193_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18511__S _18909_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12390__B1 _12359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10162_ _10162_/A _10175_/A _10162_/C vssd1 vssd1 vccd1 vccd1 _10172_/A sky130_fd_sc_hd__or3_4
XFILLER_79_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14970_ _14989_/A vssd1 vssd1 vccd1 vccd1 _14970_/X sky130_fd_sc_hd__buf_2
X_10093_ _20799_/Q vssd1 vssd1 vccd1 vccd1 _10093_/Y sky130_fd_sc_hd__inv_2
XFILLER_248_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_137_HCLK clkbuf_4_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _21374_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__20721__RESET_B repeater264/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13921_ _20642_/Q _20299_/Q _20642_/Q _20299_/Q vssd1 vssd1 vccd1 vccd1 _13921_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_208_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16640_ _19855_/Q _15289_/B _15290_/B vssd1 vssd1 vccd1 vccd1 _16640_/X sky130_fd_sc_hd__a21bo_1
X_13852_ _20309_/Q vssd1 vssd1 vccd1 vccd1 _13972_/B sky130_fd_sc_hd__inv_2
XFILLER_35_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12803_ _12803_/A vssd1 vssd1 vccd1 vccd1 _12803_/X sky130_fd_sc_hd__buf_1
X_16571_ _20001_/Q _20000_/Q vssd1 vssd1 vccd1 vccd1 _16621_/A sky130_fd_sc_hd__or2_1
X_13783_ _20619_/Q vssd1 vssd1 vccd1 vccd1 _17978_/A sky130_fd_sc_hd__inv_2
XFILLER_27_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13642__B1 _13432_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_216_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10995_ _21018_/Q _10995_/B vssd1 vssd1 vccd1 vccd1 _11896_/B sky130_fd_sc_hd__nand2_1
X_18310_ _18309_/X _14417_/Y _18897_/S vssd1 vssd1 vccd1 vccd1 _18310_/X sky130_fd_sc_hd__mux2_1
X_15522_ _19760_/Q _15516_/X _15521_/X _15519_/X vssd1 vssd1 vccd1 vccd1 _19760_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_203_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19290_ _21242_/CLK _20809_/Q vssd1 vssd1 vccd1 vccd1 _19290_/Q sky130_fd_sc_hd__dfxtp_1
X_12734_ _12734_/A _12748_/A vssd1 vssd1 vccd1 vccd1 _12738_/B sky130_fd_sc_hd__or2_1
XFILLER_231_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18241_ _20865_/Q input15/X _18242_/S vssd1 vssd1 vccd1 vccd1 _18241_/X sky130_fd_sc_hd__mux2_2
X_15453_ _19789_/Q _15449_/X _15450_/X _15452_/X vssd1 vssd1 vccd1 vccd1 _19789_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12665_ _20838_/Q _12662_/X _12663_/X _12664_/X vssd1 vssd1 vccd1 vccd1 _20838_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_repeater169_A _18849_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14404_ _14403_/Y _20218_/Q _21472_/Q _14503_/A vssd1 vssd1 vccd1 vccd1 _14404_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11616_ _20015_/Q vssd1 vssd1 vccd1 vccd1 _11617_/A sky130_fd_sc_hd__inv_2
X_18172_ _18848_/A0 _18099_/Y _18644_/S vssd1 vssd1 vccd1 vccd1 _18172_/X sky130_fd_sc_hd__mux2_1
XPHY_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15384_ _19820_/Q _15376_/X _15383_/X _15380_/X vssd1 vssd1 vccd1 vccd1 _19820_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12596_ _20876_/Q _12594_/X _18228_/X _12595_/X vssd1 vssd1 vccd1 vccd1 _20876_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17123_ _19430_/Q vssd1 vssd1 vccd1 vccd1 _17123_/Y sky130_fd_sc_hd__inv_2
X_14335_ _20229_/Q vssd1 vssd1 vccd1 vccd1 _14336_/A sky130_fd_sc_hd__inv_2
XFILLER_51_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11547_ _19912_/Q _16568_/C _16587_/A _16569_/D vssd1 vssd1 vccd1 vccd1 _11547_/X
+ sky130_fd_sc_hd__a211o_1
XPHY_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17054_ _17058_/C _17054_/B _19851_/Q vssd1 vssd1 vccd1 vccd1 _19846_/D sky130_fd_sc_hd__and3_1
X_14266_ _20248_/Q _14257_/X _13704_/X _14260_/X vssd1 vssd1 vccd1 vccd1 _20248_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_output98_A _18068_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11478_ _19101_/X _11474_/X _21157_/Q _11475_/X vssd1 vssd1 vccd1 vccd1 _21157_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19904__RESET_B repeater202/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16005_ _19531_/Q _16000_/X _15975_/X _16002_/X vssd1 vssd1 vccd1 vccd1 _19531_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_130_HCLK_A clkbuf_4_4_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13217_ _13217_/A vssd1 vssd1 vccd1 vccd1 _13217_/X sky130_fd_sc_hd__buf_1
X_10429_ _21300_/Q vssd1 vssd1 vccd1 vccd1 _10776_/A sky130_fd_sc_hd__inv_2
XANTENNA__18421__S _18874_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14197_ _14089_/A _14089_/B _14195_/Y _14193_/X vssd1 vssd1 vccd1 vccd1 _20279_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_140_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13148_ input41/X vssd1 vssd1 vccd1 vccd1 _13148_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_111_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17545__B _17807_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10392__C1 _10381_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15346__A _15424_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17956_ _18534_/X _17954_/X _18529_/X _17955_/X vssd1 vssd1 vccd1 vccd1 _17957_/D
+ sky130_fd_sc_hd__a22o_2
X_13079_ _13098_/A vssd1 vssd1 vccd1 vccd1 _13079_/X sky130_fd_sc_hd__buf_1
XFILLER_78_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16907_ _16910_/B _16906_/Y _16898_/X vssd1 vssd1 vccd1 vccd1 _16907_/X sky130_fd_sc_hd__o21a_1
X_17887_ _18498_/X _17857_/X _18489_/X _17869_/X vssd1 vssd1 vccd1 vccd1 _17887_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_226_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19626_ _19626_/CLK _19626_/D vssd1 vssd1 vccd1 vccd1 _19626_/Q sky130_fd_sc_hd__dfxtp_1
X_16838_ _16877_/A _16838_/B vssd1 vssd1 vccd1 vccd1 _16838_/Y sky130_fd_sc_hd__nor2_1
XFILLER_213_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16769_ _16769_/A vssd1 vssd1 vccd1 vccd1 _16774_/B sky130_fd_sc_hd__inv_2
X_19557_ _19777_/CLK _19557_/D vssd1 vssd1 vccd1 vccd1 _19557_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_202_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18508_ _18845_/A0 _13825_/Y _18896_/S vssd1 vssd1 vccd1 vccd1 _18508_/X sky130_fd_sc_hd__mux2_1
XFILLER_202_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19488_ _19961_/CLK _19488_/D vssd1 vssd1 vccd1 vccd1 _19488_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18439_ _18438_/X _16797_/Y _18667_/S vssd1 vssd1 vccd1 vccd1 _18439_/X sky130_fd_sc_hd__mux2_1
XFILLER_178_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21450_ _21452_/CLK _21450_/D repeater247/X vssd1 vssd1 vccd1 vccd1 _21450_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_193_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18324__A0 _17079_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_18_HCLK clkbuf_4_3_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _21021_/CLK sky130_fd_sc_hd__clkbuf_16
X_20401_ _20809_/CLK _20401_/D repeater188/X vssd1 vssd1 vccd1 vccd1 _20401_/Q sky130_fd_sc_hd__dfrtp_1
Xclkbuf_4_10_0_HCLK clkbuf_3_5_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20004_/CLK sky130_fd_sc_hd__clkbuf_1
X_21381_ _21421_/CLK _21381_/D repeater214/X vssd1 vssd1 vccd1 vccd1 _21381_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_147_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20332_ _20809_/CLK _20332_/D repeater188/X vssd1 vssd1 vccd1 vccd1 _20332_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_135_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20263_ _20724_/CLK _20263_/D repeater264/X vssd1 vssd1 vccd1 vccd1 _20263_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18627__A1 _21373_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18331__S _18748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20194_ _20626_/CLK _20194_/D repeater193/X vssd1 vssd1 vccd1 vccd1 _20194_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_163_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_52_HCLK_A clkbuf_4_14_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_245_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20132__RESET_B repeater249/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17190__B _17193_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10780_ _10780_/A _10793_/A vssd1 vssd1 vccd1 vccd1 _10781_/B sky130_fd_sc_hd__or2_1
XFILLER_25_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18563__A0 _17281_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18506__S _18644_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12450_ _12429_/A _12429_/B _12445_/X _12447_/Y vssd1 vssd1 vccd1 vccd1 _20940_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_40_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11938__B1 _11940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11401_ _11421_/A vssd1 vssd1 vccd1 vccd1 _11401_/X sky130_fd_sc_hd__buf_1
XFILLER_166_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12381_ _20957_/Q _12380_/Y _12373_/X _12312_/B vssd1 vssd1 vccd1 vccd1 _20957_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_165_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14120_ _14120_/A _14120_/B _14120_/C _14120_/D vssd1 vssd1 vccd1 vccd1 _14171_/A
+ sky130_fd_sc_hd__and4_1
X_11332_ _21169_/Q _21168_/Q _21171_/Q _21170_/Q vssd1 vssd1 vccd1 vccd1 _11367_/B
+ sky130_fd_sc_hd__or4_4
XANTENNA__11678__B _15312_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14051_ _20277_/Q vssd1 vssd1 vccd1 vccd1 _14087_/A sky130_fd_sc_hd__inv_2
XANTENNA__19402__CLK _21009_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18618__A1 _20663_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11263_ _20916_/Q _20915_/Q vssd1 vssd1 vccd1 vccd1 _11283_/C sky130_fd_sc_hd__or2_1
XANTENNA__20973__RESET_B repeater187/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18241__S _18242_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13002_ _20691_/Q _12995_/X _13001_/X _12997_/X vssd1 vssd1 vccd1 vccd1 _20691_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17826__C1 _17825_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10214_ _21383_/Q _10213_/Y _10166_/A _10205_/B vssd1 vssd1 vccd1 vccd1 _21383_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__20902__RESET_B repeater217/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11194_ _21217_/Q _11191_/X _10892_/X _11193_/X vssd1 vssd1 vccd1 vccd1 _21217_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_106_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17810_ _17810_/A _17812_/B vssd1 vssd1 vccd1 vccd1 _17810_/Y sky130_fd_sc_hd__nor2_1
X_10145_ _10145_/A vssd1 vssd1 vccd1 vccd1 _10168_/B sky130_fd_sc_hd__inv_2
X_18790_ _17448_/X _21253_/Q _20870_/Q vssd1 vssd1 vccd1 vccd1 _18790_/X sky130_fd_sc_hd__mux2_1
XANTENNA__19552__CLK _19706_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17741_ _19477_/Q vssd1 vssd1 vccd1 vccd1 _17741_/Y sky130_fd_sc_hd__inv_2
XFILLER_248_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14953_ _20107_/Q _14884_/Y _14885_/Y _14884_/A _14952_/X vssd1 vssd1 vccd1 vccd1
+ _20107_/D sky130_fd_sc_hd__o221a_1
X_10076_ _10162_/C _10163_/A _10076_/C _10168_/A vssd1 vssd1 vccd1 vccd1 _10077_/C
+ sky130_fd_sc_hd__or4_4
XANTENNA_output136_A _20982_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19072__S _19908_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13904_ _20665_/Q vssd1 vssd1 vccd1 vccd1 _13904_/Y sky130_fd_sc_hd__inv_2
XFILLER_235_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17672_ _19396_/Q vssd1 vssd1 vccd1 vccd1 _17672_/Y sky130_fd_sc_hd__inv_2
X_14884_ _14884_/A vssd1 vssd1 vccd1 vccd1 _14884_/Y sky130_fd_sc_hd__inv_2
XFILLER_47_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16623_ _16623_/A vssd1 vssd1 vccd1 vccd1 _19999_/D sky130_fd_sc_hd__inv_2
X_19411_ _21001_/CLK _19411_/D vssd1 vssd1 vccd1 vccd1 _19411_/Q sky130_fd_sc_hd__dfxtp_1
X_13835_ _13830_/Y _20177_/Q _20615_/Q _14581_/A _13834_/X vssd1 vssd1 vccd1 vccd1
+ _13836_/D sky130_fd_sc_hd__o221a_1
XFILLER_62_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13615__B1 _13550_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16554_ _16566_/C vssd1 vssd1 vccd1 vccd1 _16554_/Y sky130_fd_sc_hd__inv_2
X_19342_ _19961_/CLK _19342_/D vssd1 vssd1 vccd1 vccd1 _19342_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13766_ _20612_/Q _20189_/Q _13764_/Y _14578_/A vssd1 vssd1 vccd1 vccd1 _13766_/X
+ sky130_fd_sc_hd__o22a_1
X_10978_ _12715_/A _15884_/A vssd1 vssd1 vccd1 vccd1 _11153_/A sky130_fd_sc_hd__or2_1
XFILLER_231_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15505_ _15505_/A _15505_/B _15505_/C vssd1 vssd1 vccd1 vccd1 _15722_/C sky130_fd_sc_hd__or3_4
XANTENNA__15368__B1 _15346_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12717_ _13535_/B _13104_/B vssd1 vssd1 vccd1 vccd1 _12718_/S sky130_fd_sc_hd__or2_1
X_19273_ _17097_/Y _17098_/Y _17099_/Y _17100_/Y _19275_/S0 _21004_/Q vssd1 vssd1
+ vccd1 vccd1 _19273_/X sky130_fd_sc_hd__mux4_1
XFILLER_15_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16485_ _16485_/A vssd1 vssd1 vccd1 vccd1 _18926_/S sky130_fd_sc_hd__clkinv_8
XFILLER_231_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13697_ _20341_/Q _13693_/X _13584_/X _13694_/X vssd1 vssd1 vccd1 vccd1 _20341_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18416__S _18928_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21008__RESET_B repeater235/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18224_ _20848_/Q input28/X _18236_/S vssd1 vssd1 vccd1 vccd1 _18224_/X sky130_fd_sc_hd__mux2_1
XFILLER_175_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15436_ _15442_/A vssd1 vssd1 vccd1 vccd1 _15436_/X sky130_fd_sc_hd__buf_1
XPHY_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12648_ _17083_/A _12815_/A vssd1 vssd1 vccd1 vccd1 _12685_/A sky130_fd_sc_hd__or2_1
XANTENNA__18306__A0 _18848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18155_ _18154_/X _10588_/Y _18775_/S vssd1 vssd1 vccd1 vccd1 _18155_/X sky130_fd_sc_hd__mux2_1
X_15367_ _15367_/A vssd1 vssd1 vccd1 vccd1 _15367_/X sky130_fd_sc_hd__buf_1
XFILLER_8_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12579_ _20885_/Q _12574_/X _18237_/X _12575_/X vssd1 vssd1 vccd1 vccd1 _20885_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17106_ _19774_/Q vssd1 vssd1 vccd1 vccd1 _17106_/Y sky130_fd_sc_hd__inv_2
XFILLER_184_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14318_ _14318_/A vssd1 vssd1 vccd1 vccd1 _14318_/X sky130_fd_sc_hd__buf_1
XFILLER_117_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18086_ _18625_/X _17856_/X _18646_/X _17932_/X vssd1 vssd1 vccd1 vccd1 _18090_/A
+ sky130_fd_sc_hd__o22ai_2
X_15298_ _19864_/Q _15298_/B vssd1 vssd1 vccd1 vccd1 _15299_/B sky130_fd_sc_hd__or2_1
XFILLER_7_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17037_ _17037_/A _17038_/B vssd1 vssd1 vccd1 vccd1 _20021_/D sky130_fd_sc_hd__nor2_1
X_14249_ _14249_/A vssd1 vssd1 vccd1 vccd1 _14249_/X sky130_fd_sc_hd__buf_1
XANTENNA__18151__S _18680_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09790_ _16619_/B _09789_/Y _16620_/A _09788_/X vssd1 vssd1 vccd1 vccd1 _21459_/D
+ sky130_fd_sc_hd__a22oi_1
X_18988_ _21265_/Q _21117_/Q _18992_/S vssd1 vssd1 vccd1 vccd1 _18988_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17939_ _17974_/A vssd1 vssd1 vccd1 vccd1 _17943_/B sky130_fd_sc_hd__buf_2
XFILLER_227_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrepeater156 _18667_/S vssd1 vssd1 vccd1 vccd1 _18875_/S sky130_fd_sc_hd__buf_8
Xrepeater167 _18909_/S vssd1 vssd1 vccd1 vccd1 _18906_/S sky130_fd_sc_hd__buf_8
XFILLER_227_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20950_ _20950_/CLK _20950_/D repeater272/X vssd1 vssd1 vccd1 vccd1 _20950_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_26_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater178 _18874_/S vssd1 vssd1 vccd1 vccd1 _18666_/S sky130_fd_sc_hd__buf_8
XFILLER_39_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrepeater189 repeater270/X vssd1 vssd1 vccd1 vccd1 repeater189/X sky130_fd_sc_hd__buf_8
X_19609_ _21449_/CLK _19609_/D vssd1 vssd1 vccd1 vccd1 _19609_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20881_ _21445_/CLK _20881_/D repeater243/X vssd1 vssd1 vccd1 vccd1 _20881_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_42_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18326__S _18907_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19196__S1 _20124_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21433_ _21433_/CLK _21433_/D repeater236/X vssd1 vssd1 vccd1 vccd1 _21433_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_163_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21364_ _21367_/CLK _21364_/D repeater254/X vssd1 vssd1 vccd1 vccd1 _21364_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__19985__SET_B repeater281/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20315_ _20316_/CLK _20315_/D repeater197/X vssd1 vssd1 vccd1 vccd1 _20315_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_174_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21295_ _21302_/CLK _21295_/D repeater208/X vssd1 vssd1 vccd1 vccd1 _21295_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_150_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20246_ _21421_/CLK _20246_/D repeater214/X vssd1 vssd1 vccd1 vccd1 _20246_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17185__B _17187_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18996__S _19026_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20177_ _21485_/CLK _20177_/D repeater200/X vssd1 vssd1 vccd1 vccd1 _20177_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_190_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09988_ _20022_/Q _09988_/B vssd1 vssd1 vccd1 vccd1 _09988_/Y sky130_fd_sc_hd__nand2_1
XFILLER_67_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11950_ _19109_/X vssd1 vssd1 vccd1 vccd1 _11951_/A sky130_fd_sc_hd__inv_2
XFILLER_85_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17587__B2 _17568_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10901_ _21250_/Q _10888_/A _10900_/X _10890_/A vssd1 vssd1 vccd1 vccd1 _21250_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_29_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11881_ _11881_/A _11881_/B vssd1 vssd1 vccd1 vccd1 _11881_/Y sky130_fd_sc_hd__nand2_1
XFILLER_245_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13620_ _13626_/A vssd1 vssd1 vccd1 vccd1 _13620_/X sky130_fd_sc_hd__buf_1
X_10832_ _10760_/A _10760_/B _10827_/X _10829_/Y vssd1 vssd1 vccd1 vccd1 _21283_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_44_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14270__B1 _13710_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21172__RESET_B repeater216/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_213_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13551_ _13567_/A vssd1 vssd1 vccd1 vccd1 _13551_/X sky130_fd_sc_hd__buf_1
X_10763_ _10763_/A _10763_/B _10825_/A vssd1 vssd1 vccd1 vccd1 _10821_/A sky130_fd_sc_hd__or3_1
XFILLER_13_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18236__S _18236_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12502_ _12502_/A _12502_/B vssd1 vssd1 vccd1 vccd1 _12507_/A sky130_fd_sc_hd__or2_1
XFILLER_157_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16270_ _16270_/A vssd1 vssd1 vccd1 vccd1 _16270_/X sky130_fd_sc_hd__buf_1
X_13482_ input48/X vssd1 vssd1 vccd1 vccd1 _13482_/X sky130_fd_sc_hd__clkbuf_2
X_10694_ _10694_/A vssd1 vssd1 vccd1 vccd1 _10712_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_139_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15221_ _20472_/Q vssd1 vssd1 vccd1 vccd1 _15221_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19187__S1 _20122_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12433_ _12433_/A _12440_/A vssd1 vssd1 vccd1 vccd1 _12434_/A sky130_fd_sc_hd__or2_2
X_15152_ _20441_/Q _15093_/X _20458_/Q _15083_/A vssd1 vssd1 vccd1 vccd1 _15152_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_154_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12364_ _12364_/A vssd1 vssd1 vccd1 vccd1 _12364_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_153_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14103_ _14103_/A vssd1 vssd1 vccd1 vccd1 _14103_/X sky130_fd_sc_hd__buf_1
X_11315_ _11315_/A _20915_/Q _11315_/C vssd1 vssd1 vccd1 vccd1 _11316_/B sky130_fd_sc_hd__or3_1
XANTENNA__19067__S _19908_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14325__A1 _14313_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15083_ _15083_/A _15173_/A vssd1 vssd1 vccd1 vccd1 _15084_/B sky130_fd_sc_hd__or2_1
X_19960_ _20408_/CLK _19960_/D repeater184/X vssd1 vssd1 vccd1 vccd1 _19960_/Q sky130_fd_sc_hd__dfrtp_1
X_12295_ _20928_/Q vssd1 vssd1 vccd1 vccd1 _12476_/A sky130_fd_sc_hd__inv_2
XFILLER_181_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14034_ _14034_/A vssd1 vssd1 vccd1 vccd1 _14037_/A sky130_fd_sc_hd__inv_2
X_18911_ _17171_/Y _20243_/Q _18912_/S vssd1 vssd1 vccd1 vccd1 _18911_/X sky130_fd_sc_hd__mux2_1
X_11246_ _19059_/X _11244_/X _21193_/Q _11245_/X vssd1 vssd1 vccd1 vccd1 _21193_/D
+ sky130_fd_sc_hd__a22o_1
X_19891_ _21141_/CLK _19891_/D repeater192/X vssd1 vssd1 vccd1 vccd1 _19891_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_repeater201_A repeater205/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18842_ _18845_/A0 _10506_/Y _18896_/S vssd1 vssd1 vccd1 vccd1 _18842_/X sky130_fd_sc_hd__mux2_1
X_11177_ _15609_/A _11176_/Y _11170_/A vssd1 vssd1 vccd1 vccd1 _21220_/D sky130_fd_sc_hd__o21a_1
X_10128_ _21388_/Q _10126_/Y _10149_/A _20785_/Q _10127_/X vssd1 vssd1 vccd1 vccd1
+ _10136_/B sky130_fd_sc_hd__o221a_1
XFILLER_121_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15985_ _15985_/A _16229_/B _16325_/C vssd1 vssd1 vccd1 vccd1 _15993_/A sky130_fd_sc_hd__or3_4
X_18773_ _18772_/X _10263_/A _18841_/S vssd1 vssd1 vccd1 vccd1 _18773_/X sky130_fd_sc_hd__mux2_1
XFILLER_209_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17724_ _21142_/Q vssd1 vssd1 vccd1 vccd1 _17724_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14936_ _14914_/Y _20076_/Q _20579_/Q _14962_/B _14935_/X vssd1 vssd1 vccd1 vccd1
+ _14936_/X sky130_fd_sc_hd__a221o_1
X_10059_ _10059_/A vssd1 vssd1 vccd1 vccd1 _10157_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_63_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17578__A1 _18742_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10114__A2 _10081_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17578__B2 _17854_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17655_ _17647_/Y _17177_/B _17649_/X _17654_/X vssd1 vssd1 vccd1 vccd1 _17655_/X
+ sky130_fd_sc_hd__o211a_2
XANTENNA__15589__B1 _15588_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14867_ _14960_/C _14994_/A vssd1 vssd1 vccd1 vccd1 _14868_/B sky130_fd_sc_hd__or2_2
XFILLER_208_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13144__A input43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16606_ _16600_/Y _16605_/X _16588_/A vssd1 vssd1 vccd1 vccd1 _19989_/D sky130_fd_sc_hd__o21ai_1
X_13818_ _20620_/Q vssd1 vssd1 vccd1 vccd1 _13818_/Y sky130_fd_sc_hd__inv_2
X_17586_ _18741_/X _17569_/X _17572_/Y _17578_/X _17585_/X vssd1 vssd1 vccd1 vccd1
+ _17586_/X sky130_fd_sc_hd__o2111a_2
XANTENNA__14261__B1 _14258_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14798_ _20117_/Q vssd1 vssd1 vccd1 vccd1 _14800_/A sky130_fd_sc_hd__buf_1
XFILLER_51_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16537_ _19994_/Q vssd1 vssd1 vccd1 vccd1 _16537_/Y sky130_fd_sc_hd__inv_2
X_19325_ _21234_/CLK _19325_/D vssd1 vssd1 vccd1 vccd1 _19325_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13749_ _20626_/Q vssd1 vssd1 vccd1 vccd1 _13749_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12983__A _13012_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18146__S _18644_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19990__RESET_B repeater217/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19256_ _19252_/X _19253_/X _19254_/X _19255_/X _21005_/Q _21006_/Q vssd1 vssd1 vccd1
+ vccd1 _19256_/X sky130_fd_sc_hd__mux4_2
X_16468_ _16474_/A vssd1 vssd1 vccd1 vccd1 _16468_/X sky130_fd_sc_hd__buf_1
XFILLER_164_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19178__S1 _20122_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18207_ _18206_/X _14886_/Y _18907_/S vssd1 vssd1 vccd1 vccd1 _18207_/X sky130_fd_sc_hd__mux2_2
X_15419_ _19804_/Q _15415_/X _15383_/X _15417_/X vssd1 vssd1 vccd1 vccd1 _19804_/D
+ sky130_fd_sc_hd__a22o_1
X_19187_ _19707_/Q _19571_/Q _19563_/Q _19555_/Q _19280_/S0 _20122_/Q vssd1 vssd1
+ vccd1 vccd1 _19187_/X sky130_fd_sc_hd__mux4_2
X_16399_ _16399_/A vssd1 vssd1 vccd1 vccd1 _16399_/X sky130_fd_sc_hd__buf_1
XFILLER_191_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_3_6_0_HCLK clkbuf_3_7_0_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_6_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_18138_ _18137_/X _12221_/Y _18910_/S vssd1 vssd1 vccd1 vccd1 _18138_/X sky130_fd_sc_hd__mux2_1
XANTENNA__20824__RESET_B repeater251/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18069_ _20801_/Q vssd1 vssd1 vccd1 vccd1 _18069_/Y sky130_fd_sc_hd__inv_2
XFILLER_171_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20100_ _20101_/CLK _20100_/D repeater259/X vssd1 vssd1 vccd1 vccd1 _20100_/Q sky130_fd_sc_hd__dfrtp_1
X_09911_ _17020_/A _09899_/X _20008_/Q _20009_/Q vssd1 vssd1 vccd1 vccd1 _09912_/B
+ sky130_fd_sc_hd__a31oi_1
XFILLER_132_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21080_ _21424_/CLK _21080_/D repeater230/X vssd1 vssd1 vccd1 vccd1 _21080_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_113_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20031_ _21357_/CLK _20031_/D repeater199/X vssd1 vssd1 vccd1 vccd1 _20031_/Q sky130_fd_sc_hd__dfrtp_2
X_09842_ _21442_/Q vssd1 vssd1 vccd1 vccd1 _09847_/A sky130_fd_sc_hd__inv_2
XFILLER_140_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17805__A2 _17788_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09773_ _21461_/Q vssd1 vssd1 vccd1 vccd1 _09775_/A sky130_fd_sc_hd__inv_2
XFILLER_58_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20933_ _20944_/CLK _20933_/D repeater275/X vssd1 vssd1 vccd1 vccd1 _20933_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_227_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20864_ _21444_/CLK _20864_/D repeater246/X vssd1 vssd1 vccd1 vccd1 _20864_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_53_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18518__A0 _18848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12802__A1 _20777_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20795_ _21407_/CLK _20795_/D repeater252/X vssd1 vssd1 vccd1 vccd1 _20795_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19169__S1 _20122_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21416_ _21417_/CLK _21416_/D repeater232/X vssd1 vssd1 vccd1 vccd1 _21416_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_175_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21347_ _21349_/CLK _21347_/D repeater210/X vssd1 vssd1 vccd1 vccd1 _21347_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_190_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11100_ _11100_/A vssd1 vssd1 vccd1 vccd1 _11100_/X sky130_fd_sc_hd__buf_1
XFILLER_150_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12080_ _20960_/Q vssd1 vssd1 vccd1 vccd1 _12313_/A sky130_fd_sc_hd__inv_2
X_21278_ _21306_/CLK _21278_/D repeater207/X vssd1 vssd1 vccd1 vccd1 _21278_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__10860__B _17195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11031_ _19957_/Q _16909_/A vssd1 vssd1 vccd1 vccd1 _16913_/A sky130_fd_sc_hd__or2_2
X_20229_ _21485_/CLK _20229_/D repeater200/X vssd1 vssd1 vccd1 vccd1 _20229_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17924__A _18018_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15770_ _15770_/A vssd1 vssd1 vccd1 vccd1 _15770_/X sky130_fd_sc_hd__clkbuf_2
X_12982_ _13018_/A vssd1 vssd1 vccd1 vccd1 _13012_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_92_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input12_A HADDR[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14721_ _20149_/Q _14717_/X _14264_/X _14718_/X vssd1 vssd1 vccd1 vccd1 _20149_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__21353__RESET_B repeater255/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11933_ _11928_/Y _11930_/A _11932_/X _11929_/A vssd1 vssd1 vccd1 vccd1 _11947_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_217_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17440_ _19328_/Q vssd1 vssd1 vccd1 vccd1 _17440_/Y sky130_fd_sc_hd__inv_2
X_14652_ _20177_/Q _14651_/Y _14642_/X _14568_/B vssd1 vssd1 vccd1 vccd1 _20177_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_27_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11864_ _11864_/A vssd1 vssd1 vccd1 vccd1 _11864_/X sky130_fd_sc_hd__buf_1
XFILLER_232_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16783__A2 _16777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13603_ _17080_/A _13657_/B vssd1 vssd1 vccd1 vccd1 _13631_/A sky130_fd_sc_hd__or2_2
XPHY_3951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17371_ _21433_/Q _17536_/A vssd1 vssd1 vccd1 vccd1 _17371_/X sky130_fd_sc_hd__and2_1
X_10815_ _10815_/A vssd1 vssd1 vccd1 vccd1 _10815_/Y sky130_fd_sc_hd__inv_2
XPHY_3962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14583_ _14583_/A _14583_/B vssd1 vssd1 vccd1 vccd1 _14619_/A sky130_fd_sc_hd__or2_1
XPHY_3973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11795_ _11795_/A vssd1 vssd1 vccd1 vccd1 _12638_/A sky130_fd_sc_hd__clkbuf_2
XPHY_3984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16322_ _19376_/Q _16319_/X _16012_/X _16320_/X vssd1 vssd1 vccd1 vccd1 _19376_/D
+ sky130_fd_sc_hd__a22o_1
X_19110_ _16616_/Y _11916_/Y _19116_/S vssd1 vssd1 vccd1 vccd1 _19110_/X sky130_fd_sc_hd__mux2_1
X_13534_ _13530_/A _13530_/B _20429_/Q _13533_/X vssd1 vssd1 vccd1 vccd1 _20429_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_13_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10746_ _19935_/Q _19936_/Q _10746_/C _16843_/A vssd1 vssd1 vccd1 vccd1 _10747_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_43_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19740__CLK _19765_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19041_ _16820_/Y _20828_/Q _19046_/S vssd1 vssd1 vccd1 vccd1 _19935_/D sky130_fd_sc_hd__mux2_1
X_16253_ _19411_/Q _16248_/X _16115_/X _16250_/X vssd1 vssd1 vccd1 vccd1 _19411_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_159_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13465_ _20461_/Q _13458_/X _13274_/X _13461_/X vssd1 vssd1 vccd1 vccd1 _20461_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_repeater151_A _18902_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10677_ _10677_/A vssd1 vssd1 vccd1 vccd1 _10677_/X sky130_fd_sc_hd__buf_2
XANTENNA_repeater249_A repeater250/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12557__B1 _11741_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15204_ _15093_/X _15067_/B _15202_/Y _15193_/X vssd1 vssd1 vccd1 vccd1 _20052_/D
+ sky130_fd_sc_hd__a211oi_2
X_12416_ _12408_/C _12436_/B _12408_/A vssd1 vssd1 vccd1 vccd1 _12417_/C sky130_fd_sc_hd__o21a_1
X_16184_ _19444_/Q _16180_/X _16135_/X _16182_/X vssd1 vssd1 vccd1 vccd1 _19444_/D
+ sky130_fd_sc_hd__a22o_1
X_13396_ _20494_/Q _13390_/X _13272_/X _13393_/X vssd1 vssd1 vccd1 vccd1 _20494_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_182_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20235__RESET_B repeater203/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15135_ _15132_/Y _20049_/Q _20436_/Q _15062_/A _15134_/X vssd1 vssd1 vccd1 vccd1
+ _15144_/B sky130_fd_sc_hd__o221a_1
X_12347_ _12347_/A vssd1 vssd1 vccd1 vccd1 _12347_/Y sky130_fd_sc_hd__inv_2
XFILLER_153_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output80_A _17865_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15066_ _15066_/A _15205_/A vssd1 vssd1 vccd1 vccd1 _15067_/B sky130_fd_sc_hd__or2_2
X_19943_ _20930_/CLK _19943_/D repeater268/X vssd1 vssd1 vccd1 vccd1 _19943_/Q sky130_fd_sc_hd__dfrtp_1
X_12278_ _12262_/X _12278_/B _12278_/C _12278_/D vssd1 vssd1 vccd1 vccd1 _12302_/C
+ sky130_fd_sc_hd__and4b_1
XFILLER_4_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14017_ _14017_/A _14017_/B vssd1 vssd1 vccd1 vccd1 _14017_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__17834__A _18930_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11229_ _21198_/Q _11225_/X _10898_/X _11226_/X vssd1 vssd1 vccd1 vccd1 _21198_/D
+ sky130_fd_sc_hd__a22o_1
X_19874_ _20042_/CLK _19874_/D repeater219/X vssd1 vssd1 vccd1 vccd1 _19874_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_95_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11532__A1 _21141_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18825_ _17369_/Y _17368_/X _18926_/S vssd1 vssd1 vccd1 vccd1 _18825_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12978__A _13600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15354__A _15354_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18756_ _17535_/Y _09902_/Y _20870_/Q vssd1 vssd1 vccd1 vccd1 _18756_/X sky130_fd_sc_hd__mux2_1
X_15968_ _15978_/A vssd1 vssd1 vccd1 vccd1 _15968_/X sky130_fd_sc_hd__buf_1
XFILLER_209_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__21094__RESET_B repeater226/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17707_ _20504_/Q vssd1 vssd1 vccd1 vccd1 _17707_/Y sky130_fd_sc_hd__inv_2
XFILLER_224_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14919_ _20593_/Q vssd1 vssd1 vccd1 vccd1 _14919_/Y sky130_fd_sc_hd__inv_2
X_18687_ _18686_/X _17708_/Y _18775_/S vssd1 vssd1 vccd1 vccd1 _18687_/X sky130_fd_sc_hd__mux2_1
XFILLER_63_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15899_ _19584_/Q _15896_/X _15791_/X _15897_/X vssd1 vssd1 vccd1 vccd1 _19584_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_63_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17638_ _21077_/Q vssd1 vssd1 vccd1 vccd1 _17638_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14785__A1 _20124_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15982__B1 _15949_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17569_ _17932_/A vssd1 vssd1 vccd1 vccd1 _17569_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__12796__B1 _12699_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19308_ _21167_/CLK _19308_/D vssd1 vssd1 vccd1 vccd1 _19308_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20580_ _20946_/CLK _20580_/D repeater258/X vssd1 vssd1 vccd1 vccd1 _20580_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__09661__B1 _09659_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19239_ _17436_/Y _17437_/Y _17438_/Y _17439_/Y _20130_/Q _20131_/Q vssd1 vssd1 vccd1
+ vccd1 _19239_/X sky130_fd_sc_hd__mux4_1
XFILLER_192_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18604__S _18896_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21201_ _21255_/CLK _21201_/D repeater241/X vssd1 vssd1 vccd1 vccd1 _21201_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_117_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21132_ _21141_/CLK _21132_/D repeater192/X vssd1 vssd1 vccd1 vccd1 _21132_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_235_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21063_ _21087_/CLK _21063_/D repeater227/X vssd1 vssd1 vccd1 vccd1 _21063_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__13049__A _13262_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11523__A1 _21144_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20014_ _21120_/CLK input71/X repeater233/X vssd1 vssd1 vccd1 vccd1 _20014_/Q sky130_fd_sc_hd__dfrtp_1
X_09825_ _15873_/A _09813_/X _09824_/X _09815_/X vssd1 vssd1 vccd1 vccd1 _21450_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_input4_A HADDR[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12888__A _17178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09756_ _20156_/Q vssd1 vssd1 vccd1 vccd1 _09756_/Y sky130_fd_sc_hd__inv_2
XFILLER_246_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_170_HCLK clkbuf_opt_2_HCLK/A vssd1 vssd1 vccd1 vccd1 _19774_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_64_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_107_HCLK_A clkbuf_opt_3_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09687_ input63/X vssd1 vssd1 vccd1 vccd1 _10894_/A sky130_fd_sc_hd__buf_1
XFILLER_54_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20916_ _21196_/CLK _20916_/D repeater218/X vssd1 vssd1 vccd1 vccd1 _20916_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19841__RESET_B repeater226/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19763__CLK _19765_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20847_ _21457_/CLK _20847_/D repeater244/X vssd1 vssd1 vccd1 vccd1 _20847_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10600_ _10540_/B _20740_/Q _10534_/B _20765_/Q _10599_/X vssd1 vssd1 vccd1 vccd1
+ _10605_/C sky130_fd_sc_hd__o221a_1
XANTENNA__12787__B1 _09641_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20746__RESET_B repeater207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11580_ _16545_/A vssd1 vssd1 vccd1 vccd1 _16740_/A sky130_fd_sc_hd__buf_1
XPHY_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20778_ _21379_/CLK _20778_/D repeater214/X vssd1 vssd1 vccd1 vccd1 _20778_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10531_ _21336_/Q vssd1 vssd1 vccd1 vccd1 _10664_/C sky130_fd_sc_hd__inv_2
XFILLER_195_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18514__S _18849_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13250_ _20568_/Q _13248_/X _13166_/X _13249_/X vssd1 vssd1 vccd1 vccd1 _20568_/D
+ sky130_fd_sc_hd__a22o_1
X_10462_ _21305_/Q vssd1 vssd1 vccd1 vccd1 _10781_/A sky130_fd_sc_hd__inv_2
XFILLER_155_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12201_ _20332_/Q vssd1 vssd1 vccd1 vccd1 _12201_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17478__B1 _18795_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11211__B1 _09649_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13181_ _13528_/A _13527_/A _13181_/C _20432_/Q vssd1 vssd1 vccd1 vccd1 _13182_/C
+ sky130_fd_sc_hd__or4_4
X_10393_ _10275_/A _10275_/B _10391_/Y _10383_/X vssd1 vssd1 vccd1 vccd1 _21360_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_135_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12132_ _20975_/Q vssd1 vssd1 vccd1 vccd1 _12328_/A sky130_fd_sc_hd__inv_2
XFILLER_135_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12063_ _20956_/Q vssd1 vssd1 vccd1 vccd1 _12310_/A sky130_fd_sc_hd__inv_2
X_16940_ _16937_/Y _16938_/X _16939_/X vssd1 vssd1 vccd1 vccd1 _16940_/X sky130_fd_sc_hd__o21a_1
XANTENNA__12711__B1 _11741_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11014_ _20005_/Q vssd1 vssd1 vccd1 vccd1 _11590_/A sky130_fd_sc_hd__buf_1
XFILLER_238_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16871_ _19947_/Q vssd1 vssd1 vccd1 vccd1 _16871_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12798__A _12804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19291__D hold9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18610_ _18609_/X _14903_/Y _18907_/S vssd1 vssd1 vccd1 vccd1 _18610_/X sky130_fd_sc_hd__mux2_1
X_15822_ _19619_/Q _15817_/X _09824_/X _15819_/X vssd1 vssd1 vccd1 vccd1 _19619_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_77_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19590_ _20890_/CLK _19590_/D vssd1 vssd1 vccd1 vccd1 _19590_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18541_ _17938_/Y _20450_/Q _18784_/S vssd1 vssd1 vccd1 vccd1 _18541_/X sky130_fd_sc_hd__mux2_1
X_15753_ _19648_/Q _15750_/X _15701_/X _15751_/X vssd1 vssd1 vccd1 vccd1 _19648_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_92_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12965_ _20703_/Q _12960_/X _12884_/X _12961_/X vssd1 vssd1 vccd1 vccd1 _20703_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_161_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19080__S _19908_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17402__B1 _18829_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14704_ _14723_/A vssd1 vssd1 vccd1 vccd1 _14704_/X sky130_fd_sc_hd__buf_1
X_11916_ _21011_/Q vssd1 vssd1 vccd1 vccd1 _11916_/Y sky130_fd_sc_hd__inv_2
X_18472_ _18845_/A0 _13796_/Y _18896_/S vssd1 vssd1 vccd1 vccd1 _18472_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15684_ _19680_/Q _15681_/X _15588_/X _15682_/X vssd1 vssd1 vccd1 vccd1 _19680_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_33_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12896_ _17085_/A _12899_/A vssd1 vssd1 vccd1 vccd1 _12897_/S sky130_fd_sc_hd__or2_1
XPHY_4460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_29_HCLK_A clkbuf_opt_4_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14635_ _13738_/X _14637_/A _14575_/A vssd1 vssd1 vccd1 vccd1 _14636_/C sky130_fd_sc_hd__o21a_1
XANTENNA__14767__A1 _20132_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17423_ _21216_/Q vssd1 vssd1 vccd1 vccd1 _17423_/Y sky130_fd_sc_hd__inv_2
XPHY_4493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11847_ _11847_/A vssd1 vssd1 vccd1 vccd1 _21032_/D sky130_fd_sc_hd__inv_2
XFILLER_199_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13422__A input43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14566_ _14566_/A _14566_/B vssd1 vssd1 vccd1 vccd1 _14651_/A sky130_fd_sc_hd__or2_2
X_17354_ _19624_/Q vssd1 vssd1 vccd1 vccd1 _17354_/Y sky130_fd_sc_hd__inv_2
X_11778_ _16516_/A vssd1 vssd1 vccd1 vccd1 _16597_/A sky130_fd_sc_hd__buf_1
XFILLER_13_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19250__S0 _20130_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13517_ _20435_/Q _13514_/X _13449_/X _13515_/X vssd1 vssd1 vccd1 vccd1 _20435_/D
+ sky130_fd_sc_hd__a22o_1
X_16305_ _16305_/A vssd1 vssd1 vccd1 vccd1 _16305_/X sky130_fd_sc_hd__buf_1
XFILLER_119_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10729_ _10729_/A _10729_/B _10729_/C vssd1 vssd1 vccd1 vccd1 _21311_/D sky130_fd_sc_hd__nor3_2
X_17285_ _21073_/Q vssd1 vssd1 vccd1 vccd1 _17285_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20416__RESET_B repeater185/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17829__A _18927_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14497_ _14517_/A _14518_/B _14497_/C vssd1 vssd1 vccd1 vccd1 _14515_/A sky130_fd_sc_hd__or3_1
XANTENNA__18424__S _18784_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19024_ _16894_/Y _20399_/Q _19026_/S vssd1 vssd1 vccd1 vccd1 _19952_/D sky130_fd_sc_hd__mux2_1
X_16236_ _19420_/Q _16230_/X _16235_/X _16233_/X vssd1 vssd1 vccd1 vccd1 _19420_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_174_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13448_ _20468_/Q _13444_/X _13446_/X _13447_/X vssd1 vssd1 vccd1 vccd1 _20468_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_174_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_51_HCLK clkbuf_4_11_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _21191_/CLK sky130_fd_sc_hd__clkbuf_16
X_16167_ _16173_/A vssd1 vssd1 vccd1 vccd1 _16174_/A sky130_fd_sc_hd__inv_2
XANTENNA__15349__A input60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13379_ _20501_/Q _13377_/X _13166_/X _13378_/X vssd1 vssd1 vccd1 vccd1 _20501_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15118_ _20435_/Q _15061_/A _15115_/Y _20046_/Q _15117_/X vssd1 vssd1 vccd1 vccd1
+ _15126_/B sky130_fd_sc_hd__a221o_1
X_16098_ _19484_/Q _16094_/X _15869_/X _16096_/X vssd1 vssd1 vccd1 vccd1 _19484_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_114_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15049_ _20053_/Q vssd1 vssd1 vccd1 vccd1 _15068_/B sky130_fd_sc_hd__inv_2
X_19926_ _20841_/CLK _19926_/D repeater256/X vssd1 vssd1 vccd1 vccd1 _19926_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11505__A1 _11504_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21275__RESET_B repeater245/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19857_ _21162_/CLK _19857_/D repeater227/X vssd1 vssd1 vccd1 vccd1 _19857_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_110_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09610_ _20872_/Q _20871_/Q _13383_/A vssd1 vssd1 vccd1 vccd1 _11200_/A sky130_fd_sc_hd__or3_4
X_18808_ _18845_/A0 _10447_/Y _18896_/S vssd1 vssd1 vccd1 vccd1 _18808_/X sky130_fd_sc_hd__mux2_1
XFILLER_228_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19788_ _19789_/CLK _19788_/D vssd1 vssd1 vccd1 vccd1 _19788_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18739_ _18738_/X _19226_/X _18930_/S vssd1 vssd1 vccd1 vccd1 _18739_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20763__CLK _21342_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20701_ _21125_/CLK _20701_/D repeater190/X vssd1 vssd1 vccd1 vccd1 _20701_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_224_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12769__B1 _12668_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13332__A _13357_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20632_ _21481_/CLK _20632_/D repeater206/X vssd1 vssd1 vccd1 vccd1 _20632_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19241__S0 _20132_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20563_ _21357_/CLK _20563_/D repeater198/X vssd1 vssd1 vccd1 vccd1 _20563_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__18334__S _18903_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20494_ _20495_/CLK _20494_/D repeater274/X vssd1 vssd1 vccd1 vccd1 _20494_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_106_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11744__A1 _21056_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12941__B1 _12857_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21115_ _21120_/CLK _21115_/D repeater233/X vssd1 vssd1 vccd1 vccd1 _21115_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17880__B1 _18428_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21046_ _21193_/CLK _21046_/D repeater226/X vssd1 vssd1 vccd1 vccd1 _21046_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17193__B _17193_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09808_ _21455_/Q _09806_/Y _09806_/B _09807_/X vssd1 vssd1 vccd1 vccd1 _21455_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_75_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09739_ _11052_/C vssd1 vssd1 vccd1 vccd1 _09739_/X sky130_fd_sc_hd__buf_1
XANTENNA__18509__S _18897_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12750_ _12750_/A vssd1 vssd1 vccd1 vccd1 _12751_/A sky130_fd_sc_hd__buf_1
XPHY_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20927__RESET_B repeater267/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11701_ _21078_/Q _11697_/X _11684_/X _11699_/X vssd1 vssd1 vccd1 vccd1 _21078_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12681_ _20830_/Q _12679_/X _09630_/X _12680_/X vssd1 vssd1 vccd1 vccd1 _20830_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14420_ _14420_/A _14420_/B _14420_/C _14420_/D vssd1 vssd1 vccd1 vccd1 _14450_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_187_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11632_ _11632_/A _11632_/B vssd1 vssd1 vccd1 vccd1 _11632_/Y sky130_fd_sc_hd__nor2_1
XPHY_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19232__S0 _19275_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09625__B1 _09621_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_74_HCLK clkbuf_4_13_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20697_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14351_ _14351_/A _14351_/B _14518_/C vssd1 vssd1 vccd1 vccd1 _14497_/C sky130_fd_sc_hd__or3_1
XPHY_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11563_ input63/X vssd1 vssd1 vccd1 vccd1 _16335_/A sky130_fd_sc_hd__clkbuf_2
XPHY_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13302_ _13322_/A vssd1 vssd1 vccd1 vccd1 _13302_/X sky130_fd_sc_hd__buf_1
XFILLER_128_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17070_ _20258_/Q _20256_/Q _20257_/Q _17069_/X vssd1 vssd1 vccd1 vccd1 _19887_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_195_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10514_ _21285_/Q _17811_/A _21302_/Q _10513_/Y vssd1 vssd1 vccd1 vccd1 _10514_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_6_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14282_ _20128_/Q vssd1 vssd1 vccd1 vccd1 _15919_/A sky130_fd_sc_hd__buf_1
XPHY_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11494_ _11654_/A _17169_/D vssd1 vssd1 vccd1 vccd1 _14256_/B sky130_fd_sc_hd__or2_2
X_16021_ _16028_/A vssd1 vssd1 vccd1 vccd1 _16021_/X sky130_fd_sc_hd__buf_1
XFILLER_6_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13233_ _13248_/A vssd1 vssd1 vccd1 vccd1 _13233_/X sky130_fd_sc_hd__buf_1
X_10445_ _10761_/A _20673_/Q _21282_/Q _10441_/Y _10444_/X vssd1 vssd1 vccd1 vccd1
+ _10446_/D sky130_fd_sc_hd__o221a_1
XFILLER_124_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13164_ _20603_/Q _13158_/X _13163_/X _13159_/X vssd1 vssd1 vccd1 vccd1 _20603_/D
+ sky130_fd_sc_hd__a22o_1
X_10376_ _10285_/A _10285_/B _10375_/X _10372_/Y vssd1 vssd1 vccd1 vccd1 _21370_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_124_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19075__S _19908_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12115_ _20381_/Q vssd1 vssd1 vccd1 vccd1 _17937_/A sky130_fd_sc_hd__inv_2
XANTENNA__17871__B1 _18559_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17972_ _18210_/X _17931_/X _18300_/X _17932_/X _17971_/X vssd1 vssd1 vccd1 vccd1
+ _17973_/C sky130_fd_sc_hd__o221a_1
X_13095_ _20640_/Q _13092_/X _12954_/X _13093_/X vssd1 vssd1 vccd1 vccd1 _20640_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_78_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19711_ _19776_/CLK _19711_/D vssd1 vssd1 vccd1 vccd1 _19711_/Q sky130_fd_sc_hd__dfxtp_1
X_16923_ _19958_/Q _16913_/A _19959_/Q vssd1 vssd1 vccd1 vccd1 _16923_/X sky130_fd_sc_hd__o21a_1
X_12046_ _12305_/A _20365_/Q _20978_/Q _12045_/Y vssd1 vssd1 vccd1 vccd1 _12046_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_49_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13417__A _13444_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19642_ _20327_/CLK _19642_/D vssd1 vssd1 vccd1 vccd1 _19642_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16854_ _16858_/B _16853_/X _16831_/X vssd1 vssd1 vccd1 vccd1 _16854_/X sky130_fd_sc_hd__o21a_1
XANTENNA__14437__B1 _21477_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15805_ _19627_/Q _15800_/X _09824_/X _15802_/X vssd1 vssd1 vccd1 vccd1 _19627_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_65_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19573_ _19776_/CLK _19573_/D vssd1 vssd1 vccd1 vccd1 _19573_/Q sky130_fd_sc_hd__dfxtp_1
X_16785_ _19927_/Q vssd1 vssd1 vccd1 vccd1 _16785_/Y sky130_fd_sc_hd__inv_2
X_13997_ _20310_/Q _13996_/Y _13988_/A _13887_/B vssd1 vssd1 vccd1 vccd1 _20310_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_80_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18419__S _18903_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15632__A _15632_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18524_ _18523_/X _12284_/Y _18910_/S vssd1 vssd1 vccd1 vccd1 _18524_/X sky130_fd_sc_hd__mux2_1
XANTENNA__20668__RESET_B repeater207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15736_ _15736_/A vssd1 vssd1 vccd1 vccd1 _15736_/X sky130_fd_sc_hd__buf_1
X_12948_ _12960_/A vssd1 vssd1 vccd1 vccd1 _12948_/X sky130_fd_sc_hd__buf_1
XFILLER_234_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09630__A input48/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_221_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11671__B1 _11516_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_153_HCLK_A clkbuf_opt_1_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18455_ _17901_/Y _20787_/Q _18885_/S vssd1 vssd1 vccd1 vccd1 _18455_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15667_ _15667_/A vssd1 vssd1 vccd1 vccd1 _15667_/X sky130_fd_sc_hd__buf_1
X_12879_ _13710_/A vssd1 vssd1 vccd1 vccd1 _12879_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_233_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17406_ _17158_/X _17384_/X _17170_/X _17393_/X _17405_/X vssd1 vssd1 vccd1 vccd1
+ _17406_/Y sky130_fd_sc_hd__o221ai_4
X_14618_ _14585_/A _14585_/B _14607_/X _14616_/Y vssd1 vssd1 vccd1 vccd1 _20196_/D
+ sky130_fd_sc_hd__a211oi_2
X_18386_ _18385_/X _12296_/Y _18910_/S vssd1 vssd1 vccd1 vccd1 _18386_/X sky130_fd_sc_hd__mux2_1
X_15598_ _15604_/A vssd1 vssd1 vccd1 vccd1 _15598_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__19223__S0 _19275_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14549_ _15798_/B _20130_/Q _14747_/B _14548_/X _19121_/X vssd1 vssd1 vccd1 vccd1
+ _14549_/Y sky130_fd_sc_hd__o221ai_1
X_17337_ _19408_/Q vssd1 vssd1 vccd1 vccd1 _17337_/Y sky130_fd_sc_hd__inv_2
XFILLER_186_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18154__S _18896_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12991__A input59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17268_ _19350_/Q vssd1 vssd1 vccd1 vccd1 _17268_/Y sky130_fd_sc_hd__inv_2
XFILLER_128_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19007_ _16968_/X _20416_/Q _19019_/S vssd1 vssd1 vccd1 vccd1 _19969_/D sky130_fd_sc_hd__mux2_1
X_16219_ _19429_/Q _16216_/X _16109_/X _16218_/X vssd1 vssd1 vccd1 vccd1 _19429_/D
+ sky130_fd_sc_hd__a22o_1
X_17199_ _17323_/A vssd1 vssd1 vccd1 vccd1 _17933_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__21456__RESET_B repeater245/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12923__B1 _12922_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19909_ _21338_/CLK _19909_/D repeater221/X vssd1 vssd1 vccd1 vccd1 _19909_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_29_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18329__S _18896_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13100__B1 _12875_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_97_HCLK clkbuf_4_13_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20293_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__17917__B2 _17326_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19214__S0 _19275_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_12_HCLK_A clkbuf_opt_2_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_75_HCLK_A clkbuf_4_13_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20615_ _20622_/CLK _20615_/D repeater195/X vssd1 vssd1 vccd1 vccd1 _20615_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_138_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_rebuffer2_A _20027_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_0_HCLK_A clkbuf_opt_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20546_ _20947_/CLK _20546_/D repeater266/X vssd1 vssd1 vccd1 vccd1 _20546_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_126_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18999__S _19026_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_3_HCLK clkbuf_opt_2_HCLK/A vssd1 vssd1 vccd1 vccd1 _19812_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_153_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20477_ _20480_/CLK _20477_/D repeater183/X vssd1 vssd1 vccd1 vccd1 _20477_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_193_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12914__B1 _12670_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10230_ _21373_/Q vssd1 vssd1 vccd1 vccd1 _10288_/A sky130_fd_sc_hd__inv_2
XFILLER_134_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10161_ _10161_/A _10161_/B vssd1 vssd1 vccd1 vccd1 _10175_/A sky130_fd_sc_hd__or2_2
XFILLER_126_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10092_ _10199_/A _20773_/Q _21376_/Q _10089_/Y _10091_/X vssd1 vssd1 vccd1 vccd1
+ _10098_/C sky130_fd_sc_hd__o221a_1
XFILLER_248_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17605__B1 _11932_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21029_ _21255_/CLK _21029_/D repeater242/X vssd1 vssd1 vccd1 vccd1 _21029_/Q sky130_fd_sc_hd__dfrtp_1
X_13920_ _20641_/Q _20298_/Q _13919_/Y _14014_/A vssd1 vssd1 vccd1 vccd1 _13922_/C
+ sky130_fd_sc_hd__o22a_1
XFILLER_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12141__A _20393_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13851_ _20310_/Q vssd1 vssd1 vccd1 vccd1 _13972_/A sky130_fd_sc_hd__inv_2
XANTENNA__18239__S _18242_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12802_ _20777_/Q _12797_/X _11733_/X _12798_/X vssd1 vssd1 vccd1 vccd1 _20777_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16570_ _21093_/Q _21092_/Q vssd1 vssd1 vccd1 vccd1 _19841_/D sky130_fd_sc_hd__or2_1
XANTENNA__20761__RESET_B repeater205/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13782_ _20609_/Q vssd1 vssd1 vccd1 vccd1 _13782_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10994_ _21019_/Q vssd1 vssd1 vccd1 vccd1 _10994_/X sky130_fd_sc_hd__buf_1
XFILLER_231_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20079__RESET_B repeater259/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15521_ _15588_/A vssd1 vssd1 vccd1 vccd1 _15521_/X sky130_fd_sc_hd__buf_1
X_12733_ _20805_/Q vssd1 vssd1 vccd1 vccd1 _12748_/A sky130_fd_sc_hd__inv_2
XFILLER_43_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18240_ _20864_/Q input14/X _18242_/S vssd1 vssd1 vccd1 vccd1 _18240_/X sky130_fd_sc_hd__mux2_1
X_15452_ _15460_/A vssd1 vssd1 vccd1 vccd1 _15452_/X sky130_fd_sc_hd__buf_1
XANTENNA__20008__RESET_B repeater238/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12664_ _12680_/A vssd1 vssd1 vccd1 vccd1 _12664_/X sky130_fd_sc_hd__buf_1
XANTENNA__19205__S0 _19275_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14403_ _21472_/Q vssd1 vssd1 vccd1 vccd1 _14403_/Y sky130_fd_sc_hd__inv_2
XFILLER_175_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11615_ _21111_/Q _11614_/B _11623_/B _11614_/Y vssd1 vssd1 vccd1 vccd1 _21111_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15383_ _15661_/A vssd1 vssd1 vccd1 vccd1 _15383_/X sky130_fd_sc_hd__buf_1
X_18171_ _18170_/X _10291_/Y _18886_/S vssd1 vssd1 vccd1 vccd1 _18171_/X sky130_fd_sc_hd__mux2_1
XPHY_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12595_ _12601_/A vssd1 vssd1 vccd1 vccd1 _12595_/X sky130_fd_sc_hd__buf_1
XPHY_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14334_ _20230_/Q vssd1 vssd1 vccd1 vccd1 _14460_/A sky130_fd_sc_hd__inv_2
X_17122_ _19486_/Q vssd1 vssd1 vccd1 vccd1 _17122_/Y sky130_fd_sc_hd__inv_2
XPHY_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11546_ _11280_/A _11542_/Y _12504_/B _12501_/B _11545_/X vssd1 vssd1 vccd1 vccd1
+ _16569_/D sky130_fd_sc_hd__a2111o_1
XPHY_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_183_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17053_ _19851_/D vssd1 vssd1 vccd1 vccd1 _17058_/C sky130_fd_sc_hd__inv_2
XFILLER_184_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14265_ _20249_/Q _14257_/X _14264_/X _14260_/X vssd1 vssd1 vccd1 vccd1 _20249_/D
+ sky130_fd_sc_hd__a22o_1
X_11477_ _19100_/X _11474_/X _21158_/Q _11475_/X vssd1 vssd1 vccd1 vccd1 _21158_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_183_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16004_ _19532_/Q _16000_/X _15973_/X _16002_/X vssd1 vssd1 vccd1 vccd1 _19532_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_7_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13216_ input48/X vssd1 vssd1 vccd1 vccd1 _13216_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__12905__B1 _12651_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10428_ _20684_/Q vssd1 vssd1 vccd1 vccd1 _10428_/Y sky130_fd_sc_hd__inv_2
X_14196_ _20280_/Q _14195_/Y _14183_/X _14091_/B vssd1 vssd1 vccd1 vccd1 _20280_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_124_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13147_ _20612_/Q _13139_/X _13146_/X _13142_/X vssd1 vssd1 vccd1 vccd1 _20612_/D
+ sky130_fd_sc_hd__a22o_1
X_10359_ _10261_/A _20704_/Q _21360_/Q _10355_/Y _10358_/X vssd1 vssd1 vccd1 vccd1
+ _10360_/D sky130_fd_sc_hd__o221a_1
XANTENNA__14531__A _15832_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19944__RESET_B repeater251/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17955_ _17955_/A vssd1 vssd1 vccd1 vccd1 _17955_/X sky130_fd_sc_hd__buf_1
X_13078_ _13078_/A vssd1 vssd1 vccd1 vccd1 _13098_/A sky130_fd_sc_hd__buf_1
XFILLER_39_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_239_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12029_ _12029_/A vssd1 vssd1 vccd1 vccd1 _12029_/X sky130_fd_sc_hd__buf_1
X_16906_ _16906_/A _16906_/B vssd1 vssd1 vccd1 vccd1 _16906_/Y sky130_fd_sc_hd__nor2_1
XFILLER_39_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17886_ _09719_/Y _17853_/X _10956_/Y _17854_/X vssd1 vssd1 vccd1 vccd1 _17886_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19625_ _21449_/CLK _19625_/D vssd1 vssd1 vccd1 vccd1 _19625_/Q sky130_fd_sc_hd__dfxtp_1
X_16837_ _16834_/A _16829_/A _16836_/Y vssd1 vssd1 vccd1 vccd1 _16838_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__18149__S _18904_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19556_ _19776_/CLK _19556_/D vssd1 vssd1 vccd1 vccd1 _19556_/Q sky130_fd_sc_hd__dfxtp_1
X_16768_ _19923_/Q vssd1 vssd1 vccd1 vccd1 _16770_/A sky130_fd_sc_hd__inv_2
XFILLER_19_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_202_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18507_ _18506_/X _10275_/A _18886_/S vssd1 vssd1 vccd1 vccd1 _18507_/X sky130_fd_sc_hd__mux2_1
XFILLER_179_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15719_ _19664_/Q _15716_/X _15701_/X _15717_/X vssd1 vssd1 vccd1 vccd1 _19664_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__20431__RESET_B repeater235/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19487_ _20890_/CLK _19487_/D vssd1 vssd1 vccd1 vccd1 _19487_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_221_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16699_ _19894_/Q _14234_/B _14235_/B vssd1 vssd1 vccd1 vccd1 _16699_/X sky130_fd_sc_hd__a21bo_1
XFILLER_22_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18438_ _18848_/A0 _17876_/Y _18666_/S vssd1 vssd1 vccd1 vccd1 _18438_/X sky130_fd_sc_hd__mux2_1
XFILLER_221_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13397__B1 _13274_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_221_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17289__A _21081_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18369_ _17982_/Y _20793_/Q _18885_/S vssd1 vssd1 vccd1 vccd1 _18369_/X sky130_fd_sc_hd__mux2_1
XFILLER_187_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20400_ _21234_/CLK _20400_/D repeater270/X vssd1 vssd1 vccd1 vccd1 _20400_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_108_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21380_ _21421_/CLK _21380_/D repeater214/X vssd1 vssd1 vccd1 vccd1 _21380_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__13149__B1 _13148_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20331_ _20331_/CLK _20331_/D repeater190/X vssd1 vssd1 vccd1 vccd1 _20331_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_134_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18612__S _18680_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__21290__RESET_B repeater210/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20262_ _20724_/CLK _20262_/D repeater264/X vssd1 vssd1 vccd1 vccd1 _20262_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_143_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20193_ _20626_/CLK _20193_/D repeater200/X vssd1 vssd1 vccd1 vccd1 _20193_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_115_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10438__B2 _20690_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20172__RESET_B repeater248/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20101__RESET_B repeater259/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11400_ _11402_/B vssd1 vssd1 vccd1 vccd1 _11421_/A sky130_fd_sc_hd__buf_1
XFILLER_21_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12380_ _12380_/A vssd1 vssd1 vccd1 vccd1 _12380_/Y sky130_fd_sc_hd__inv_2
XFILLER_166_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11331_ _21179_/Q vssd1 vssd1 vccd1 vccd1 _11363_/A sky130_fd_sc_hd__buf_1
XFILLER_166_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20529_ _20944_/CLK _20529_/D repeater274/X vssd1 vssd1 vccd1 vccd1 _20529_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__17927__A _18020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18522__S _18908_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14888__B1 _20594_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14050_ _20278_/Q vssd1 vssd1 vccd1 vccd1 _14088_/A sky130_fd_sc_hd__inv_2
X_11262_ _20909_/Q vssd1 vssd1 vccd1 vccd1 _11313_/B sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_104_HCLK clkbuf_4_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20590_/CLK sky130_fd_sc_hd__clkbuf_16
X_13001_ input55/X vssd1 vssd1 vccd1 vccd1 _13001_/X sky130_fd_sc_hd__buf_2
XANTENNA__17826__B1 _18289_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10213_ _10213_/A vssd1 vssd1 vccd1 vccd1 _10213_/Y sky130_fd_sc_hd__inv_2
XFILLER_134_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11193_ _11193_/A vssd1 vssd1 vccd1 vccd1 _11193_/X sky130_fd_sc_hd__buf_1
XFILLER_239_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input42_A HWDATA[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10144_ _20736_/Q _10185_/A vssd1 vssd1 vccd1 vccd1 _10145_/A sky130_fd_sc_hd__or2_1
XFILLER_239_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13312__B1 _13311_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17740_ _19701_/Q vssd1 vssd1 vccd1 vccd1 _17740_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20942__RESET_B repeater278/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14952_ _14978_/A vssd1 vssd1 vccd1 vccd1 _14952_/X sky130_fd_sc_hd__buf_1
X_10075_ _10148_/B _10075_/B _10075_/C vssd1 vssd1 vccd1 vccd1 _10168_/A sky130_fd_sc_hd__or3_1
XFILLER_87_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18251__A0 _18250_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13903_ _20645_/Q vssd1 vssd1 vccd1 vccd1 _13903_/Y sky130_fd_sc_hd__inv_2
X_17671_ _19428_/Q vssd1 vssd1 vccd1 vccd1 _17671_/Y sky130_fd_sc_hd__inv_2
X_14883_ _14883_/A _14883_/B vssd1 vssd1 vccd1 vccd1 _14884_/A sky130_fd_sc_hd__or2_1
XANTENNA_output129_A _21103_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19410_ _21001_/CLK _19410_/D vssd1 vssd1 vccd1 vccd1 _19410_/Q sky130_fd_sc_hd__dfxtp_1
X_16622_ _16508_/A _16621_/Y _16501_/X _11748_/B _16494_/X vssd1 vssd1 vccd1 vccd1
+ _16623_/A sky130_fd_sc_hd__o32a_1
XFILLER_35_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13834_ _20630_/Q _13832_/Y _20623_/Q _14589_/A vssd1 vssd1 vccd1 vccd1 _13834_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_62_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19341_ _19961_/CLK _19341_/D vssd1 vssd1 vccd1 vccd1 _19341_/Q sky130_fd_sc_hd__dfxtp_1
X_16553_ _16553_/A _16584_/B vssd1 vssd1 vccd1 vccd1 _16566_/C sky130_fd_sc_hd__or2_2
X_13765_ _20189_/Q vssd1 vssd1 vccd1 vccd1 _14578_/A sky130_fd_sc_hd__inv_2
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12969__A3 _10985_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10977_ _20868_/Q _20867_/Q vssd1 vssd1 vccd1 vccd1 _15884_/A sky130_fd_sc_hd__or2_4
XFILLER_203_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15504_ _19766_/Q _15499_/X _15431_/X _15500_/X vssd1 vssd1 vccd1 vccd1 _19766_/D
+ sky130_fd_sc_hd__a22o_1
X_12716_ _17639_/A _12716_/B _12716_/C _20875_/Q vssd1 vssd1 vccd1 vccd1 _13104_/B
+ sky130_fd_sc_hd__or4b_4
X_19272_ _17093_/Y _17094_/Y _17095_/Y _17096_/Y _19275_/S0 _21004_/Q vssd1 vssd1
+ vccd1 vccd1 _19272_/X sky130_fd_sc_hd__mux4_2
XFILLER_231_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16484_ _16484_/A _16484_/B vssd1 vssd1 vccd1 vccd1 _16484_/Y sky130_fd_sc_hd__nor2_1
X_13696_ _20342_/Q _13693_/X _12863_/A _13694_/X vssd1 vssd1 vccd1 vccd1 _20342_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_31_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13379__B1 _13166_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_231_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18223_ _20847_/Q input27/X _18236_/S vssd1 vssd1 vccd1 vccd1 _18223_/X sky130_fd_sc_hd__mux2_4
XPHY_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15435_ _15441_/A vssd1 vssd1 vccd1 vccd1 _15442_/A sky130_fd_sc_hd__inv_2
X_12647_ _13328_/A _17323_/A vssd1 vssd1 vccd1 vccd1 _12815_/A sky130_fd_sc_hd__or2_2
XFILLER_31_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14526__A _20208_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13430__A _13447_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18154_ _18845_/A0 _10472_/Y _18896_/S vssd1 vssd1 vccd1 vccd1 _18154_/X sky130_fd_sc_hd__mux2_1
X_15366_ _15366_/A vssd1 vssd1 vccd1 vccd1 _15366_/X sky130_fd_sc_hd__buf_1
XANTENNA__16317__B1 _16237_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12578_ _20886_/Q _12574_/X _18238_/X _12575_/X vssd1 vssd1 vccd1 vccd1 _20886_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17105_ _19710_/Q vssd1 vssd1 vccd1 vccd1 _17105_/Y sky130_fd_sc_hd__inv_2
X_11529_ _11535_/A vssd1 vssd1 vccd1 vccd1 _11529_/X sky130_fd_sc_hd__buf_1
X_14317_ _16451_/B _15490_/A vssd1 vssd1 vccd1 vccd1 _14318_/A sky130_fd_sc_hd__or2_1
XFILLER_8_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15297_ _19863_/Q _15297_/B vssd1 vssd1 vccd1 vccd1 _15298_/B sky130_fd_sc_hd__or2_1
XFILLER_156_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18085_ _20426_/Q _18085_/B vssd1 vssd1 vccd1 vccd1 _18085_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__18432__S _18906_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14248_ _20257_/Q _14246_/X _20256_/Q _18946_/S vssd1 vssd1 vccd1 vccd1 _20257_/D
+ sky130_fd_sc_hd__a22o_1
X_17036_ _17036_/A _17038_/B vssd1 vssd1 vccd1 vccd1 _20020_/D sky130_fd_sc_hd__nor2_1
X_14179_ _14179_/A vssd1 vssd1 vccd1 vccd1 _14179_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19377__CLK _19706_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18490__A0 _17079_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18987_ _21266_/Q _21118_/Q _18992_/S vssd1 vssd1 vccd1 vccd1 _18987_/X sky130_fd_sc_hd__mux2_1
XFILLER_239_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13303__B1 _13140_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17572__A _18748_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20683__RESET_B repeater208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17938_ _17938_/A _17938_/B vssd1 vssd1 vccd1 vccd1 _17938_/Y sky130_fd_sc_hd__nor2_1
XFILLER_227_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater146 _19026_/S vssd1 vssd1 vccd1 vccd1 _19019_/S sky130_fd_sc_hd__buf_8
Xrepeater157 _18886_/S vssd1 vssd1 vccd1 vccd1 _18667_/S sky130_fd_sc_hd__buf_8
Xrepeater168 _18874_/S vssd1 vssd1 vccd1 vccd1 _18909_/S sky130_fd_sc_hd__buf_8
X_17869_ _17869_/A vssd1 vssd1 vccd1 vccd1 _17869_/X sky130_fd_sc_hd__buf_1
Xrepeater179 _18242_/S vssd1 vssd1 vccd1 vccd1 _18236_/S sky130_fd_sc_hd__buf_8
XFILLER_227_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19608_ _20890_/CLK _19608_/D vssd1 vssd1 vccd1 vccd1 _19608_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13605__A _13625_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20880_ _21459_/CLK _20880_/D repeater243/X vssd1 vssd1 vccd1 vccd1 _20880_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_226_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19539_ _21462_/CLK _19539_/D vssd1 vssd1 vccd1 vccd1 _19539_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18607__S _18928_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11125__A _21004_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_195_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21471__RESET_B repeater204/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21432_ _21438_/CLK _21432_/D repeater236/X vssd1 vssd1 vccd1 vccd1 _21432_/Q sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_127_HCLK clkbuf_4_4_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20422_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__17169__D _17169_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21363_ _21367_/CLK _21363_/D repeater254/X vssd1 vssd1 vccd1 vccd1 _21363_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_175_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18342__S _18908_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19866__RESET_B repeater217/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20314_ _20316_/CLK _20314_/D repeater197/X vssd1 vssd1 vccd1 vccd1 _20314_/Q sky130_fd_sc_hd__dfrtp_1
X_21294_ _21294_/CLK _21294_/D repeater209/X vssd1 vssd1 vccd1 vccd1 _21294_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_190_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11795__A _11795_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13542__B1 _13538_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20245_ _21421_/CLK _20245_/D repeater214/X vssd1 vssd1 vccd1 vccd1 _20245_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18481__A0 _18848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20176_ _21485_/CLK _20176_/D repeater200/X vssd1 vssd1 vccd1 vccd1 _20176_/Q sky130_fd_sc_hd__dfrtp_4
X_09987_ _09987_/A vssd1 vssd1 vccd1 vccd1 _09988_/B sky130_fd_sc_hd__inv_2
XFILLER_76_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17587__A2 _17559_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10900_ _11743_/A vssd1 vssd1 vccd1 vccd1 _10900_/X sky130_fd_sc_hd__buf_2
XFILLER_245_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11880_ _11878_/Y _10983_/A _21021_/Q _11883_/A vssd1 vssd1 vccd1 vccd1 _11881_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_123_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10858__B _20887_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10831_ _21284_/Q _10829_/Y _10830_/X _10762_/B vssd1 vssd1 vccd1 vccd1 _21284_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_16_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18517__S _18617_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15730__A _16235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13550_ input57/X vssd1 vssd1 vccd1 vccd1 _13550_/X sky130_fd_sc_hd__buf_4
XFILLER_213_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10762_ _10762_/A _10762_/B vssd1 vssd1 vccd1 vccd1 _10825_/A sky130_fd_sc_hd__or2_2
XFILLER_197_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12501_ _16568_/B _12501_/B _16569_/C vssd1 vssd1 vccd1 vccd1 _12525_/B sky130_fd_sc_hd__or3_4
XFILLER_200_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13481_ _13481_/A vssd1 vssd1 vccd1 vccd1 _13481_/X sky130_fd_sc_hd__buf_1
X_10693_ _10693_/A vssd1 vssd1 vccd1 vccd1 _10693_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15220_ _18078_/A _15029_/A _20474_/Q _15068_/B _15219_/X vssd1 vssd1 vccd1 vccd1
+ _15232_/A sky130_fd_sc_hd__o221a_1
X_12432_ _12432_/A _12443_/A _12432_/C vssd1 vssd1 vccd1 vccd1 _12440_/A sky130_fd_sc_hd__or3_4
XFILLER_200_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15151_ _20449_/Q vssd1 vssd1 vccd1 vccd1 _15151_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12363_ _20967_/Q _12362_/Y _12359_/X _12321_/B vssd1 vssd1 vccd1 vccd1 _20967_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__18252__S _18680_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14102_ _20561_/Q vssd1 vssd1 vccd1 vccd1 _14102_/Y sky130_fd_sc_hd__inv_2
X_11314_ _12500_/B _12502_/B _11314_/C _12504_/B vssd1 vssd1 vccd1 vccd1 _11317_/C
+ sky130_fd_sc_hd__or4_4
X_15082_ _15104_/A _15082_/B vssd1 vssd1 vccd1 vccd1 _15173_/A sky130_fd_sc_hd__or2_1
X_12294_ _20947_/Q _12289_/Y _20920_/Q _12290_/Y _12293_/X vssd1 vssd1 vccd1 vccd1
+ _12301_/C sky130_fd_sc_hd__o221a_1
X_18910_ _18909_/X _17172_/Y _18910_/S vssd1 vssd1 vccd1 vccd1 _18910_/X sky130_fd_sc_hd__mux2_1
X_14033_ _14033_/A _14033_/B _14037_/C vssd1 vssd1 vccd1 vccd1 _20294_/D sky130_fd_sc_hd__nor3_1
X_11245_ _11251_/A vssd1 vssd1 vccd1 vccd1 _11245_/X sky130_fd_sc_hd__buf_1
XFILLER_4_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19890_ _21141_/CLK _19890_/D repeater192/X vssd1 vssd1 vccd1 vccd1 _19890_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_122_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18472__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18841_ _18840_/X _10261_/A _18841_/S vssd1 vssd1 vccd1 vccd1 _18841_/X sky130_fd_sc_hd__mux2_1
X_11176_ _11176_/A _11176_/B vssd1 vssd1 vccd1 vccd1 _11176_/Y sky130_fd_sc_hd__nor2_1
XFILLER_121_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15286__B1 _20043_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10127_ _10151_/A _20787_/Q _10056_/A _20787_/Q vssd1 vssd1 vccd1 vccd1 _10127_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_18772_ _18771_/X _17450_/Y _18879_/S vssd1 vssd1 vccd1 vccd1 _18772_/X sky130_fd_sc_hd__mux2_1
X_15984_ _16451_/B vssd1 vssd1 vccd1 vccd1 _16229_/B sky130_fd_sc_hd__buf_1
XFILLER_209_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17723_ _17721_/Y _17639_/X _17722_/Y _17162_/B vssd1 vssd1 vccd1 vccd1 _17723_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_57_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14935_ _20576_/Q _20087_/Q _14934_/Y _14863_/C vssd1 vssd1 vccd1 vccd1 _14935_/X
+ sky130_fd_sc_hd__o22a_1
X_10058_ _21396_/Q vssd1 vssd1 vccd1 vccd1 _10059_/A sky130_fd_sc_hd__inv_2
XFILLER_209_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18000__B _18001_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17654_ _17650_/Y _17376_/A _17651_/Y _17150_/X _17653_/X vssd1 vssd1 vccd1 vccd1
+ _17654_/X sky130_fd_sc_hd__o221a_1
X_14866_ _14960_/D _14866_/B vssd1 vssd1 vccd1 vccd1 _14994_/A sky130_fd_sc_hd__or2_1
XFILLER_35_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16605_ _16541_/A _16546_/A _16537_/Y _16604_/X vssd1 vssd1 vccd1 vccd1 _16605_/X
+ sky130_fd_sc_hd__o31a_1
X_13817_ _20603_/Q _14570_/A _13813_/Y _20179_/Q _13816_/X vssd1 vssd1 vccd1 vccd1
+ _13836_/A sky130_fd_sc_hd__o221a_1
XFILLER_63_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17585_ _12605_/A _17579_/X _17582_/Y _17584_/X vssd1 vssd1 vccd1 vccd1 _17585_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__14261__A1 _16720_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14797_ _14797_/A vssd1 vssd1 vccd1 vccd1 _19125_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__18427__S _18835_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19991__SET_B repeater220/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19324_ _19626_/CLK _19324_/D vssd1 vssd1 vccd1 vccd1 _19324_/Q sky130_fd_sc_hd__dfxtp_1
X_16536_ _19993_/Q vssd1 vssd1 vccd1 vccd1 _16737_/A sky130_fd_sc_hd__buf_1
XFILLER_50_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13748_ _20617_/Q _14583_/A _13744_/Y _20199_/Q _13747_/X vssd1 vssd1 vccd1 vccd1
+ _13761_/B sky130_fd_sc_hd__o221a_1
XANTENNA_clkbuf_opt_3_HCLK_A clkbuf_opt_3_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21229__RESET_B repeater249/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19255_ _17342_/Y _17343_/Y _17344_/Y _17345_/Y _19275_/S0 _21004_/Q vssd1 vssd1
+ vccd1 vccd1 _19255_/X sky130_fd_sc_hd__mux4_2
XFILLER_149_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16467_ _16473_/A vssd1 vssd1 vccd1 vccd1 _16474_/A sky130_fd_sc_hd__inv_2
X_13679_ _13679_/A vssd1 vssd1 vccd1 vccd1 _13679_/X sky130_fd_sc_hd__buf_1
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18206_ _18205_/X _15097_/Y _18784_/S vssd1 vssd1 vccd1 vccd1 _18206_/X sky130_fd_sc_hd__mux2_1
X_15418_ _19805_/Q _15415_/X _15378_/X _15417_/X vssd1 vssd1 vccd1 vccd1 _19805_/D
+ sky130_fd_sc_hd__a22o_1
X_19186_ _19182_/X _19183_/X _19184_/X _19185_/X _20123_/Q _20124_/Q vssd1 vssd1 vccd1
+ vccd1 _19186_/X sky130_fd_sc_hd__mux4_2
X_16398_ _19337_/Q _16392_/X _16332_/X _16394_/X vssd1 vssd1 vccd1 vccd1 _19337_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_157_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18137_ _18136_/X _12183_/Y _18787_/S vssd1 vssd1 vccd1 vccd1 _18137_/X sky130_fd_sc_hd__mux2_2
XFILLER_117_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15349_ input60/X vssd1 vssd1 vccd1 vccd1 _15588_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__18162__S _18748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18068_ _18018_/X _18068_/B _18068_/C vssd1 vssd1 vccd1 vccd1 _18068_/Y sky130_fd_sc_hd__nand3b_4
XFILLER_132_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09910_ _21253_/Q _17020_/A _09907_/Y _09908_/Y _09909_/Y vssd1 vssd1 vccd1 vccd1
+ _09910_/X sky130_fd_sc_hd__o221a_1
X_17019_ _17019_/A vssd1 vssd1 vccd1 vccd1 _17023_/B sky130_fd_sc_hd__buf_1
XFILLER_208_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09841_ _20033_/Q vssd1 vssd1 vccd1 vccd1 _09861_/B sky130_fd_sc_hd__inv_2
X_20030_ _21357_/CLK _20030_/D repeater199/X vssd1 vssd1 vccd1 vccd1 _20030_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_101_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09772_ _09777_/B vssd1 vssd1 vccd1 vccd1 _09781_/B sky130_fd_sc_hd__buf_1
XFILLER_140_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_246_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09813__A _09827_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18766__A1 _19236_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20932_ _20943_/CLK _20932_/D repeater275/X vssd1 vssd1 vccd1 vccd1 _20932_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_4119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_240_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20863_ _21444_/CLK _20863_/D repeater246/X vssd1 vssd1 vccd1 vccd1 _20863_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_242_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18337__S _18897_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_230_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15550__A _15663_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20794_ _21407_/CLK _20794_/D repeater252/X vssd1 vssd1 vccd1 vccd1 _20794_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12893__B _12899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21415_ _21419_/CLK _21415_/D repeater232/X vssd1 vssd1 vccd1 vccd1 _21415_/Q sky130_fd_sc_hd__dfrtp_1
X_21346_ _21349_/CLK _21346_/D repeater210/X vssd1 vssd1 vccd1 vccd1 _21346_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_2_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21277_ _21306_/CLK _21277_/D repeater205/X vssd1 vssd1 vccd1 vccd1 _21277_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_118_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18800__S _18930_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11030_ _19956_/Q _16905_/A vssd1 vssd1 vccd1 vccd1 _16909_/A sky130_fd_sc_hd__or2_1
X_20228_ _21485_/CLK _20228_/D repeater200/X vssd1 vssd1 vccd1 vccd1 _20228_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__15725__A _16231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20159_ _20159_/CLK _20159_/D repeater189/X vssd1 vssd1 vccd1 vccd1 _20159_/Q sky130_fd_sc_hd__dfrtp_1
X_12981_ _12981_/A _13261_/A vssd1 vssd1 vccd1 vccd1 _13018_/A sky130_fd_sc_hd__or2_2
X_14720_ _20150_/Q _14717_/X _14262_/X _14718_/X vssd1 vssd1 vccd1 vccd1 _20150_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13245__A _14264_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11932_ _21008_/Q vssd1 vssd1 vccd1 vccd1 _11932_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_150_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14651_ _14651_/A vssd1 vssd1 vccd1 vccd1 _14651_/Y sky130_fd_sc_hd__inv_2
X_11863_ _11863_/A vssd1 vssd1 vccd1 vccd1 _11863_/X sky130_fd_sc_hd__buf_1
XANTENNA__15440__B1 _15421_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10814_ _10769_/A _10769_/B _10809_/X _10811_/Y vssd1 vssd1 vccd1 vccd1 _21293_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_60_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13602_ _13600_/X _20396_/Q _13602_/S vssd1 vssd1 vccd1 vccd1 _20396_/D sky130_fd_sc_hd__mux2_1
XPHY_3952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17370_ _17370_/A vssd1 vssd1 vccd1 vccd1 _17536_/A sky130_fd_sc_hd__buf_1
XPHY_3963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14582_ _14582_/A _14623_/A vssd1 vssd1 vccd1 vccd1 _14583_/B sky130_fd_sc_hd__or2_2
X_11794_ _11794_/A vssd1 vssd1 vccd1 vccd1 _11795_/A sky130_fd_sc_hd__inv_2
XFILLER_198_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16321_ _19377_/Q _16319_/X _16009_/X _16320_/X vssd1 vssd1 vccd1 vccd1 _19377_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10745_ _19939_/Q _19938_/Q _19940_/Q vssd1 vssd1 vccd1 vccd1 _16843_/A sky130_fd_sc_hd__or3_1
X_13533_ _16525_/A _11974_/X _13520_/Y vssd1 vssd1 vccd1 vccd1 _13533_/X sky130_fd_sc_hd__o21a_1
XFILLER_43_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19040_ _16825_/X _20829_/Q _19046_/S vssd1 vssd1 vccd1 vccd1 _19936_/D sky130_fd_sc_hd__mux2_1
X_13464_ _20462_/Q _13458_/X _13272_/X _13461_/X vssd1 vssd1 vccd1 vccd1 _20462_/D
+ sky130_fd_sc_hd__a22o_1
X_16252_ _19412_/Q _16248_/X _16113_/X _16250_/X vssd1 vssd1 vccd1 vccd1 _19412_/D
+ sky130_fd_sc_hd__a22o_1
X_10676_ _10664_/A _10675_/A _21335_/Q _10675_/Y _10642_/X vssd1 vssd1 vccd1 vccd1
+ _21335_/D sky130_fd_sc_hd__o221a_1
XFILLER_9_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19078__S _19908_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15203_ _15068_/B _15202_/A _15092_/X _15202_/Y _15160_/X vssd1 vssd1 vccd1 vccd1
+ _20053_/D sky130_fd_sc_hd__o221a_1
X_12415_ _12415_/A vssd1 vssd1 vccd1 vccd1 _12436_/B sky130_fd_sc_hd__inv_2
XFILLER_139_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16183_ _19445_/Q _16180_/X _16131_/X _16182_/X vssd1 vssd1 vccd1 vccd1 _19445_/D
+ sky130_fd_sc_hd__a22o_1
X_13395_ _20495_/Q _13390_/X _13270_/X _13393_/X vssd1 vssd1 vccd1 vccd1 _20495_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_127_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12346_ _12329_/A _12329_/B _12376_/A _12342_/Y vssd1 vssd1 vccd1 vccd1 _20976_/D
+ sky130_fd_sc_hd__a211oi_2
X_15134_ _20456_/Q _15081_/A _15133_/Y _20056_/Q vssd1 vssd1 vccd1 vccd1 _15134_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_153_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15065_ _15065_/A _15065_/B vssd1 vssd1 vccd1 vccd1 _15205_/A sky130_fd_sc_hd__or2_1
XFILLER_4_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19942_ _21372_/CLK _19942_/D repeater251/X vssd1 vssd1 vccd1 vccd1 _19942_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_126_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12277_ _20943_/Q _12273_/Y _20932_/Q _12274_/Y _12276_/X vssd1 vssd1 vccd1 vccd1
+ _12278_/D sky130_fd_sc_hd__o221a_1
XANTENNA__09617__B _12898_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18710__S _18875_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14016_ _14016_/A _14020_/A vssd1 vssd1 vccd1 vccd1 _14017_/B sky130_fd_sc_hd__or2_2
X_11228_ _21199_/Q _11225_/X _10896_/X _11226_/X vssd1 vssd1 vccd1 vccd1 _21199_/D
+ sky130_fd_sc_hd__a22o_1
X_19873_ _21164_/CLK _19873_/D repeater225/X vssd1 vssd1 vccd1 vccd1 _19873_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17834__B _18929_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18824_ _17371_/X _21252_/Q _20870_/Q vssd1 vssd1 vccd1 vccd1 _18824_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11159_ _20432_/Q vssd1 vssd1 vccd1 vccd1 _11160_/D sky130_fd_sc_hd__inv_2
XFILLER_228_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09633__A input47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18755_ _17537_/Y _10003_/Y _20870_/Q vssd1 vssd1 vccd1 vccd1 _18755_/X sky130_fd_sc_hd__mux2_1
X_15967_ _15985_/A _15967_/B _16451_/C vssd1 vssd1 vccd1 vccd1 _15978_/A sky130_fd_sc_hd__or3_4
XFILLER_48_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17706_ _17777_/A _20115_/Q vssd1 vssd1 vccd1 vccd1 _17706_/Y sky130_fd_sc_hd__nand2_1
XFILLER_209_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14918_ _14918_/A _14918_/B _14918_/C _14918_/D vssd1 vssd1 vccd1 vccd1 _14949_/B
+ sky130_fd_sc_hd__and4_1
X_18686_ _18845_/A0 _10466_/Y _18896_/S vssd1 vssd1 vccd1 vccd1 _18686_/X sky130_fd_sc_hd__mux2_1
XFILLER_63_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_236_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15898_ _19585_/Q _15896_/X _15788_/X _15897_/X vssd1 vssd1 vccd1 vccd1 _19585_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_236_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17637_ _21061_/Q vssd1 vssd1 vccd1 vccd1 _17637_/Y sky130_fd_sc_hd__inv_2
XFILLER_224_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14849_ _20080_/Q vssd1 vssd1 vccd1 vccd1 _15000_/A sky130_fd_sc_hd__inv_2
XANTENNA__16466__A _16473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18157__S _18775_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_212_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17568_ _16550_/Y _17550_/X _17561_/Y _17376_/X _17567_/X vssd1 vssd1 vccd1 vccd1
+ _17568_/X sky130_fd_sc_hd__o221a_2
XANTENNA__19565__CLK _19706_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19307_ _20241_/CLK _19307_/D vssd1 vssd1 vccd1 vccd1 _19307_/Q sky130_fd_sc_hd__dfxtp_1
X_16519_ _21094_/Q vssd1 vssd1 vccd1 vccd1 _16519_/Y sky130_fd_sc_hd__inv_2
XFILLER_189_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17499_ _19402_/Q vssd1 vssd1 vccd1 vccd1 _17499_/Y sky130_fd_sc_hd__inv_2
XFILLER_210_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_220_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19238_ _17432_/Y _17433_/Y _17434_/Y _17435_/Y _20130_/Q _20131_/Q vssd1 vssd1 vccd1
+ vccd1 _19238_/X sky130_fd_sc_hd__mux4_2
XFILLER_164_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19169_ _19727_/Q _19367_/Q _19783_/Q _19767_/Q _19280_/S0 _20122_/Q vssd1 vssd1
+ vccd1 vccd1 _19169_/X sky130_fd_sc_hd__mux4_2
XFILLER_145_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21200_ _21255_/CLK _21200_/D repeater240/X vssd1 vssd1 vccd1 vccd1 _21200_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_172_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15498__B1 _15421_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21131_ _21134_/CLK _21131_/D repeater192/X vssd1 vssd1 vccd1 vccd1 _21131_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18620__S _18896_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21062_ _21134_/CLK _21062_/D repeater227/X vssd1 vssd1 vccd1 vccd1 _21062_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20013_ _21438_/CLK _20013_/D repeater236/X vssd1 vssd1 vccd1 vccd1 _20013_/Q sky130_fd_sc_hd__dfrtp_1
X_09824_ _15871_/A vssd1 vssd1 vccd1 vccd1 _09824_/X sky130_fd_sc_hd__buf_1
XANTENNA__12888__B _12899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09755_ _11052_/D _20147_/Q _11062_/A _20157_/Q _09754_/X vssd1 vssd1 vccd1 vccd1
+ _09768_/B sky130_fd_sc_hd__o221a_1
XANTENNA__18739__A1 _19226_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15670__B1 _15590_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_227_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09686_ _21467_/Q _09673_/X _09685_/X _09678_/X vssd1 vssd1 vccd1 vccd1 _21467_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_55_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20915_ _20915_/CLK _20915_/D repeater218/X vssd1 vssd1 vccd1 vccd1 _20915_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_199_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15422__B1 _15421_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20846_ _20857_/CLK _20846_/D repeater243/X vssd1 vssd1 vccd1 vccd1 _20846_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_120_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20777_ _21147_/CLK _20777_/D repeater215/X vssd1 vssd1 vccd1 vccd1 _20777_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10530_ _20699_/Q vssd1 vssd1 vccd1 vccd1 _10722_/A sky130_fd_sc_hd__inv_2
XPHY_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10461_ _20694_/Q vssd1 vssd1 vccd1 vccd1 _10461_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12200_ _12081_/X _20342_/Q _12105_/X _20352_/Q _12199_/X vssd1 vssd1 vccd1 vccd1
+ _12204_/C sky130_fd_sc_hd__o221a_1
XFILLER_109_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13180_ _13180_/A vssd1 vssd1 vccd1 vccd1 _13528_/A sky130_fd_sc_hd__buf_1
XFILLER_202_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10392_ _21361_/Q _10391_/Y _10277_/B _10381_/X vssd1 vssd1 vccd1 vccd1 _21361_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__20715__RESET_B repeater254/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12131_ _20389_/Q vssd1 vssd1 vccd1 vccd1 _12131_/Y sky130_fd_sc_hd__inv_2
XFILLER_123_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21329_ _21477_/CLK _21329_/D repeater204/X vssd1 vssd1 vccd1 vccd1 _21329_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_150_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18530__S _18644_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18427__A0 _17281_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12062_ _20377_/Q vssd1 vssd1 vccd1 vccd1 _12062_/Y sky130_fd_sc_hd__inv_2
XFILLER_238_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11013_ _19108_/X _19115_/S _10985_/Y _11012_/X vssd1 vssd1 vccd1 vccd1 _21245_/D
+ sky130_fd_sc_hd__a22oi_1
X_16870_ _16877_/A _16870_/B vssd1 vssd1 vccd1 vccd1 _16870_/Y sky130_fd_sc_hd__nor2_1
XFILLER_238_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15821_ _19620_/Q _15817_/X _09821_/X _15819_/X vssd1 vssd1 vccd1 vccd1 _19620_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_46_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18540_ _18539_/X _16951_/A _18680_/S vssd1 vssd1 vccd1 vccd1 _18540_/X sky130_fd_sc_hd__mux2_2
XFILLER_58_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15752_ _19649_/Q _15750_/X _15697_/X _15751_/X vssd1 vssd1 vccd1 vccd1 _19649_/D
+ sky130_fd_sc_hd__a22o_1
X_12964_ _20704_/Q _12960_/X _12881_/X _12961_/X vssd1 vssd1 vccd1 vccd1 _20704_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_234_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14703_ _14705_/A vssd1 vssd1 vccd1 vccd1 _14723_/A sky130_fd_sc_hd__clkbuf_2
X_18471_ _18470_/X _16944_/Y _18680_/S vssd1 vssd1 vccd1 vccd1 _18471_/X sky130_fd_sc_hd__mux2_2
X_11915_ _11913_/A _15396_/B _11913_/Y vssd1 vssd1 vccd1 vccd1 _21012_/D sky130_fd_sc_hd__a21oi_1
XFILLER_206_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15683_ _19681_/Q _15681_/X _15585_/X _15682_/X vssd1 vssd1 vccd1 vccd1 _19681_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12895_ _13108_/B vssd1 vssd1 vccd1 vccd1 _17085_/A sky130_fd_sc_hd__buf_4
XPHY_4461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19969__RESET_B repeater184/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17422_ _19401_/Q vssd1 vssd1 vccd1 vccd1 _17422_/Y sky130_fd_sc_hd__inv_2
X_14634_ _20187_/Q _14636_/B _14624_/X _14577_/B vssd1 vssd1 vccd1 vccd1 _20187_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__20565__CLK _20592_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11846_ _11842_/B _11827_/A _11845_/X _11834_/X _11845_/A vssd1 vssd1 vccd1 vccd1
+ _11847_/A sky130_fd_sc_hd__o32a_1
XPHY_4494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17353_ _19343_/Q vssd1 vssd1 vccd1 vccd1 _17353_/Y sky130_fd_sc_hd__inv_2
X_11777_ _16507_/A vssd1 vssd1 vccd1 vccd1 _16516_/A sky130_fd_sc_hd__buf_1
XFILLER_202_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14565_ _14526_/Y _19121_/X _14534_/X _14564_/X vssd1 vssd1 vccd1 vccd1 _20208_/D
+ sky130_fd_sc_hd__o22ai_1
XANTENNA_repeater261_A repeater262/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19250__S1 _20131_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18705__S _18926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16304_ _19386_/Q _16298_/X _16285_/X _16300_/X vssd1 vssd1 vccd1 vccd1 _19386_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_202_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10728_ _10723_/A _10723_/B _10723_/C vssd1 vssd1 vccd1 vccd1 _10729_/B sky130_fd_sc_hd__o21a_1
X_13516_ _20436_/Q _13514_/X _13446_/X _13515_/X vssd1 vssd1 vccd1 vccd1 _20436_/D
+ sky130_fd_sc_hd__a22o_1
X_17284_ _20398_/Q vssd1 vssd1 vccd1 vccd1 _17284_/Y sky130_fd_sc_hd__inv_2
X_14496_ _14496_/A vssd1 vssd1 vccd1 vccd1 _14518_/B sky130_fd_sc_hd__buf_1
X_19023_ _16899_/X _20400_/Q _19026_/S vssd1 vssd1 vccd1 vccd1 _19953_/D sky130_fd_sc_hd__mux2_1
X_16235_ _16235_/A vssd1 vssd1 vccd1 vccd1 _16235_/X sky130_fd_sc_hd__buf_2
X_10659_ _10659_/A _10659_/B vssd1 vssd1 vccd1 vccd1 _10683_/A sky130_fd_sc_hd__or2_1
X_13447_ _13447_/A vssd1 vssd1 vccd1 vccd1 _13447_/X sky130_fd_sc_hd__buf_1
XFILLER_6_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09628__A input50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16166_ _16173_/A vssd1 vssd1 vccd1 vccd1 _16166_/X sky130_fd_sc_hd__buf_1
X_13378_ _13378_/A vssd1 vssd1 vccd1 vccd1 _13378_/X sky130_fd_sc_hd__buf_1
XFILLER_126_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15117_ _20446_/Q _20057_/Q _15116_/Y _15071_/A vssd1 vssd1 vccd1 vccd1 _15117_/X
+ sky130_fd_sc_hd__o22a_1
X_12329_ _12329_/A _12329_/B vssd1 vssd1 vccd1 vccd1 _12342_/A sky130_fd_sc_hd__or2_1
X_16097_ _19485_/Q _16094_/X _15865_/X _16096_/X vssd1 vssd1 vccd1 vccd1 _19485_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18440__S _18909_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_113_HCLK_A clkbuf_opt_3_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19925_ _21342_/CLK _19925_/D repeater211/X vssd1 vssd1 vccd1 vccd1 _19925_/Q sky130_fd_sc_hd__dfrtp_1
X_15048_ _20054_/Q vssd1 vssd1 vccd1 vccd1 _15068_/A sky130_fd_sc_hd__inv_2
XANTENNA__12989__A input61/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19856_ _21162_/CLK _19856_/D repeater227/X vssd1 vssd1 vccd1 vccd1 _19856_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_84_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18807_ _18806_/X _10262_/A _18841_/S vssd1 vssd1 vccd1 vccd1 _18807_/X sky130_fd_sc_hd__mux2_1
X_19787_ _19789_/CLK _19787_/D vssd1 vssd1 vccd1 vccd1 _19787_/Q sky130_fd_sc_hd__dfxtp_1
X_16999_ _16999_/A _16999_/B vssd1 vssd1 vccd1 vccd1 _16999_/Y sky130_fd_sc_hd__nor2_1
XFILLER_37_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18738_ _18737_/X _17607_/Y _18929_/S vssd1 vssd1 vccd1 vccd1 _18738_/X sky130_fd_sc_hd__mux2_1
XFILLER_243_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18669_ _18668_/X _14442_/Y _18669_/S vssd1 vssd1 vccd1 vccd1 _18669_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15404__B1 _15343_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20700_ _21294_/CLK _20700_/D repeater209/X vssd1 vssd1 vccd1 vccd1 _20700_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_24_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13613__A _13625_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_211_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20631_ _21481_/CLK _20631_/D repeater206/X vssd1 vssd1 vccd1 vccd1 _20631_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18615__S _18928_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19241__S1 _20133_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15168__C1 _15201_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20562_ _20724_/CLK _20562_/D repeater264/X vssd1 vssd1 vccd1 vccd1 _20562_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_220_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20493_ _20495_/CLK _20493_/D repeater273/X vssd1 vssd1 vccd1 vccd1 _20493_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_164_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20197__RESET_B repeater193/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20126__RESET_B repeater247/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18350__S _18886_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21114_ _21120_/CLK _21114_/D repeater233/X vssd1 vssd1 vccd1 vccd1 _21114_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12899__A _12899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21045_ _21193_/CLK _21045_/D repeater224/X vssd1 vssd1 vccd1 vccd1 _21045_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_115_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09807_ _09804_/A _09806_/A _21459_/Q _16620_/B vssd1 vssd1 vccd1 vccd1 _09807_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_75_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_98_HCLK_A clkbuf_4_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_12_0_HCLK_A clkbuf_3_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09738_ _21226_/Q vssd1 vssd1 vccd1 vccd1 _11052_/C sky130_fd_sc_hd__inv_2
XFILLER_216_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09669_ _15377_/A vssd1 vssd1 vccd1 vccd1 _12544_/A sky130_fd_sc_hd__clkbuf_4
XPHY_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11700_ _21079_/Q _11697_/X _11680_/X _11699_/X vssd1 vssd1 vccd1 vccd1 _21079_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12680_ _12680_/A vssd1 vssd1 vccd1 vccd1 _12680_/X sky130_fd_sc_hd__buf_1
XPHY_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11631_ _14813_/C _11631_/B vssd1 vssd1 vccd1 vccd1 _11632_/B sky130_fd_sc_hd__nand2_1
XFILLER_24_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20829_ _20841_/CLK _20829_/D repeater251/X vssd1 vssd1 vccd1 vccd1 _20829_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09625__A1 _21485_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20967__RESET_B repeater186/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18525__S _18908_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19232__S1 _21004_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14350_ _20210_/Q vssd1 vssd1 vccd1 vccd1 _14518_/C sky130_fd_sc_hd__inv_2
X_11562_ _11562_/A vssd1 vssd1 vccd1 vccd1 _11562_/X sky130_fd_sc_hd__buf_1
XPHY_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10513_ _20691_/Q vssd1 vssd1 vccd1 vccd1 _10513_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13709__B1 _13707_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13301_ _13301_/A vssd1 vssd1 vccd1 vccd1 _13322_/A sky130_fd_sc_hd__buf_1
XFILLER_210_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14281_ _20128_/Q vssd1 vssd1 vccd1 vccd1 _16451_/A sky130_fd_sc_hd__inv_2
XPHY_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11493_ _13327_/A _13327_/B _14303_/C vssd1 vssd1 vccd1 vccd1 _17169_/D sky130_fd_sc_hd__or3_4
XFILLER_183_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13232_ _20577_/Q _13226_/X _13148_/X _13228_/X vssd1 vssd1 vccd1 vccd1 _20577_/D
+ sky130_fd_sc_hd__a22o_1
X_16020_ _16297_/A _16107_/B _16344_/C vssd1 vssd1 vccd1 vccd1 _16028_/A sky130_fd_sc_hd__or3_4
XANTENNA_input72_A MSI_S3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10444_ _10782_/A _20695_/Q _21284_/Q _10443_/Y vssd1 vssd1 vccd1 vccd1 _10444_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_108_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11196__B1 _10896_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13163_ _13163_/A vssd1 vssd1 vccd1 vccd1 _13163_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__18260__S _18787_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10375_ _10397_/A vssd1 vssd1 vccd1 vccd1 _10375_/X sky130_fd_sc_hd__buf_2
XFILLER_123_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12114_ _20971_/Q vssd1 vssd1 vccd1 vccd1 _12324_/A sky130_fd_sc_hd__inv_2
XFILLER_69_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17971_ _18204_/X _17963_/X _18302_/X _17947_/A vssd1 vssd1 vccd1 vccd1 _17971_/X
+ sky130_fd_sc_hd__o22a_1
X_13094_ _20641_/Q _13092_/X _12950_/X _13093_/X vssd1 vssd1 vccd1 vccd1 _20641_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_2_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19710_ _19776_/CLK _19710_/D vssd1 vssd1 vccd1 vccd1 _19710_/Q sky130_fd_sc_hd__dfxtp_1
X_16922_ _16922_/A vssd1 vssd1 vccd1 vccd1 _16927_/B sky130_fd_sc_hd__inv_2
X_12045_ _20392_/Q vssd1 vssd1 vccd1 vccd1 _12045_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12696__B1 _09659_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18820__A0 _17079_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20241__D _20241_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19641_ _20326_/CLK _19641_/D vssd1 vssd1 vccd1 vccd1 _19641_/Q sky130_fd_sc_hd__dfxtp_1
X_16853_ _19942_/Q _16853_/B vssd1 vssd1 vccd1 vccd1 _16853_/X sky130_fd_sc_hd__and2_1
XFILLER_37_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19091__S _19870_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15634__B1 _15585_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15804_ _19628_/Q _15800_/X _09821_/X _15802_/X vssd1 vssd1 vccd1 vccd1 _19628_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_1_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19572_ _19776_/CLK _19572_/D vssd1 vssd1 vccd1 vccd1 _19572_/Q sky130_fd_sc_hd__dfxtp_1
X_16784_ _16820_/A _16784_/B vssd1 vssd1 vccd1 vccd1 _16784_/Y sky130_fd_sc_hd__nor2_1
XFILLER_225_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13996_ _13996_/A vssd1 vssd1 vccd1 vccd1 _13996_/Y sky130_fd_sc_hd__inv_2
XFILLER_218_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18523_ _18522_/X _12165_/Y _18787_/S vssd1 vssd1 vccd1 vccd1 _18523_/X sky130_fd_sc_hd__mux2_2
X_15735_ _19658_/Q _15723_/X _15694_/X _15727_/X vssd1 vssd1 vccd1 vccd1 _19658_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12947_ _20711_/Q _12942_/X _12699_/X _12943_/X vssd1 vssd1 vccd1 vccd1 _20711_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11671__A1 _16654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18454_ _18453_/X _10766_/A _18617_/S vssd1 vssd1 vccd1 vccd1 _18454_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15666_ _15666_/A vssd1 vssd1 vccd1 vccd1 _15666_/X sky130_fd_sc_hd__buf_1
XPHY_4280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12878_ _16338_/A vssd1 vssd1 vccd1 vccd1 _13710_/A sky130_fd_sc_hd__clkbuf_4
XPHY_4291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17405_ _17060_/B _17396_/X _17400_/X _17403_/X _17404_/X vssd1 vssd1 vccd1 vccd1
+ _17405_/X sky130_fd_sc_hd__o2111a_1
X_14617_ _20197_/Q _14616_/Y _14610_/X _14587_/B vssd1 vssd1 vccd1 vccd1 _20197_/D
+ sky130_fd_sc_hd__o211a_1
X_18385_ _18384_/X _12154_/Y _18909_/S vssd1 vssd1 vccd1 vccd1 _18385_/X sky130_fd_sc_hd__mux2_1
X_11829_ _21036_/Q _11829_/B vssd1 vssd1 vccd1 vccd1 _11829_/Y sky130_fd_sc_hd__nor2_1
X_15597_ _15603_/A vssd1 vssd1 vccd1 vccd1 _15604_/A sky130_fd_sc_hd__inv_2
XANTENNA__18435__S _18884_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19223__S1 _21004_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17336_ _19392_/Q vssd1 vssd1 vccd1 vccd1 _17336_/Y sky130_fd_sc_hd__inv_2
X_14548_ _14751_/B vssd1 vssd1 vccd1 vccd1 _14548_/X sky130_fd_sc_hd__buf_1
X_17267_ _19615_/Q vssd1 vssd1 vccd1 vccd1 _17267_/Y sky130_fd_sc_hd__inv_2
X_14479_ _14463_/D _14374_/B _14476_/Y _14474_/X vssd1 vssd1 vccd1 vccd1 _20231_/D
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__14264__A _14264_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19006_ _16974_/Y _20417_/Q _19019_/S vssd1 vssd1 vccd1 vccd1 _19970_/D sky130_fd_sc_hd__mux2_1
X_16218_ _16224_/A vssd1 vssd1 vccd1 vccd1 _16218_/X sky130_fd_sc_hd__buf_1
XFILLER_127_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_160_HCLK clkbuf_opt_0_HCLK/A vssd1 vssd1 vccd1 vccd1 _19828_/CLK sky130_fd_sc_hd__clkbuf_16
X_17198_ _17194_/Y _17196_/X _17197_/Y _17169_/D vssd1 vssd1 vccd1 vccd1 _17235_/A
+ sky130_fd_sc_hd__o22a_2
XANTENNA__18103__A2 _17862_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16149_ _19462_/Q _16141_/X _15916_/X _16143_/X vssd1 vssd1 vccd1 vccd1 _19462_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17847__D1 _17846_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18170__S _18644_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19908_ _21185_/CLK _19908_/D repeater221/X vssd1 vssd1 vccd1 vccd1 _19908_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__13608__A _13626_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_216_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18811__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19839_ _21151_/CLK _19839_/D repeater223/X vssd1 vssd1 vccd1 vccd1 _19839_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_110_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13100__A1 _20637_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17917__A2 _18020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_213_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11662__A1 _11504_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18345__S _18908_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16654__A _16654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19214__S1 _21004_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20614_ _20622_/CLK _20614_/D repeater196/X vssd1 vssd1 vccd1 vccd1 _20614_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_177_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20378__RESET_B repeater185/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20545_ _20724_/CLK _20545_/D repeater263/X vssd1 vssd1 vccd1 vccd1 _20545_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_153_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20476_ _20476_/CLK _20476_/D repeater280/X vssd1 vssd1 vccd1 vccd1 _20476_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_118_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20260__CLK _20592_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10160_ _10160_/A _10179_/A vssd1 vssd1 vccd1 vccd1 _10161_/B sky130_fd_sc_hd__or2_2
XFILLER_106_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12678__B1 _09628_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10091_ _21397_/Q _10090_/Y _10034_/B _20800_/Q vssd1 vssd1 vccd1 vccd1 _10091_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_126_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19150__S0 _19285_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21166__RESET_B repeater225/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21028_ _21255_/CLK _21028_/D repeater241/X vssd1 vssd1 vccd1 vccd1 _21028_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17605__A1 _11940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15733__A _16237_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13850_ _20311_/Q vssd1 vssd1 vccd1 vccd1 _13971_/B sky130_fd_sc_hd__inv_2
XFILLER_235_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12801_ _20778_/Q _12797_/X _12550_/X _12798_/X vssd1 vssd1 vccd1 vccd1 _20778_/D
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_41_HCLK clkbuf_4_11_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20908_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_62_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13781_ _20182_/Q vssd1 vssd1 vccd1 vccd1 _14572_/A sky130_fd_sc_hd__inv_2
X_10993_ _21019_/Q vssd1 vssd1 vccd1 vccd1 _10993_/Y sky130_fd_sc_hd__inv_2
X_15520_ _19761_/Q _15516_/X _15518_/X _15519_/X vssd1 vssd1 vccd1 vccd1 _19761_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_243_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12732_ _20806_/Q vssd1 vssd1 vccd1 vccd1 _12734_/A sky130_fd_sc_hd__inv_2
XFILLER_35_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16041__B1 _16006_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15451_ _15459_/A vssd1 vssd1 vccd1 vccd1 _15460_/A sky130_fd_sc_hd__inv_2
XFILLER_231_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12663_ input57/X vssd1 vssd1 vccd1 vccd1 _12663_/X sky130_fd_sc_hd__clkbuf_4
XPHY_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18255__S _18898_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19205__S1 _21004_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14402_ _21476_/Q vssd1 vssd1 vccd1 vccd1 _14402_/Y sky130_fd_sc_hd__inv_2
XPHY_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11614_ _21111_/Q _11614_/B vssd1 vssd1 vccd1 vccd1 _11614_/Y sky130_fd_sc_hd__nand2_1
XPHY_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18170_ _18169_/X _10086_/Y _18644_/S vssd1 vssd1 vccd1 vccd1 _18170_/X sky130_fd_sc_hd__mux2_1
XPHY_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15382_ _15382_/A vssd1 vssd1 vccd1 vccd1 _15661_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__20730__RESET_B repeater257/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12594_ _12600_/A vssd1 vssd1 vccd1 vccd1 _12594_/X sky130_fd_sc_hd__buf_1
XPHY_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17121_ _19574_/Q vssd1 vssd1 vccd1 vccd1 _17121_/Y sky130_fd_sc_hd__inv_2
XPHY_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14333_ _14333_/A vssd1 vssd1 vccd1 vccd1 _14463_/D sky130_fd_sc_hd__buf_1
X_11545_ _11545_/A _11545_/B vssd1 vssd1 vccd1 vccd1 _11545_/X sky130_fd_sc_hd__or2_1
XPHY_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17052_ _20042_/Q _20040_/Q _20041_/Q _17051_/X vssd1 vssd1 vccd1 vccd1 _19849_/D
+ sky130_fd_sc_hd__a22o_1
X_11476_ _19099_/X _11474_/X _21159_/Q _11475_/X vssd1 vssd1 vccd1 vccd1 _21159_/D
+ sky130_fd_sc_hd__a22o_1
X_14264_ _14264_/A vssd1 vssd1 vccd1 vccd1 _14264_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_167_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16003_ _19533_/Q _16000_/X _15969_/X _16002_/X vssd1 vssd1 vccd1 vccd1 _19533_/D
+ sky130_fd_sc_hd__a22o_1
X_10427_ _10422_/Y _20697_/Q _21286_/Q _10423_/Y _10426_/X vssd1 vssd1 vccd1 vccd1
+ _10446_/A sky130_fd_sc_hd__o221a_1
X_13215_ _13215_/A vssd1 vssd1 vccd1 vccd1 _13215_/X sky130_fd_sc_hd__buf_1
XANTENNA_repeater224_A repeater226/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14195_ _14195_/A vssd1 vssd1 vccd1 vccd1 _14195_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20753__CLK _21342_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13146_ input42/X vssd1 vssd1 vccd1 vccd1 _13146_/X sky130_fd_sc_hd__clkbuf_4
X_10358_ _21375_/Q _10356_/Y _21368_/Q _18035_/A vssd1 vssd1 vccd1 vccd1 _10358_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_2_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15855__B1 _15785_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18003__B _18006_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13428__A _13444_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17954_ _17954_/A vssd1 vssd1 vccd1 vccd1 _17954_/X sky130_fd_sc_hd__buf_1
X_13077_ _20650_/Q _13072_/X _12932_/X _13073_/X vssd1 vssd1 vccd1 vccd1 _20650_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_239_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12669__B1 _12668_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10289_ _10289_/A _10289_/B vssd1 vssd1 vccd1 vccd1 _10290_/A sky130_fd_sc_hd__or2_1
X_12028_ _19078_/X _12023_/X _20987_/Q _12024_/X vssd1 vssd1 vccd1 vccd1 _20987_/D
+ sky130_fd_sc_hd__a22o_1
X_16905_ _16905_/A vssd1 vssd1 vccd1 vccd1 _16910_/B sky130_fd_sc_hd__inv_2
XFILLER_66_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17885_ _20410_/Q vssd1 vssd1 vccd1 vccd1 _17885_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19984__RESET_B repeater185/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19624_ _20890_/CLK _19624_/D vssd1 vssd1 vccd1 vccd1 _19624_/Q sky130_fd_sc_hd__dfxtp_1
X_16836_ _19938_/Q _16843_/B vssd1 vssd1 vccd1 vccd1 _16836_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_81_HCLK_A clkbuf_4_13_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19913__RESET_B repeater220/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09641__A _12849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19555_ _19706_/CLK _19555_/D vssd1 vssd1 vccd1 vccd1 _19555_/Q sky130_fd_sc_hd__dfxtp_1
X_16767_ _16770_/B _16766_/Y _16762_/X vssd1 vssd1 vccd1 vccd1 _16767_/X sky130_fd_sc_hd__o21a_1
XANTENNA__13094__B1 _12950_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20889__RESET_B repeater185/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13979_ _13979_/A vssd1 vssd1 vccd1 vccd1 _13979_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13163__A _13163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18506_ _18505_/X _10095_/Y _18644_/S vssd1 vssd1 vccd1 vccd1 _18506_/X sky130_fd_sc_hd__mux2_1
X_15718_ _19665_/Q _15716_/X _15697_/X _15717_/X vssd1 vssd1 vccd1 vccd1 _19665_/D
+ sky130_fd_sc_hd__a22o_1
X_19486_ _19961_/CLK _19486_/D vssd1 vssd1 vccd1 vccd1 _19486_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_202_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16698_ _16700_/A _18943_/X vssd1 vssd1 vccd1 vccd1 _19893_/D sky130_fd_sc_hd__and2_1
XANTENNA__20818__RESET_B repeater211/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18437_ _18436_/X _10272_/A _18841_/S vssd1 vssd1 vccd1 vccd1 _18437_/X sky130_fd_sc_hd__mux2_1
X_15649_ _19697_/Q _15647_/X _15480_/X _15648_/X vssd1 vssd1 vccd1 vccd1 _19697_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16474__A _16474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18165__S _18904_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_221_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18368_ _18367_/X _21297_/Q _18617_/S vssd1 vssd1 vccd1 vccd1 _18368_/X sky130_fd_sc_hd__mux2_1
XFILLER_221_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17319_ _17732_/A vssd1 vssd1 vccd1 vccd1 _17319_/X sky130_fd_sc_hd__buf_1
XFILLER_186_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20400__RESET_B repeater270/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18299_ _17281_/X _17968_/Y _18835_/S vssd1 vssd1 vccd1 vccd1 _18299_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13149__A1 _20611_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20330_ _20331_/CLK _20330_/D repeater190/X vssd1 vssd1 vccd1 vccd1 _20330_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_116_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20261_ _21366_/CLK _20261_/D repeater264/X vssd1 vssd1 vccd1 vccd1 _20261_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__10907__B1 _21248_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20192_ _20626_/CLK _20192_/D repeater200/X vssd1 vssd1 vccd1 vccd1 _20192_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_88_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19132__S0 _19285_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_64_HCLK clkbuf_4_11_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _21338_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_56_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10135__B2 _10132_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_229_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12896__B _12899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13085__B1 _12857_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13073__A _13073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_225_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12832__B1 _12666_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19199__S0 _20130_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20141__RESET_B repeater250/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18803__S _18879_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11330_ _11375_/A vssd1 vssd1 vccd1 vccd1 _11357_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_166_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20528_ _20944_/CLK _20528_/D repeater274/X vssd1 vssd1 vccd1 vccd1 _20528_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_181_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11261_ _20911_/Q vssd1 vssd1 vccd1 vccd1 _11286_/C sky130_fd_sc_hd__buf_1
XFILLER_181_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20459_ _20937_/CLK _20459_/D repeater276/X vssd1 vssd1 vccd1 vccd1 _20459_/Q sky130_fd_sc_hd__dfrtp_1
X_13000_ _20692_/Q _12995_/X _12999_/X _12997_/X vssd1 vssd1 vccd1 vccd1 _20692_/D
+ sky130_fd_sc_hd__a22o_1
X_10212_ _10205_/A _10205_/B _10210_/Y _10177_/X vssd1 vssd1 vccd1 vccd1 _21384_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_97_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21347__RESET_B repeater210/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11192_ _11192_/A vssd1 vssd1 vccd1 vccd1 _11193_/A sky130_fd_sc_hd__inv_2
XFILLER_106_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10143_ _10177_/A vssd1 vssd1 vccd1 vccd1 _10227_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA_input35_A HSEL vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14951_ _15059_/B vssd1 vssd1 vccd1 vccd1 _14978_/A sky130_fd_sc_hd__buf_1
XFILLER_88_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10074_ _10160_/A _10159_/A _10162_/A _10161_/A vssd1 vssd1 vccd1 vccd1 _10075_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_102_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13902_ _20640_/Q _14013_/A _20661_/Q _13894_/B _13901_/X vssd1 vssd1 vccd1 vccd1
+ _13914_/A sky130_fd_sc_hd__o221a_1
X_17670_ _19364_/Q vssd1 vssd1 vccd1 vccd1 _17670_/Y sky130_fd_sc_hd__inv_2
X_14882_ _14882_/A _14957_/A vssd1 vssd1 vccd1 vccd1 _14883_/B sky130_fd_sc_hd__or2_1
XFILLER_247_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16621_ _16621_/A vssd1 vssd1 vccd1 vccd1 _16621_/Y sky130_fd_sc_hd__inv_2
X_13833_ _20200_/Q vssd1 vssd1 vccd1 vccd1 _14589_/A sky130_fd_sc_hd__inv_2
XANTENNA__20982__RESET_B repeater187/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13076__B1 _12930_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19340_ _20142_/CLK _19340_/D vssd1 vssd1 vccd1 vccd1 _19340_/Q sky130_fd_sc_hd__dfxtp_1
X_16552_ _16547_/Y _16550_/Y _16551_/Y _19913_/Q vssd1 vssd1 vccd1 vccd1 _16584_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_189_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20911__RESET_B repeater218/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13764_ _20612_/Q vssd1 vssd1 vccd1 vccd1 _13764_/Y sky130_fd_sc_hd__inv_2
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10976_ _20870_/Q _20869_/Q _11200_/A vssd1 vssd1 vccd1 vccd1 _12715_/A sky130_fd_sc_hd__or3_4
XFILLER_43_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15503_ _19767_/Q _15499_/X _15429_/X _15500_/X vssd1 vssd1 vccd1 vccd1 _19767_/D
+ sky130_fd_sc_hd__a22o_1
X_19271_ _19267_/X _19268_/X _19269_/X _19270_/X _20132_/Q _20133_/Q vssd1 vssd1 vccd1
+ vccd1 _19271_/X sky130_fd_sc_hd__mux4_2
X_12715_ _12715_/A vssd1 vssd1 vccd1 vccd1 _17639_/A sky130_fd_sc_hd__buf_4
XANTENNA__20229__RESET_B repeater200/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16483_ _20129_/Q vssd1 vssd1 vccd1 vccd1 _16483_/Y sky130_fd_sc_hd__inv_2
X_13695_ _20343_/Q _13693_/X _12860_/A _13694_/X vssd1 vssd1 vccd1 vccd1 _20343_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_repeater174_A _18885_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18222_ _20846_/Q input26/X _18236_/S vssd1 vssd1 vccd1 vccd1 _18222_/X sky130_fd_sc_hd__mux2_4
XANTENNA__13379__A1 _20501_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15434_ _15441_/A vssd1 vssd1 vccd1 vccd1 _15434_/X sky130_fd_sc_hd__buf_1
XFILLER_175_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12646_ _12753_/A _12713_/B _13047_/C vssd1 vssd1 vccd1 vccd1 _17323_/A sky130_fd_sc_hd__or3_1
XPHY_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18153_ _18152_/X _20587_/Q _18907_/S vssd1 vssd1 vccd1 vccd1 _18153_/X sky130_fd_sc_hd__mux2_1
XFILLER_168_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15365_ _19826_/Q _15359_/X _15343_/X _15361_/X vssd1 vssd1 vccd1 vccd1 _19826_/D
+ sky130_fd_sc_hd__a22o_1
X_12577_ _20887_/Q _12574_/X _18239_/X _12575_/X vssd1 vssd1 vccd1 vccd1 _20887_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18713__S _18884_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17104_ _19718_/Q vssd1 vssd1 vccd1 vccd1 _17104_/Y sky130_fd_sc_hd__inv_2
X_14316_ _20127_/Q vssd1 vssd1 vccd1 vccd1 _16451_/B sky130_fd_sc_hd__inv_2
XPHY_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11528_ _11534_/A vssd1 vssd1 vccd1 vccd1 _11535_/A sky130_fd_sc_hd__inv_2
X_18084_ _20840_/Q _18084_/B vssd1 vssd1 vccd1 vccd1 _18084_/Y sky130_fd_sc_hd__nand2_1
X_15296_ _19862_/Q _15296_/B vssd1 vssd1 vccd1 vccd1 _15297_/B sky130_fd_sc_hd__or2_1
XFILLER_183_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17035_ _17035_/A _17035_/B vssd1 vssd1 vccd1 vccd1 _20019_/D sky130_fd_sc_hd__nor2_1
X_14247_ _20258_/Q _14246_/X _20257_/Q _18946_/S vssd1 vssd1 vccd1 vccd1 _20258_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13000__B1 _12999_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11459_ _11459_/A _19870_/D vssd1 vssd1 vccd1 vccd1 _11462_/A sky130_fd_sc_hd__or2_2
XFILLER_113_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09636__A input46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14178_ _14099_/A _14099_/B _14100_/Y _14215_/B vssd1 vssd1 vccd1 vccd1 _20289_/D
+ sky130_fd_sc_hd__a211oi_2
Xclkbuf_leaf_87_HCLK clkbuf_4_12_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _21407_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_97_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21017__RESET_B repeater238/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13129_ _20621_/Q _13126_/X _12918_/X _13127_/X vssd1 vssd1 vccd1 vccd1 _20621_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_98_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18986_ _21267_/Q _21119_/Q _18992_/S vssd1 vssd1 vccd1 vccd1 _18986_/X sky130_fd_sc_hd__mux2_1
XFILLER_239_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17937_ _17937_/A _17938_/B vssd1 vssd1 vccd1 vccd1 _17937_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__12997__A _13013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10117__B2 _20795_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15373__A _15505_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_239_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater147 _19058_/S vssd1 vssd1 vccd1 vccd1 _19046_/S sky130_fd_sc_hd__buf_8
X_17868_ _18573_/X _17853_/X _18557_/X _17854_/X vssd1 vssd1 vccd1 vccd1 _17868_/X
+ sky130_fd_sc_hd__o22a_1
Xrepeater158 _18850_/S vssd1 vssd1 vccd1 vccd1 _18904_/S sky130_fd_sc_hd__buf_8
XFILLER_227_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater169 _18849_/S vssd1 vssd1 vccd1 vccd1 _18903_/S sky130_fd_sc_hd__buf_8
XFILLER_94_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19607_ _20890_/CLK _19607_/D vssd1 vssd1 vccd1 vccd1 _19607_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16819_ _16822_/A _16822_/C _16818_/Y _16814_/Y vssd1 vssd1 vccd1 vccd1 _16820_/B
+ sky130_fd_sc_hd__o22a_1
X_17799_ _18676_/X _17216_/A _18380_/X _17223_/A vssd1 vssd1 vccd1 vccd1 _17799_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_242_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12814__A0 _12809_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19538_ _19789_/CLK _19538_/D vssd1 vssd1 vccd1 vccd1 _19538_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__19941__CLK _20930_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19469_ _19834_/CLK _19469_/D vssd1 vssd1 vccd1 vccd1 _19469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21431_ _21431_/CLK _21431_/D repeater236/X vssd1 vssd1 vccd1 vccd1 _21431_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18623__S _18666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_238_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21362_ _21368_/CLK _21362_/D repeater254/X vssd1 vssd1 vccd1 vccd1 _21362_/Q sky130_fd_sc_hd__dfrtp_1
X_20313_ _20316_/CLK _20313_/D repeater197/X vssd1 vssd1 vccd1 vccd1 _20313_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__15548__A _15661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21293_ _21294_/CLK _21293_/D repeater211/X vssd1 vssd1 vccd1 vccd1 _21293_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__10980__A _15505_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20244_ _21421_/CLK _20244_/D repeater214/X vssd1 vssd1 vccd1 vccd1 _20244_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_162_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20175_ _20241_/CLK _20175_/D repeater249/X vssd1 vssd1 vccd1 vccd1 _20175_/Q sky130_fd_sc_hd__dfrtp_4
X_09986_ _20021_/Q _09986_/B vssd1 vssd1 vccd1 vccd1 _09987_/A sky130_fd_sc_hd__nand2_1
XFILLER_77_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16244__B1 _16014_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13058__B1 _12991_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10830_ _10830_/A vssd1 vssd1 vccd1 vccd1 _10830_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__12805__B1 _11736_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10761_ _10761_/A _10829_/A vssd1 vssd1 vccd1 vccd1 _10762_/B sky130_fd_sc_hd__or2_2
XANTENNA__20322__RESET_B repeater262/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12500_ _12500_/A _12500_/B vssd1 vssd1 vccd1 vccd1 _16569_/C sky130_fd_sc_hd__or2_1
XFILLER_197_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10692_ _10655_/A _10655_/B _10685_/X _10690_/Y vssd1 vssd1 vccd1 vccd1 _21326_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_157_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13480_ _20453_/Q _13472_/X _13479_/X _13473_/X vssd1 vssd1 vccd1 vccd1 _20453_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_232_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12431_ _12431_/A _12431_/B vssd1 vssd1 vccd1 vccd1 _12443_/A sky130_fd_sc_hd__or2_2
XANTENNA__13230__B1 _13144_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18533__S _18903_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15150_ _15148_/Y _20065_/Q _15091_/Y _15092_/X _15149_/X vssd1 vssd1 vccd1 vccd1
+ _15157_/B sky130_fd_sc_hd__o221a_1
X_12362_ _12362_/A vssd1 vssd1 vccd1 vccd1 _12362_/Y sky130_fd_sc_hd__inv_2
XFILLER_193_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10595__B2 _10592_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14101_ _20290_/Q vssd1 vssd1 vccd1 vccd1 _14101_/Y sky130_fd_sc_hd__inv_2
X_11313_ _11287_/C _11313_/B _11313_/C vssd1 vssd1 vccd1 vccd1 _12504_/B sky130_fd_sc_hd__and3b_1
XFILLER_154_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15081_ _15081_/A _15176_/A vssd1 vssd1 vccd1 vccd1 _15082_/B sky130_fd_sc_hd__or2_2
XFILLER_5_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12293_ _20946_/Q _12291_/Y _12471_/A _20503_/Q vssd1 vssd1 vccd1 vccd1 _12293_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__21181__RESET_B repeater216/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11244_ _11250_/A vssd1 vssd1 vccd1 vccd1 _11244_/X sky130_fd_sc_hd__buf_1
XFILLER_4_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14032_ _13865_/B _14034_/A _13865_/A vssd1 vssd1 vccd1 vccd1 _14033_/B sky130_fd_sc_hd__o21a_1
XFILLER_107_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11175_ _11141_/X _11170_/Y _11173_/X vssd1 vssd1 vccd1 vccd1 _21221_/D sky130_fd_sc_hd__o21a_1
X_18840_ _18839_/X _17282_/Y _18885_/S vssd1 vssd1 vccd1 vccd1 _18840_/X sky130_fd_sc_hd__mux2_1
XANTENNA__15286__B2 _15160_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10126_ _20785_/Q vssd1 vssd1 vccd1 vccd1 _10126_/Y sky130_fd_sc_hd__inv_2
X_18771_ _18845_/A0 _10329_/Y _18884_/S vssd1 vssd1 vccd1 vccd1 _18771_/X sky130_fd_sc_hd__mux2_1
XANTENNA_output141_A _21185_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15983_ _19542_/Q _15978_/X _15951_/X _15979_/X vssd1 vssd1 vccd1 vccd1 _19542_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_94_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17722_ _19883_/Q vssd1 vssd1 vccd1 vccd1 _17722_/Y sky130_fd_sc_hd__inv_2
X_14934_ _20576_/Q vssd1 vssd1 vccd1 vccd1 _14934_/Y sky130_fd_sc_hd__inv_2
X_10057_ _21397_/Q vssd1 vssd1 vccd1 vccd1 _10158_/A sky130_fd_sc_hd__inv_2
XFILLER_209_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17653_ _16547_/Y _17550_/A _17652_/Y _17154_/X vssd1 vssd1 vccd1 vccd1 _17653_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_48_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14865_ _14997_/A _14963_/A vssd1 vssd1 vccd1 vccd1 _14866_/B sky130_fd_sc_hd__or2_2
XFILLER_224_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18708__S _18926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16604_ _16602_/Y _16603_/X _16585_/C _16541_/A vssd1 vssd1 vccd1 vccd1 _16604_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_217_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13816_ _20611_/Q _14577_/A _20619_/Q _14585_/A vssd1 vssd1 vccd1 vccd1 _13816_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__15921__A _15927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17584_ _18752_/X _17821_/A _18761_/X _17226_/A vssd1 vssd1 vccd1 vccd1 _17584_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_14796_ _14796_/A vssd1 vssd1 vccd1 vccd1 _14797_/A sky130_fd_sc_hd__inv_2
XFILLER_16_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19323_ _19626_/CLK _19323_/D vssd1 vssd1 vccd1 vccd1 _19323_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16535_ _16583_/A vssd1 vssd1 vccd1 vccd1 _16535_/X sky130_fd_sc_hd__buf_1
X_13747_ _20618_/Q _14584_/A _17898_/A _20190_/Q vssd1 vssd1 vccd1 vccd1 _13747_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_32_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20063__RESET_B repeater281/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17735__B1 _18691_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10959_ _21032_/Q vssd1 vssd1 vccd1 vccd1 _11845_/A sky130_fd_sc_hd__inv_2
XFILLER_189_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13441__A input64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19254_ _17338_/Y _17339_/Y _17340_/Y _17341_/Y _19275_/S0 _21004_/Q vssd1 vssd1
+ vccd1 vccd1 _19254_/X sky130_fd_sc_hd__mux4_2
XFILLER_231_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16466_ _16473_/A vssd1 vssd1 vccd1 vccd1 _16466_/X sky130_fd_sc_hd__buf_1
XFILLER_177_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13678_ _20352_/Q _13673_/X _13479_/X _13674_/X vssd1 vssd1 vccd1 vccd1 _20352_/D
+ sky130_fd_sc_hd__a22o_1
X_18205_ _17079_/Y _15262_/Y _18908_/S vssd1 vssd1 vccd1 vccd1 _18205_/X sky130_fd_sc_hd__mux2_1
X_15417_ _15425_/A vssd1 vssd1 vccd1 vccd1 _15417_/X sky130_fd_sc_hd__buf_1
XPHY_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12629_ input2/X _12625_/X _20853_/Q _12626_/X vssd1 vssd1 vccd1 vccd1 _20853_/D
+ sky130_fd_sc_hd__o22a_1
X_19185_ _19304_/Q _19826_/Q _19834_/Q _19418_/Q _19280_/S0 _20122_/Q vssd1 vssd1
+ vccd1 vccd1 _19185_/X sky130_fd_sc_hd__mux4_2
XANTENNA__18443__S _18787_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16397_ _19338_/Q _16392_/X _16237_/X _16394_/X vssd1 vssd1 vccd1 vccd1 _19338_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18136_ _17079_/Y _12057_/Y _18908_/S vssd1 vssd1 vccd1 vccd1 _18136_/X sky130_fd_sc_hd__mux2_1
X_15348_ _19833_/Q _15345_/X _15346_/X _15347_/X vssd1 vssd1 vccd1 vccd1 _19833_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_129_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18067_ _18386_/X _18024_/X _18512_/X _18064_/X _18066_/X vssd1 vssd1 vccd1 vccd1
+ _18068_/C sky130_fd_sc_hd__o221a_1
X_15279_ _15277_/Y _20074_/Q _15278_/Y _20057_/Q vssd1 vssd1 vccd1 vccd1 _15279_/X
+ sky130_fd_sc_hd__o22a_1
X_17018_ _20160_/Q _12743_/B _12743_/A _16526_/B vssd1 vssd1 vccd1 vccd1 _20003_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_208_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14721__B1 _14264_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09840_ _20034_/Q vssd1 vssd1 vccd1 vccd1 _09840_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_112_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09771_ _09783_/A _09812_/A _18963_/X _09771_/D vssd1 vssd1 vccd1 vccd1 _09777_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_58_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18969_ _11316_/B _12506_/B _20917_/Q vssd1 vssd1 vccd1 vccd1 _18969_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20931_ _20947_/CLK _20931_/D repeater266/X vssd1 vssd1 vccd1 vccd1 _20931_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18618__S _18903_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_240_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20862_ _21444_/CLK _20862_/D repeater246/X vssd1 vssd1 vccd1 vccd1 _20862_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_81_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14252__A2 _14246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_242_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20793_ _21407_/CLK _20793_/D repeater252/X vssd1 vssd1 vccd1 vccd1 _20793_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18353__S _18849_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21414_ _21419_/CLK _21414_/D repeater232/X vssd1 vssd1 vccd1 vccd1 _21414_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_194_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21345_ _21368_/CLK _21345_/D repeater255/X vssd1 vssd1 vccd1 vccd1 _21345_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_118_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21276_ _21445_/CLK _21276_/D repeater245/X vssd1 vssd1 vccd1 vccd1 _21276_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_2_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_8_0_HCLK clkbuf_4_9_0_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_opt_4_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_118_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20227_ _21485_/CLK _20227_/D repeater200/X vssd1 vssd1 vccd1 vccd1 _20227_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_104_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20158_ _20159_/CLK _20158_/D repeater189/X vssd1 vssd1 vccd1 vccd1 _20158_/Q sky130_fd_sc_hd__dfrtp_1
X_09969_ _09969_/A vssd1 vssd1 vccd1 vccd1 _09976_/A sky130_fd_sc_hd__inv_2
XFILLER_76_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13279__B1 _13277_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_218_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18206__A1 _15097_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12980_ _12978_/X _20698_/Q _12980_/S vssd1 vssd1 vccd1 vccd1 _20698_/D sky130_fd_sc_hd__mux2_1
XFILLER_57_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20089_ _20496_/CLK _20089_/D repeater273/X vssd1 vssd1 vccd1 vccd1 _20089_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_182_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11931_ _21007_/Q vssd1 vssd1 vccd1 vccd1 _11947_/A sky130_fd_sc_hd__buf_1
XFILLER_73_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20503__RESET_B repeater267/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17940__B _17943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18528__S _18669_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17965__B1 _18201_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14650_ _14568_/A _14568_/B _14639_/X _14648_/Y vssd1 vssd1 vccd1 vccd1 _20178_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_72_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11862_ _11862_/A vssd1 vssd1 vccd1 vccd1 _21028_/D sky130_fd_sc_hd__inv_2
XFILLER_33_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13601_ _13657_/B _13601_/B vssd1 vssd1 vccd1 vccd1 _13602_/S sky130_fd_sc_hd__or2_1
X_10813_ _21294_/Q _10811_/Y _10812_/X _10771_/B vssd1 vssd1 vccd1 vccd1 _21294_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_3942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14581_ _14581_/A _14581_/B vssd1 vssd1 vccd1 vccd1 _14623_/A sky130_fd_sc_hd__or2_1
XFILLER_14_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11793_ _12619_/A vssd1 vssd1 vccd1 vccd1 _11793_/X sky130_fd_sc_hd__buf_1
XPHY_3964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16320_ _16320_/A vssd1 vssd1 vccd1 vccd1 _16320_/X sky130_fd_sc_hd__buf_1
XANTENNA__13261__A _13261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13532_ _20430_/Q _13530_/Y _13530_/B _13531_/X vssd1 vssd1 vccd1 vccd1 _20430_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_43_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10744_ _19934_/Q _19937_/Q _19941_/Q vssd1 vssd1 vccd1 vccd1 _10746_/C sky130_fd_sc_hd__or3_2
XPHY_3997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18390__A0 _17079_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16251_ _19413_/Q _16248_/X _16109_/X _16250_/X vssd1 vssd1 vccd1 vccd1 _19413_/D
+ sky130_fd_sc_hd__a22o_1
X_13463_ _20463_/Q _13458_/X _13270_/X _13461_/X vssd1 vssd1 vccd1 vccd1 _20463_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13203__B1 _12999_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10675_ _10675_/A vssd1 vssd1 vccd1 vccd1 _10675_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18263__S _18903_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15202_ _15202_/A vssd1 vssd1 vccd1 vccd1 _15202_/Y sky130_fd_sc_hd__inv_2
X_12414_ _20396_/Q _12453_/A vssd1 vssd1 vccd1 vccd1 _12415_/A sky130_fd_sc_hd__or2_1
XANTENNA__21362__RESET_B repeater254/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18142__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16182_ _16188_/A vssd1 vssd1 vccd1 vccd1 _16182_/X sky130_fd_sc_hd__clkbuf_2
X_13394_ _20496_/Q _13390_/X _13265_/X _13393_/X vssd1 vssd1 vccd1 vccd1 _20496_/D
+ sky130_fd_sc_hd__a22o_1
X_15133_ _20445_/Q vssd1 vssd1 vccd1 vccd1 _15133_/Y sky130_fd_sc_hd__inv_2
X_12345_ _20977_/Q _12342_/Y _12344_/X _12331_/B vssd1 vssd1 vccd1 vccd1 _20977_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__18693__A1 _13939_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12605__A _12605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15064_ _15064_/A _15208_/A vssd1 vssd1 vccd1 vccd1 _15065_/B sky130_fd_sc_hd__or2_1
X_19941_ _20930_/CLK _19941_/D repeater268/X vssd1 vssd1 vccd1 vccd1 _19941_/Q sky130_fd_sc_hd__dfrtp_1
X_12276_ _12258_/A _20518_/Q _12407_/C _20527_/Q vssd1 vssd1 vccd1 vccd1 _12276_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_175_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11517__B1 _11516_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19094__S _19870_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14015_ _14015_/A _14015_/B vssd1 vssd1 vccd1 vccd1 _14020_/A sky130_fd_sc_hd__or2_1
X_11227_ _21200_/Q _11225_/X _10894_/X _11226_/X vssd1 vssd1 vccd1 vccd1 _21200_/D
+ sky130_fd_sc_hd__a22o_1
X_19872_ _21151_/CLK _19872_/D repeater223/X vssd1 vssd1 vccd1 vccd1 _19872_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__16456__B1 _11502_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18823_ _17372_/X _21414_/Q _20870_/Q vssd1 vssd1 vccd1 vccd1 _18823_/X sky130_fd_sc_hd__mux2_1
X_11158_ _20431_/Q vssd1 vssd1 vccd1 vccd1 _13181_/C sky130_fd_sc_hd__inv_2
XFILLER_1_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13436__A _13444_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10109_ _20780_/Q vssd1 vssd1 vccd1 vccd1 _10109_/Y sky130_fd_sc_hd__inv_2
X_11089_ _11089_/A vssd1 vssd1 vccd1 vccd1 _11090_/B sky130_fd_sc_hd__inv_2
X_15966_ _19550_/Q _15961_/X _15951_/X _15962_/X vssd1 vssd1 vccd1 vccd1 _19550_/D
+ sky130_fd_sc_hd__a22o_1
X_18754_ _18753_/X _20502_/Q _18910_/S vssd1 vssd1 vccd1 vccd1 _18754_/X sky130_fd_sc_hd__mux2_2
XFILLER_48_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_117_HCLK clkbuf_opt_3_HCLK/A vssd1 vssd1 vccd1 vccd1 _20943_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__17405__C1 _17403_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14917_ _14914_/Y _20076_/Q _14915_/Y _20091_/Q _14916_/X vssd1 vssd1 vccd1 vccd1
+ _14918_/D sky130_fd_sc_hd__o221a_1
X_17705_ _21437_/Q _17776_/B vssd1 vssd1 vccd1 vccd1 _17705_/Y sky130_fd_sc_hd__nand2_1
XFILLER_48_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13690__B1 _12853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18438__S _18666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15897_ _15897_/A vssd1 vssd1 vccd1 vccd1 _15897_/X sky130_fd_sc_hd__buf_1
X_18685_ _18684_/X _10266_/A _18841_/S vssd1 vssd1 vccd1 vccd1 _18685_/X sky130_fd_sc_hd__mux2_1
XANTENNA__16747__A _16835_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_224_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17636_ _20402_/Q vssd1 vssd1 vccd1 vccd1 _17636_/Y sky130_fd_sc_hd__inv_2
X_14848_ _20497_/Q vssd1 vssd1 vccd1 vccd1 _14997_/A sky130_fd_sc_hd__inv_2
XFILLER_36_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17567_ _17562_/Y _17553_/X _17563_/Y _17387_/X _17566_/X vssd1 vssd1 vccd1 vccd1
+ _17567_/X sky130_fd_sc_hd__o221a_1
XFILLER_63_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14779_ _14779_/A _14779_/B vssd1 vssd1 vccd1 vccd1 _14779_/Y sky130_fd_sc_hd__nor2_1
XFILLER_51_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13171__A _13171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_136_HCLK_A clkbuf_4_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16518_ _21092_/Q vssd1 vssd1 vccd1 vccd1 _16518_/Y sky130_fd_sc_hd__inv_2
X_19306_ _20172_/CLK _19306_/D vssd1 vssd1 vccd1 vccd1 _19306_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18381__A0 _17079_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17498_ _19296_/Q vssd1 vssd1 vccd1 vccd1 _17498_/Y sky130_fd_sc_hd__inv_2
XFILLER_189_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16449_ _17055_/B _19850_/Q vssd1 vssd1 vccd1 vccd1 _16449_/X sky130_fd_sc_hd__or2_1
X_19237_ _17428_/Y _17429_/Y _17430_/Y _17431_/Y _20130_/Q _20131_/Q vssd1 vssd1 vccd1
+ vccd1 _19237_/X sky130_fd_sc_hd__mux4_1
XANTENNA__18173__S _18886_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19168_ _19543_/Q _19535_/Q _19527_/Q _19511_/Q _19280_/S0 _20122_/Q vssd1 vssd1
+ vccd1 vccd1 _19168_/X sky130_fd_sc_hd__mux4_2
XFILLER_118_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18119_ vssd1 vssd1 vccd1 vccd1 _18119_/HI _18119_/LO sky130_fd_sc_hd__conb_1
XFILLER_145_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21032__RESET_B repeater242/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20837__CLK _20930_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18684__A1 _10081_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19099_ _16671_/X _21079_/Q _19870_/D vssd1 vssd1 vccd1 vccd1 _19099_/X sky130_fd_sc_hd__mux2_1
XANTENNA__18901__S _18901_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21130_ _21134_/CLK _21130_/D repeater192/X vssd1 vssd1 vccd1 vccd1 _21130_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17892__C1 _17891_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21061_ _21191_/CLK _21061_/D repeater227/X vssd1 vssd1 vccd1 vccd1 _21061_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18436__A1 _10132_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20012_ _21438_/CLK _20012_/D repeater237/X vssd1 vssd1 vccd1 vccd1 _20012_/Q sky130_fd_sc_hd__dfrtp_1
X_09823_ _21450_/Q vssd1 vssd1 vccd1 vccd1 _15873_/A sky130_fd_sc_hd__buf_1
XFILLER_86_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09754_ _21227_/Q _09752_/Y _11093_/A _20152_/Q vssd1 vssd1 vccd1 vccd1 _09754_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_228_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09685_ _10892_/A vssd1 vssd1 vccd1 vccd1 _09685_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_55_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18348__S _18884_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20914_ _21196_/CLK _20914_/D repeater218/X vssd1 vssd1 vccd1 vccd1 _20914_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13433__B1 _13432_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20845_ _20857_/CLK _20845_/D repeater243/X vssd1 vssd1 vccd1 vccd1 _20845_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20776_ _21379_/CLK _20776_/D repeater213/X vssd1 vssd1 vccd1 vccd1 _20776_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_11_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_58_HCLK_A clkbuf_4_14_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10460_ _21296_/Q vssd1 vssd1 vccd1 vccd1 _10772_/A sky130_fd_sc_hd__inv_2
XFILLER_108_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12716__D_N _20875_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10391_ _10391_/A vssd1 vssd1 vccd1 vccd1 _10391_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18811__S _18896_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12130_ _20955_/Q _12125_/Y _20970_/Q _17975_/A _12129_/X vssd1 vssd1 vccd1 vccd1
+ _12144_/B sky130_fd_sc_hd__o221a_1
X_21328_ _21341_/CLK _21328_/D repeater201/X vssd1 vssd1 vccd1 vccd1 _21328_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17883__C1 _17882_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12061_ _20367_/Q vssd1 vssd1 vccd1 vccd1 _12061_/Y sky130_fd_sc_hd__inv_2
X_21259_ _21390_/CLK _21259_/D repeater239/X vssd1 vssd1 vccd1 vccd1 _21259_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__20755__RESET_B repeater205/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16438__B1 _11502_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11012_ _11012_/A _11012_/B _11012_/C _11983_/C vssd1 vssd1 vccd1 vccd1 _11012_/X
+ sky130_fd_sc_hd__or4b_4
XFILLER_49_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15820_ _19621_/Q _15817_/X _09818_/X _15819_/X vssd1 vssd1 vccd1 vccd1 _19621_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_93_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15751_ _15751_/A vssd1 vssd1 vccd1 vccd1 _15751_/X sky130_fd_sc_hd__buf_1
X_12963_ _20705_/Q _12960_/X _12879_/X _12961_/X vssd1 vssd1 vccd1 vccd1 _20705_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18258__S _18748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13672__B1 _13557_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14702_ _14702_/A _16433_/A vssd1 vssd1 vccd1 vccd1 _14705_/A sky130_fd_sc_hd__or2_1
XANTENNA__15471__A _15481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18470_ _17281_/X _17913_/Y _18835_/S vssd1 vssd1 vccd1 vccd1 _18470_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11914_ _15505_/A _11913_/Y _11906_/A vssd1 vssd1 vccd1 vccd1 _21013_/D sky130_fd_sc_hd__o21a_1
XFILLER_61_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15682_ _15682_/A vssd1 vssd1 vccd1 vccd1 _15682_/X sky130_fd_sc_hd__buf_1
XPHY_4440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12894_ _12891_/X _20736_/Q _12894_/S vssd1 vssd1 vccd1 vccd1 _20736_/D sky130_fd_sc_hd__mux2_1
XFILLER_73_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17421_ _19295_/Q vssd1 vssd1 vccd1 vccd1 _17421_/Y sky130_fd_sc_hd__inv_2
XPHY_4462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14633_ _14633_/A vssd1 vssd1 vccd1 vccd1 _14636_/B sky130_fd_sc_hd__inv_2
XFILLER_72_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11845_ _11845_/A _11845_/B vssd1 vssd1 vccd1 vccd1 _11845_/X sky130_fd_sc_hd__and2_1
XPHY_4484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output104_A _17483_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17352_ _19319_/Q vssd1 vssd1 vccd1 vccd1 _17352_/Y sky130_fd_sc_hd__inv_2
XPHY_3772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14564_ _14535_/Y _14544_/X _14549_/Y _14555_/Y _14563_/X vssd1 vssd1 vccd1 vccd1
+ _14564_/X sky130_fd_sc_hd__a2111o_1
X_11776_ _16683_/A _11776_/B vssd1 vssd1 vccd1 vccd1 _11776_/X sky130_fd_sc_hd__and2_1
XPHY_3783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16303_ _19387_/Q _16298_/X _16283_/X _16300_/X vssd1 vssd1 vccd1 vccd1 _19387_/D
+ sky130_fd_sc_hd__a22o_1
X_13515_ _13515_/A vssd1 vssd1 vccd1 vccd1 _13515_/X sky130_fd_sc_hd__buf_1
XFILLER_13_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10727_ _10540_/B _10726_/A _21312_/Q _10729_/A _10670_/X vssd1 vssd1 vccd1 vccd1
+ _21312_/D sky130_fd_sc_hd__o221a_1
X_17283_ _20812_/Q vssd1 vssd1 vccd1 vccd1 _17283_/Y sky130_fd_sc_hd__inv_2
X_14495_ _14460_/D _14364_/B _14493_/Y _14488_/X vssd1 vssd1 vccd1 vccd1 _20221_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_158_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_repeater254_A repeater255/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17829__C _18926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19022_ _16903_/X _20401_/Q _19026_/S vssd1 vssd1 vccd1 vccd1 _19954_/D sky130_fd_sc_hd__mux2_1
XFILLER_158_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16234_ _19421_/Q _16230_/X _16231_/X _16233_/X vssd1 vssd1 vccd1 vccd1 _19421_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_146_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13446_ _15424_/A vssd1 vssd1 vccd1 vccd1 _13446_/X sky130_fd_sc_hd__buf_2
XFILLER_70_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10658_ _10658_/A _10687_/A vssd1 vssd1 vccd1 vccd1 _10659_/B sky130_fd_sc_hd__or2_2
XANTENNA__11738__B1 _11736_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18115__B1 _13560_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18006__B _18006_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16165_ _16419_/A _16165_/B _16194_/C vssd1 vssd1 vccd1 vccd1 _16173_/A sky130_fd_sc_hd__or3_4
XANTENNA__18666__A1 _18069_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13377_ _13377_/A vssd1 vssd1 vccd1 vccd1 _13377_/X sky130_fd_sc_hd__buf_1
XFILLER_126_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10589_ _10661_/A _20760_/Q _21331_/Q _10588_/Y vssd1 vssd1 vccd1 vccd1 _10589_/X
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__18721__S _18898_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15116_ _20446_/Q vssd1 vssd1 vccd1 vccd1 _15116_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12328_ _12328_/A _12347_/A vssd1 vssd1 vccd1 vccd1 _12329_/B sky130_fd_sc_hd__or2_2
XANTENNA__17874__C1 _17873_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16096_ _16102_/A vssd1 vssd1 vccd1 vccd1 _16096_/X sky130_fd_sc_hd__buf_1
XFILLER_154_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19924_ _21342_/CLK _19924_/D repeater212/X vssd1 vssd1 vccd1 vccd1 _19924_/Q sky130_fd_sc_hd__dfrtp_1
X_15047_ _20055_/Q vssd1 vssd1 vccd1 vccd1 _15069_/A sky130_fd_sc_hd__inv_2
X_12259_ _20937_/Q vssd1 vssd1 vccd1 vccd1 _12426_/A sky130_fd_sc_hd__inv_2
XFILLER_96_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09644__A input43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19091__A1 _21087_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19855_ _21162_/CLK _19855_/D repeater228/X vssd1 vssd1 vccd1 vccd1 _19855_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__20425__RESET_B repeater270/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15101__B1 _20456_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17861__A _17861_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13166__A _13166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18806_ _18805_/X _10100_/Y _18879_/S vssd1 vssd1 vccd1 vccd1 _18806_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19786_ _19828_/CLK _19786_/D vssd1 vssd1 vccd1 vccd1 _19786_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_228_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16998_ _16998_/A vssd1 vssd1 vccd1 vccd1 _16998_/Y sky130_fd_sc_hd__inv_2
X_18737_ _17610_/Y _10925_/Y _18928_/S vssd1 vssd1 vccd1 vccd1 _18737_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18168__S _18617_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13663__B1 _13538_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15949_ _16340_/A vssd1 vssd1 vccd1 vccd1 _15949_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_92_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18668_ _18845_/A0 _13777_/Y _18896_/S vssd1 vssd1 vccd1 vccd1 _18668_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17619_ _19491_/Q vssd1 vssd1 vccd1 vccd1 _17619_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19682__CLK _19813_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18599_ _18598_/X _10346_/X _18886_/S vssd1 vssd1 vccd1 vccd1 _18599_/X sky130_fd_sc_hd__mux2_1
XFILLER_224_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__21284__RESET_B repeater207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20630_ _20697_/CLK _20630_/D repeater196/X vssd1 vssd1 vccd1 vccd1 _20630_/Q sky130_fd_sc_hd__dfrtp_1
X_20561_ _20592_/CLK _20561_/D repeater260/X vssd1 vssd1 vccd1 vccd1 _20561_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_32_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20492_ _20495_/CLK _20492_/D repeater274/X vssd1 vssd1 vccd1 vccd1 _20492_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_192_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18657__A1 _20030_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14391__B2 _20031_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18631__S _18896_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17865__C1 _17864_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21113_ _21433_/CLK _21113_/D repeater233/X vssd1 vssd1 vccd1 vccd1 _21113_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18409__A1 _21477_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15340__B1 _14258_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12899__B _13261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21044_ _21193_/CLK _21044_/D repeater224/X vssd1 vssd1 vccd1 vccd1 _21044_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09806_ _09806_/A _09806_/B vssd1 vssd1 vccd1 vccd1 _09806_/Y sky130_fd_sc_hd__nor2_1
XFILLER_115_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09737_ _11096_/A _20151_/Q _21231_/Q _20151_/Q vssd1 vssd1 vccd1 vccd1 _09742_/C
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_39_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13654__B1 _13449_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09668_ input67/X vssd1 vssd1 vccd1 vccd1 _15377_/A sky130_fd_sc_hd__buf_1
XPHY_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17396__B2 _17232_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_231_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13406__B1 _13287_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_203_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09599_ _19982_/Q vssd1 vssd1 vccd1 vccd1 _10973_/C sky130_fd_sc_hd__inv_2
XANTENNA__18806__S _18879_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11630_ _14813_/B _11625_/B _11613_/A vssd1 vssd1 vccd1 vccd1 _11631_/B sky130_fd_sc_hd__o21ai_1
XPHY_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18345__A0 _17079_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20828_ _20841_/CLK _20828_/D repeater251/X vssd1 vssd1 vccd1 vccd1 _20828_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11561_ _21131_/Q _11552_/X _11560_/X _11554_/X vssd1 vssd1 vccd1 vccd1 _21131_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20759_ _21477_/CLK _20759_/D repeater201/X vssd1 vssd1 vccd1 vccd1 _20759_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_168_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13300_ _13321_/A vssd1 vssd1 vccd1 vccd1 _13300_/X sky130_fd_sc_hd__buf_1
X_10512_ _20674_/Q vssd1 vssd1 vccd1 vccd1 _17811_/A sky130_fd_sc_hd__inv_2
XFILLER_128_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14280_ _14283_/B vssd1 vssd1 vccd1 vccd1 _14280_/X sky130_fd_sc_hd__buf_1
XPHY_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11492_ _12713_/B vssd1 vssd1 vccd1 vccd1 _13327_/B sky130_fd_sc_hd__buf_1
XFILLER_11_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13231_ _20578_/Q _13226_/X _13146_/X _13228_/X vssd1 vssd1 vccd1 vccd1 _20578_/D
+ sky130_fd_sc_hd__a22o_1
X_10443_ _20673_/Q vssd1 vssd1 vccd1 vccd1 _10443_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18541__S _18784_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13162_ _20604_/Q _13158_/X _12957_/X _13159_/X vssd1 vssd1 vccd1 vccd1 _20604_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_input65_A HWDATA[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10374_ _21371_/Q _10372_/Y _10373_/X _10287_/B vssd1 vssd1 vccd1 vccd1 _21371_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_163_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12113_ _20378_/Q vssd1 vssd1 vccd1 vccd1 _17895_/A sky130_fd_sc_hd__inv_2
XANTENNA__15331__B1 _13553_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17970_ _18207_/X _17926_/X _18181_/X _17927_/X _17969_/X vssd1 vssd1 vccd1 vccd1
+ _17973_/B sky130_fd_sc_hd__o221a_2
XFILLER_124_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13093_ _13099_/A vssd1 vssd1 vccd1 vccd1 _13093_/X sky130_fd_sc_hd__buf_1
XANTENNA__19555__CLK _19706_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19073__A1 _21137_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16921_ _19959_/Q vssd1 vssd1 vccd1 vccd1 _16921_/Y sky130_fd_sc_hd__inv_2
X_12044_ _20951_/Q vssd1 vssd1 vccd1 vccd1 _12305_/A sky130_fd_sc_hd__inv_2
XFILLER_77_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_238_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19640_ _20326_/CLK _19640_/D vssd1 vssd1 vccd1 vccd1 _19640_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16852_ _16856_/B vssd1 vssd1 vccd1 vccd1 _16858_/B sky130_fd_sc_hd__inv_2
XFILLER_77_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15803_ _19629_/Q _15800_/X _09818_/X _15802_/X vssd1 vssd1 vccd1 vccd1 _19629_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_225_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19571_ _19812_/CLK _19571_/D vssd1 vssd1 vccd1 vccd1 _19571_/Q sky130_fd_sc_hd__dfxtp_1
X_16783_ _19926_/Q _16777_/A _16781_/Y _16777_/Y vssd1 vssd1 vccd1 vccd1 _16784_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_18_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13995_ _13971_/B _13887_/B _13993_/Y _13991_/X vssd1 vssd1 vccd1 vccd1 _20311_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_81_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18522_ _17079_/Y _12037_/Y _18908_/S vssd1 vssd1 vccd1 vccd1 _18522_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13714__A _13714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15734_ _19659_/Q _15723_/X _15733_/X _15727_/X vssd1 vssd1 vccd1 vccd1 _19659_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_246_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12946_ _20712_/Q _12942_/X _12697_/X _12943_/X vssd1 vssd1 vccd1 vccd1 _20712_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_206_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15665_ _19690_/Q _15656_/X _15582_/X _15659_/X vssd1 vssd1 vccd1 vccd1 _19690_/D
+ sky130_fd_sc_hd__a22o_1
X_18453_ _18452_/X _10592_/Y _18775_/S vssd1 vssd1 vccd1 vccd1 _18453_/X sky130_fd_sc_hd__mux2_1
X_12877_ _20741_/Q _12874_/X _12875_/X _12876_/X vssd1 vssd1 vccd1 vccd1 _20741_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11671__A2 _11657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18716__S _18896_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14616_ _14616_/A vssd1 vssd1 vccd1 vccd1 _14616_/Y sky130_fd_sc_hd__inv_2
X_17404_ _18804_/X _17324_/X _18813_/X _17326_/X vssd1 vssd1 vccd1 vccd1 _17404_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_21_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18384_ _17079_/Y _12038_/Y _18908_/S vssd1 vssd1 vccd1 vccd1 _18384_/X sky130_fd_sc_hd__mux2_1
X_11828_ _11828_/A vssd1 vssd1 vccd1 vccd1 _11829_/B sky130_fd_sc_hd__inv_2
XFILLER_221_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18336__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15596_ _15603_/A vssd1 vssd1 vccd1 vccd1 _15596_/X sky130_fd_sc_hd__buf_1
XPHY_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17335_ _19424_/Q vssd1 vssd1 vccd1 vccd1 _17335_/Y sky130_fd_sc_hd__inv_2
X_14547_ _20130_/Q vssd1 vssd1 vccd1 vccd1 _14751_/B sky130_fd_sc_hd__inv_2
XFILLER_60_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11759_ _11761_/A _11771_/A vssd1 vssd1 vccd1 vccd1 _11759_/X sky130_fd_sc_hd__or2_1
XFILLER_41_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17266_ _19431_/Q vssd1 vssd1 vccd1 vccd1 _17266_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14478_ _20232_/Q _14476_/Y _14376_/B _14477_/X vssd1 vssd1 vccd1 vccd1 _20232_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA_clkbuf_leaf_41_HCLK_A clkbuf_4_11_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19005_ _16977_/Y _20418_/Q _19019_/S vssd1 vssd1 vccd1 vccd1 _19971_/D sky130_fd_sc_hd__mux2_1
X_16217_ _16223_/A vssd1 vssd1 vccd1 vccd1 _16224_/A sky130_fd_sc_hd__inv_2
XFILLER_174_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13429_ input40/X vssd1 vssd1 vccd1 vccd1 _13429_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__17856__A _17856_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18451__S _18841_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17197_ _18911_/X vssd1 vssd1 vccd1 vccd1 _17197_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20677__RESET_B repeater208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16148_ _19463_/Q _16141_/X _16147_/X _16143_/X vssd1 vssd1 vccd1 vccd1 _19463_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17847__C1 _17843_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15322__B1 _13538_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15376__A _15389_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16079_ _16179_/A _16165_/B _16405_/C vssd1 vssd1 vccd1 vccd1 _16087_/A sky130_fd_sc_hd__or3_4
XFILLER_114_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19907_ _19907_/CLK _19907_/D repeater202/X vssd1 vssd1 vccd1 vccd1 _19907_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_216_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_229_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19838_ _21390_/CLK _19838_/D repeater239/X vssd1 vssd1 vccd1 vccd1 _19838_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_69_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput1 HADDR[0] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_1
XFILLER_68_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13636__B1 _13422_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19769_ _19784_/CLK _19769_/D vssd1 vssd1 vccd1 vccd1 _19769_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_232_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__21465__RESET_B repeater205/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_225_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18626__S _18885_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10870__B1 _09685_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20613_ _20693_/CLK _20613_/D repeater196/X vssd1 vssd1 vccd1 vccd1 _20613_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_138_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20544_ _20724_/CLK _20544_/D repeater264/X vssd1 vssd1 vccd1 vccd1 _20544_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_137_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20475_ _20476_/CLK _20475_/D repeater183/X vssd1 vssd1 vccd1 vccd1 _20475_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18361__S _18667_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15313__A0 _13600_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20555__CLK _20592_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10090_ _20794_/Q vssd1 vssd1 vccd1 vccd1 _10090_/Y sky130_fd_sc_hd__inv_2
XFILLER_102_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19150__S1 _21017_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21027_ _21207_/CLK _21027_/D repeater242/X vssd1 vssd1 vccd1 vccd1 _21027_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_102_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12800_ _20779_/Q _12797_/X _12548_/X _12798_/X vssd1 vssd1 vccd1 vccd1 _20779_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_228_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13780_ _20617_/Q vssd1 vssd1 vccd1 vccd1 _13780_/Y sky130_fd_sc_hd__inv_2
XFILLER_142_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10992_ _10995_/B vssd1 vssd1 vccd1 vccd1 _10992_/X sky130_fd_sc_hd__buf_1
XFILLER_27_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12731_ _20701_/Q vssd1 vssd1 vccd1 vccd1 _12740_/B sky130_fd_sc_hd__buf_1
XFILLER_55_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18536__S _18667_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_243_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15450_ _15657_/A vssd1 vssd1 vccd1 vccd1 _15450_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_187_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12662_ _12679_/A vssd1 vssd1 vccd1 vccd1 _12662_/X sky130_fd_sc_hd__buf_1
XPHY_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14401_ _14401_/A _14401_/B _14401_/C _14400_/X vssd1 vssd1 vccd1 vccd1 _14401_/X
+ sky130_fd_sc_hd__or4b_4
XPHY_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11613_ _11613_/A vssd1 vssd1 vccd1 vccd1 _11623_/B sky130_fd_sc_hd__buf_1
XPHY_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12602__A1 _20872_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15381_ _19821_/Q _15376_/X _15378_/X _15380_/X vssd1 vssd1 vccd1 vccd1 _19821_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18869__A1 _10985_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12602__B2 _12601_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12593_ _20877_/Q _12588_/X _18229_/X _12589_/X vssd1 vssd1 vccd1 vccd1 _20877_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17120_ _19590_/Q vssd1 vssd1 vccd1 vccd1 _17120_/Y sky130_fd_sc_hd__inv_2
XPHY_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14332_ _20231_/Q vssd1 vssd1 vccd1 vccd1 _14333_/A sky130_fd_sc_hd__inv_2
XPHY_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11544_ _11544_/A _11544_/B vssd1 vssd1 vccd1 vccd1 _12501_/B sky130_fd_sc_hd__nand2_1
XFILLER_51_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17051_ _20042_/Q _20040_/Q vssd1 vssd1 vccd1 vccd1 _17051_/X sky130_fd_sc_hd__or2_1
XFILLER_183_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14263_ _20250_/Q _14257_/X _14262_/X _14260_/X vssd1 vssd1 vccd1 vccd1 _20250_/D
+ sky130_fd_sc_hd__a22o_1
X_11475_ _11481_/A vssd1 vssd1 vccd1 vccd1 _11475_/X sky130_fd_sc_hd__buf_1
XANTENNA__18271__S _18880_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16002_ _16010_/A vssd1 vssd1 vccd1 vccd1 _16002_/X sky130_fd_sc_hd__buf_1
X_13214_ _20585_/Q _13206_/X _13213_/X _13207_/X vssd1 vssd1 vccd1 vccd1 _20585_/D
+ sky130_fd_sc_hd__a22o_1
X_10426_ _10762_/A _20674_/Q _10770_/A _20683_/Q vssd1 vssd1 vccd1 vccd1 _10426_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_143_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14194_ _14091_/A _14091_/B _14190_/Y _14193_/X vssd1 vssd1 vccd1 vccd1 _20281_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_3_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13145_ _20613_/Q _13139_/X _13144_/X _13142_/X vssd1 vssd1 vccd1 vccd1 _20613_/D
+ sky130_fd_sc_hd__a22o_1
X_10357_ _20727_/Q vssd1 vssd1 vccd1 vccd1 _18035_/A sky130_fd_sc_hd__inv_2
XFILLER_98_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_repeater217_A repeater218/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17953_ _18538_/X _17951_/X _18542_/X _17952_/X vssd1 vssd1 vccd1 vccd1 _17957_/C
+ sky130_fd_sc_hd__a22o_1
X_13076_ _20651_/Q _13072_/X _12930_/X _13073_/X vssd1 vssd1 vccd1 vccd1 _20651_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_183_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10288_ _10288_/A _10369_/A vssd1 vssd1 vccd1 vccd1 _10289_/B sky130_fd_sc_hd__or2_2
XFILLER_78_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12027_ _19077_/X _12023_/X _20988_/Q _12024_/X vssd1 vssd1 vccd1 vccd1 _20988_/D
+ sky130_fd_sc_hd__a22o_1
X_16904_ _19955_/Q vssd1 vssd1 vccd1 vccd1 _16906_/A sky130_fd_sc_hd__inv_2
XFILLER_239_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17884_ _20824_/Q vssd1 vssd1 vccd1 vccd1 _17884_/Y sky130_fd_sc_hd__inv_2
XFILLER_120_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19623_ _20890_/CLK _19623_/D vssd1 vssd1 vccd1 vccd1 _19623_/Q sky130_fd_sc_hd__dfxtp_1
X_16835_ _16835_/A vssd1 vssd1 vccd1 vccd1 _16877_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__13618__B1 _13557_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13444__A _13444_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19554_ _19706_/CLK _19554_/D vssd1 vssd1 vccd1 vccd1 _19554_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_207_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16766_ _16766_/A _16766_/B vssd1 vssd1 vccd1 vccd1 _16766_/Y sky130_fd_sc_hd__nor2_1
XFILLER_34_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13978_ _20319_/Q _13977_/X _13969_/X _13895_/A vssd1 vssd1 vccd1 vccd1 _20319_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_80_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18505_ _18848_/A0 _10355_/Y _18884_/S vssd1 vssd1 vccd1 vccd1 _18505_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15717_ _15717_/A vssd1 vssd1 vccd1 vccd1 _15717_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_12929_ _20721_/Q _12924_/X _12928_/X _12926_/X vssd1 vssd1 vccd1 vccd1 _20721_/D
+ sky130_fd_sc_hd__a22o_1
X_16697_ _19893_/Q _14233_/B _14234_/B vssd1 vssd1 vccd1 vccd1 _16697_/X sky130_fd_sc_hd__a21bo_1
X_19485_ _19626_/CLK _19485_/D vssd1 vssd1 vccd1 vccd1 _19485_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__18446__S _18884_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18436_ _18435_/X _10132_/Y _18885_/S vssd1 vssd1 vccd1 vccd1 _18436_/X sky130_fd_sc_hd__mux2_1
XANTENNA__18309__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15648_ _15648_/A vssd1 vssd1 vccd1 vccd1 _15648_/X sky130_fd_sc_hd__buf_1
XFILLER_15_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15579_ _19733_/Q _15576_/X _15544_/X _15578_/X vssd1 vssd1 vccd1 vccd1 _19733_/D
+ sky130_fd_sc_hd__a22o_1
X_18367_ _17981_/Y _20758_/Q _18775_/S vssd1 vssd1 vccd1 vccd1 _18367_/X sky130_fd_sc_hd__mux2_1
XANTENNA__20858__RESET_B repeater243/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17318_ _18844_/X _17861_/A _18841_/X _17862_/A _17317_/X vssd1 vssd1 vccd1 vccd1
+ _17318_/X sky130_fd_sc_hd__o221a_1
X_18298_ _18297_/X _10285_/A _18886_/S vssd1 vssd1 vccd1 vccd1 _18298_/X sky130_fd_sc_hd__mux2_1
XFILLER_186_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17249_ _19775_/Q vssd1 vssd1 vccd1 vccd1 _17249_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18181__S _18904_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20260_ _20592_/CLK _20260_/D repeater262/X vssd1 vssd1 vccd1 vccd1 _20260_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_116_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13619__A _13625_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20191_ _20626_/CLK _20191_/D repeater200/X vssd1 vssd1 vccd1 vccd1 _20191_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_89_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19132__S1 _21017_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13609__B1 _13538_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10978__A _12715_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12832__A1 _20764_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_225_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18356__S _18849_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19199__S1 _20131_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20527_ _20946_/CLK _20527_/D repeater275/X vssd1 vssd1 vccd1 vccd1 _20527_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__15534__B1 _15456_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11260_ _20912_/Q vssd1 vssd1 vccd1 vccd1 _11270_/B sky130_fd_sc_hd__inv_2
XANTENNA__20181__RESET_B repeater200/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20458_ _20937_/CLK _20458_/D repeater276/X vssd1 vssd1 vccd1 vccd1 _20458_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_4_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10211_ _21385_/Q _10210_/Y _10207_/B _10140_/X vssd1 vssd1 vccd1 vccd1 _21385_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_106_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11191_ _11192_/A vssd1 vssd1 vccd1 vccd1 _11191_/X sky130_fd_sc_hd__buf_1
X_20389_ _20950_/CLK _20389_/D repeater278/X vssd1 vssd1 vccd1 vccd1 _20389_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_106_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10142_ _10185_/A vssd1 vssd1 vccd1 vccd1 _10177_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__17943__B _17943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14950_ _14950_/A vssd1 vssd1 vccd1 vccd1 _15059_/B sky130_fd_sc_hd__inv_2
X_10073_ _21400_/Q vssd1 vssd1 vccd1 vccd1 _10161_/A sky130_fd_sc_hd__inv_2
XFILLER_48_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21387__RESET_B repeater252/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11323__A1 _21185_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13901_ _13900_/Y _20316_/Q _20659_/Q _13893_/A vssd1 vssd1 vccd1 vccd1 _13901_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_247_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input28_A HADDR[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14881_ _14881_/A _14881_/B _14968_/A vssd1 vssd1 vccd1 vccd1 _14957_/A sky130_fd_sc_hd__or3_1
XFILLER_248_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13832_ _20207_/Q vssd1 vssd1 vccd1 vccd1 _13832_/Y sky130_fd_sc_hd__inv_2
X_16620_ _16620_/A _16620_/B _16620_/C vssd1 vssd1 vccd1 vccd1 _16620_/X sky130_fd_sc_hd__and3_1
XFILLER_235_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18539__A0 _17281_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_150_HCLK clkbuf_opt_1_HCLK/A vssd1 vssd1 vccd1 vccd1 _20137_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_204_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16551_ _21150_/Q vssd1 vssd1 vccd1 vccd1 _16551_/Y sky130_fd_sc_hd__inv_2
XFILLER_204_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13763_ _20601_/Q vssd1 vssd1 vccd1 vccd1 _13763_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10975_ _10975_/A _17315_/A vssd1 vssd1 vccd1 vccd1 _11190_/A sky130_fd_sc_hd__or2_1
XANTENNA__18266__S _18903_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15502_ _19768_/Q _15499_/X _15427_/X _15500_/X vssd1 vssd1 vccd1 vccd1 _19768_/D
+ sky130_fd_sc_hd__a22o_1
X_12714_ _13328_/A _17316_/A vssd1 vssd1 vccd1 vccd1 _13535_/B sky130_fd_sc_hd__or2_2
X_19270_ _17126_/Y _17127_/Y _17128_/Y _17129_/Y _20130_/Q _20131_/Q vssd1 vssd1 vccd1
+ vccd1 _19270_/X sky130_fd_sc_hd__mux4_2
X_16482_ _16482_/A vssd1 vssd1 vccd1 vccd1 _19123_/S sky130_fd_sc_hd__inv_2
X_13694_ _13708_/A vssd1 vssd1 vccd1 vccd1 _13694_/X sky130_fd_sc_hd__buf_1
XFILLER_43_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18221_ _20845_/Q input23/X _18236_/S vssd1 vssd1 vccd1 vccd1 _18221_/X sky130_fd_sc_hd__mux2_4
X_15433_ _15528_/A _15655_/B _15708_/C vssd1 vssd1 vccd1 vccd1 _15441_/A sky130_fd_sc_hd__or3_4
XFILLER_203_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12645_ _14304_/A vssd1 vssd1 vccd1 vccd1 _13328_/A sky130_fd_sc_hd__buf_1
XPHY_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_repeater167_A _18909_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18152_ _18001_/Y _20455_/Q _18784_/S vssd1 vssd1 vccd1 vccd1 _18152_/X sky130_fd_sc_hd__mux2_2
XPHY_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15364_ _19827_/Q _15359_/X _14264_/X _15361_/X vssd1 vssd1 vccd1 vccd1 _19827_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_12_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12576_ _20888_/Q _12574_/X _18240_/X _12575_/X vssd1 vssd1 vccd1 vccd1 _20888_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__20269__RESET_B repeater263/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18711__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19097__S _19870_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14315_ _14315_/A vssd1 vssd1 vccd1 vccd1 _14315_/Y sky130_fd_sc_hd__inv_2
XPHY_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17103_ _19502_/Q vssd1 vssd1 vccd1 vccd1 _17103_/Y sky130_fd_sc_hd__inv_2
X_11527_ _11534_/A vssd1 vssd1 vccd1 vccd1 _11527_/X sky130_fd_sc_hd__buf_1
XPHY_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18083_ _18083_/A _18083_/B vssd1 vssd1 vccd1 vccd1 _18083_/Y sky130_fd_sc_hd__nor2_1
X_15295_ _19861_/Q _15295_/B vssd1 vssd1 vccd1 vccd1 _15296_/B sky130_fd_sc_hd__or2_1
XFILLER_172_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17034_ _17034_/A _17035_/B vssd1 vssd1 vccd1 vccd1 _20018_/D sky130_fd_sc_hd__nor2_1
X_14246_ _14246_/A vssd1 vssd1 vccd1 vccd1 _14246_/X sky130_fd_sc_hd__buf_1
XFILLER_183_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output96_A _18051_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11458_ _21167_/Q _11454_/X _21071_/Q _11457_/X vssd1 vssd1 vccd1 vccd1 _19870_/D
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__13000__A1 _20692_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18014__B _18014_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11011__B1 _21017_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10409_ _10409_/A vssd1 vssd1 vccd1 vccd1 _10409_/Y sky130_fd_sc_hd__inv_2
X_14177_ _14207_/A vssd1 vssd1 vccd1 vccd1 _14215_/B sky130_fd_sc_hd__buf_2
X_11389_ _11389_/A _11389_/B _11389_/C vssd1 vssd1 vccd1 vccd1 _11412_/B sky130_fd_sc_hd__or3_1
XFILLER_113_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13128_ _20622_/Q _13126_/X _13006_/X _13127_/X vssd1 vssd1 vccd1 vccd1 _20622_/D
+ sky130_fd_sc_hd__a22o_1
X_18985_ _11618_/Y _11614_/Y _20015_/Q vssd1 vssd1 vccd1 vccd1 _20015_/D sky130_fd_sc_hd__mux2_1
XFILLER_100_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17936_ _17925_/X _17936_/B _17936_/C vssd1 vssd1 vccd1 vccd1 _17936_/Y sky130_fd_sc_hd__nand3b_4
X_13059_ _20662_/Q _13052_/X _12993_/X _13055_/X vssd1 vssd1 vccd1 vccd1 _20662_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09652__A _12857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_239_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17867_ _20408_/Q vssd1 vssd1 vccd1 vccd1 _17867_/Y sky130_fd_sc_hd__inv_2
Xrepeater148 _18848_/A0 vssd1 vssd1 vccd1 vccd1 _18845_/A0 sky130_fd_sc_hd__clkbuf_16
Xrepeater159 _18850_/S vssd1 vssd1 vccd1 vccd1 _18886_/S sky130_fd_sc_hd__buf_6
X_19606_ _21449_/CLK _19606_/D vssd1 vssd1 vccd1 vccd1 _19606_/Q sky130_fd_sc_hd__dfxtp_1
X_16818_ _16822_/A vssd1 vssd1 vccd1 vccd1 _16818_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17798_ _18672_/X _17472_/X _18671_/X _17474_/X vssd1 vssd1 vccd1 vccd1 _17798_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_207_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19537_ _21462_/CLK _19537_/D vssd1 vssd1 vccd1 vccd1 _19537_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12814__A1 _16779_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16749_ _16758_/A _16749_/B vssd1 vssd1 vccd1 vccd1 _19058_/S sky130_fd_sc_hd__nor2_8
XFILLER_235_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18176__S _18896_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19468_ _20241_/CLK _19468_/D vssd1 vssd1 vccd1 vccd1 _19468_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18419_ _17897_/Y _20648_/Q _18903_/S vssd1 vssd1 vccd1 vccd1 _18419_/X sky130_fd_sc_hd__mux2_1
XFILLER_179_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19399_ _19812_/CLK _19399_/D vssd1 vssd1 vccd1 vccd1 _19399_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__18904__S _18904_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21430_ _21433_/CLK _21430_/D repeater236/X vssd1 vssd1 vccd1 vccd1 _21430_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_147_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21361_ _21367_/CLK _21361_/D repeater254/X vssd1 vssd1 vccd1 vccd1 _21361_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_190_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20312_ _20316_/CLK _20312_/D repeater197/X vssd1 vssd1 vccd1 vccd1 _20312_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__09827__A _09827_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput70 HWRITE vssd1 vssd1 vccd1 vccd1 input70/X sky130_fd_sc_hd__buf_2
XFILLER_116_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21292_ _21357_/CLK _21292_/D repeater199/X vssd1 vssd1 vccd1 vccd1 _21292_/Q sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_31_HCLK clkbuf_opt_4_HCLK/A vssd1 vssd1 vccd1 vccd1 _21120_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_116_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20243_ _21421_/CLK _20243_/D repeater214/X vssd1 vssd1 vccd1 vccd1 _20243_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_171_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20174_ _20241_/CLK _20174_/D repeater249/X vssd1 vssd1 vccd1 vccd1 _20174_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_115_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09985_ _09985_/A vssd1 vssd1 vccd1 vccd1 _09986_/B sky130_fd_sc_hd__inv_2
XANTENNA__18769__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19875__RESET_B repeater226/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_229_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13058__A1 _20663_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14312__A1_N _14275_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10760_ _10760_/A _10760_/B vssd1 vssd1 vccd1 vccd1 _10829_/A sky130_fd_sc_hd__or2_1
XANTENNA__20709__RESET_B repeater210/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10691_ _21327_/Q _10690_/Y _10680_/X _10657_/B vssd1 vssd1 vccd1 vccd1 _21327_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__18814__S _18902_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12430_ _12430_/A _12447_/A vssd1 vssd1 vccd1 vccd1 _12431_/B sky130_fd_sc_hd__or2_1
XFILLER_200_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17938__B _17938_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12361_ _12321_/A _12321_/B _12350_/X _12358_/Y vssd1 vssd1 vccd1 vccd1 _20968_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_165_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14100_ _14100_/A vssd1 vssd1 vccd1 vccd1 _14100_/Y sky130_fd_sc_hd__inv_2
X_11312_ _11312_/A _12503_/B _16568_/B vssd1 vssd1 vccd1 vccd1 _11314_/C sky130_fd_sc_hd__or3_2
XFILLER_165_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15080_ _15129_/A _15080_/B vssd1 vssd1 vccd1 vccd1 _15176_/A sky130_fd_sc_hd__or2_1
XFILLER_4_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12292_ _20923_/Q vssd1 vssd1 vccd1 vccd1 _12471_/A sky130_fd_sc_hd__inv_2
XFILLER_5_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14031_ _14031_/A _14031_/B _14031_/C vssd1 vssd1 vccd1 vccd1 _14034_/A sky130_fd_sc_hd__or3_4
X_11243_ _19910_/Q _11243_/B vssd1 vssd1 vccd1 vccd1 _21194_/D sky130_fd_sc_hd__or2_1
XFILLER_107_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11174_ _15610_/A _11141_/X _11170_/Y _15756_/A _11173_/X vssd1 vssd1 vccd1 vccd1
+ _21222_/D sky130_fd_sc_hd__a32o_1
XFILLER_106_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10125_ _10221_/C _20774_/Q _21381_/Q _10123_/Y _10124_/X vssd1 vssd1 vccd1 vccd1
+ _10125_/X sky130_fd_sc_hd__a221o_1
X_18770_ _18769_/X _16759_/Y _18880_/S vssd1 vssd1 vccd1 vccd1 _18770_/X sky130_fd_sc_hd__mux2_1
X_15982_ _19543_/Q _15978_/X _15949_/X _15979_/X vssd1 vssd1 vccd1 vccd1 _19543_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13297__A1 _20547_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17721_ _20899_/Q vssd1 vssd1 vccd1 vccd1 _17721_/Y sky130_fd_sc_hd__inv_2
XFILLER_236_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14933_ _14933_/A _14933_/B _14933_/C _14933_/D vssd1 vssd1 vccd1 vccd1 _14949_/C
+ sky130_fd_sc_hd__and4_1
X_10056_ _10056_/A vssd1 vssd1 vccd1 vccd1 _10151_/A sky130_fd_sc_hd__buf_1
XANTENNA_output134_A _17042_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11507__A _20251_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17652_ _21191_/Q vssd1 vssd1 vccd1 vccd1 _17652_/Y sky130_fd_sc_hd__inv_2
XFILLER_224_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14864_ _15000_/A _14999_/C _14864_/C _14864_/D vssd1 vssd1 vccd1 vccd1 _14963_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_90_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16603_ _19994_/Q _19991_/Q _16603_/C vssd1 vssd1 vccd1 vccd1 _16603_/X sky130_fd_sc_hd__or3_2
X_13815_ _20196_/Q vssd1 vssd1 vccd1 vccd1 _14585_/A sky130_fd_sc_hd__inv_2
X_14795_ _20118_/Q vssd1 vssd1 vccd1 vccd1 _14795_/Y sky130_fd_sc_hd__inv_2
X_17583_ _17732_/A vssd1 vssd1 vccd1 vccd1 _17821_/A sky130_fd_sc_hd__inv_2
XFILLER_217_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19322_ _19626_/CLK _19322_/D vssd1 vssd1 vccd1 vccd1 _19322_/Q sky130_fd_sc_hd__dfxtp_1
X_16534_ _16556_/A vssd1 vssd1 vccd1 vccd1 _16583_/A sky130_fd_sc_hd__buf_1
X_13746_ _20613_/Q vssd1 vssd1 vccd1 vccd1 _17898_/A sky130_fd_sc_hd__inv_2
XFILLER_31_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19280__S0 _19280_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12272__A2 _20502_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10958_ _21205_/Q vssd1 vssd1 vccd1 vccd1 _10958_/Y sky130_fd_sc_hd__inv_2
XFILLER_189_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18009__B _18084_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19253_ _17334_/Y _17335_/Y _17336_/Y _17337_/Y _19275_/S0 _21004_/Q vssd1 vssd1
+ vccd1 vccd1 _19253_/X sky130_fd_sc_hd__mux4_2
XFILLER_189_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13677_ _20353_/Q _13673_/X _13477_/X _13674_/X vssd1 vssd1 vccd1 vccd1 _20353_/D
+ sky130_fd_sc_hd__a22o_1
X_16465_ _16465_/A _16465_/B _16465_/C vssd1 vssd1 vccd1 vccd1 _16473_/A sky130_fd_sc_hd__or3_4
XFILLER_189_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18724__S _18850_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10889_ _12550_/A vssd1 vssd1 vccd1 vccd1 _10889_/X sky130_fd_sc_hd__buf_2
XFILLER_176_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18204_ _18203_/X _10278_/A _18886_/S vssd1 vssd1 vccd1 vccd1 _18204_/X sky130_fd_sc_hd__mux2_1
XPHY_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12628_ input3/X _12625_/X _20854_/Q _12626_/X vssd1 vssd1 vccd1 vccd1 _20854_/D
+ sky130_fd_sc_hd__o22a_1
X_15416_ _15423_/A vssd1 vssd1 vccd1 vccd1 _15425_/A sky130_fd_sc_hd__inv_2
XFILLER_169_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19184_ _19730_/Q _19370_/Q _19786_/Q _19770_/Q _19280_/S0 _20122_/Q vssd1 vssd1
+ vccd1 vccd1 _19184_/X sky130_fd_sc_hd__mux4_1
X_16396_ _19339_/Q _16392_/X _16235_/X _16394_/X vssd1 vssd1 vccd1 vccd1 _19339_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_54_HCLK clkbuf_4_12_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _21379_/CLK sky130_fd_sc_hd__clkbuf_16
X_15347_ _15347_/A vssd1 vssd1 vccd1 vccd1 _15347_/X sky130_fd_sc_hd__buf_1
X_18135_ _18134_/X _16865_/Y _18667_/S vssd1 vssd1 vccd1 vccd1 _18135_/X sky130_fd_sc_hd__mux2_1
X_12559_ _20892_/Q _12527_/X _12512_/Y vssd1 vssd1 vccd1 vccd1 _20892_/D sky130_fd_sc_hd__o21a_1
XANTENNA__20032__RESET_B repeater205/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10586__A2 _10584_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_184_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15278_ _20478_/Q vssd1 vssd1 vccd1 vccd1 _15278_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18066_ _18284_/X _18048_/X _18135_/X _18065_/X vssd1 vssd1 vccd1 vccd1 _18066_/X
+ sky130_fd_sc_hd__o22a_1
X_17017_ _21269_/Q _09840_/X _09861_/B vssd1 vssd1 vccd1 vccd1 _20004_/D sky130_fd_sc_hd__a21o_4
XANTENNA__13169__A _13710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14229_ _20260_/Q _14228_/Y _14072_/B _14191_/X vssd1 vssd1 vccd1 vccd1 _20260_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_172_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_159_HCLK_A clkbuf_opt_1_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09770_ _09812_/B _09770_/B _16617_/B _14309_/A vssd1 vssd1 vccd1 vccd1 _09771_/D
+ sky130_fd_sc_hd__and4b_1
X_18968_ _11784_/X _11375_/B _21184_/Q vssd1 vssd1 vccd1 vccd1 _18968_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17919_ _17852_/A _17914_/X _17916_/X _17918_/X vssd1 vssd1 vccd1 vccd1 _17919_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_39_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18899_ _17180_/Y _14031_/A _18899_/S vssd1 vssd1 vccd1 vccd1 _18899_/X sky130_fd_sc_hd__mux2_1
XFILLER_226_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20930_ _20930_/CLK _20930_/D repeater268/X vssd1 vssd1 vccd1 vccd1 _20930_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_226_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20766__CLK _21342_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_214_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20861_ _21444_/CLK _20861_/D repeater246/X vssd1 vssd1 vccd1 vccd1 _20861_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_240_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12799__B1 _12544_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_240_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09664__B1 _09663_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19271__S0 _20132_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20792_ _21374_/CLK _20792_/D repeater253/X vssd1 vssd1 vccd1 vccd1 _20792_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__20802__RESET_B repeater252/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18634__S _18896_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11152__A _19986_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21413_ _21417_/CLK _21413_/D repeater234/X vssd1 vssd1 vccd1 vccd1 _21413_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__11223__B1 _10889_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21344_ _21374_/CLK _21344_/D repeater255/X vssd1 vssd1 vccd1 vccd1 _21344_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_118_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21275_ _21462_/CLK _21275_/D repeater245/X vssd1 vssd1 vccd1 vccd1 _21275_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_78_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20226_ _21484_/CLK _20226_/D repeater202/X vssd1 vssd1 vccd1 vccd1 _20226_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_103_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09968_ _09975_/A vssd1 vssd1 vccd1 vccd1 _09968_/X sky130_fd_sc_hd__buf_1
X_20157_ _21242_/CLK _20157_/D repeater189/X vssd1 vssd1 vccd1 vccd1 _20157_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_103_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_18_HCLK_A clkbuf_4_3_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20088_ _20088_/CLK _20088_/D repeater273/X vssd1 vssd1 vccd1 vccd1 _20088_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_100_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09899_ _20007_/Q vssd1 vssd1 vccd1 vccd1 _09899_/X sky130_fd_sc_hd__buf_1
XANTENNA__18809__S _18879_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11930_ _11930_/A vssd1 vssd1 vccd1 vccd1 _19116_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_leaf_6_HCLK_A clkbuf_opt_2_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11861_ _11856_/B _11860_/Y _11803_/X _11852_/X _11805_/A vssd1 vssd1 vccd1 vccd1
+ _11862_/A sky130_fd_sc_hd__o32a_1
XFILLER_150_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13600_ _13600_/A vssd1 vssd1 vccd1 vccd1 _13600_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_214_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10812_ _10812_/A vssd1 vssd1 vccd1 vccd1 _10812_/X sky130_fd_sc_hd__clkbuf_2
XPHY_3932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14580_ _14580_/A _14627_/A vssd1 vssd1 vccd1 vccd1 _14581_/B sky130_fd_sc_hd__or2_2
XFILLER_150_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11792_ _12637_/A vssd1 vssd1 vccd1 vccd1 _12619_/A sky130_fd_sc_hd__buf_1
XANTENNA__19262__S0 _19275_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20543__RESET_B repeater264/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_77_HCLK clkbuf_4_13_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20657_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_3965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13531_ _13528_/A _13530_/A _13175_/A _11974_/X vssd1 vssd1 vccd1 vccd1 _13531_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_213_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10743_ _19933_/Q _19932_/Q _16801_/A vssd1 vssd1 vccd1 vccd1 _16813_/B sky130_fd_sc_hd__or3_4
XPHY_3987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18544__S _18896_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_240_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16250_ _16256_/A vssd1 vssd1 vccd1 vccd1 _16250_/X sky130_fd_sc_hd__buf_1
X_13462_ _20464_/Q _13458_/X _13265_/X _13461_/X vssd1 vssd1 vccd1 vccd1 _20464_/D
+ sky130_fd_sc_hd__a22o_1
X_10674_ _21336_/Q _10669_/C _10670_/X _10672_/A vssd1 vssd1 vccd1 vccd1 _21336_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_174_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15201_ _15201_/A _15201_/B _15201_/C vssd1 vssd1 vccd1 vccd1 _20054_/D sky130_fd_sc_hd__nor3_2
X_12413_ _12445_/A vssd1 vssd1 vccd1 vccd1 _12496_/C sky130_fd_sc_hd__buf_2
X_16181_ _16187_/A vssd1 vssd1 vccd1 vccd1 _16188_/A sky130_fd_sc_hd__inv_2
XFILLER_154_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13393_ _13411_/A vssd1 vssd1 vccd1 vccd1 _13393_/X sky130_fd_sc_hd__buf_1
X_15132_ _20438_/Q vssd1 vssd1 vccd1 vccd1 _15132_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12962__B1 _12875_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12344_ _12359_/A vssd1 vssd1 vccd1 vccd1 _12344_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_175_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15063_ _15128_/A _15063_/B vssd1 vssd1 vccd1 vccd1 _15208_/A sky130_fd_sc_hd__or2_1
X_19940_ _20428_/CLK _19940_/D repeater269/X vssd1 vssd1 vccd1 vccd1 _19940_/Q sky130_fd_sc_hd__dfrtp_1
X_12275_ _20947_/Q vssd1 vssd1 vccd1 vccd1 _12407_/C sky130_fd_sc_hd__inv_2
XANTENNA__15900__B1 _15793_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14014_ _14014_/A _14023_/A vssd1 vssd1 vccd1 vccd1 _14015_/B sky130_fd_sc_hd__or2_2
X_11226_ _11226_/A vssd1 vssd1 vccd1 vccd1 _11226_/X sky130_fd_sc_hd__buf_1
X_19871_ _20042_/CLK _19871_/D repeater219/X vssd1 vssd1 vccd1 vccd1 _19871_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__21331__RESET_B repeater204/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18822_ _18821_/X _12290_/Y _18910_/S vssd1 vssd1 vccd1 vccd1 _18822_/X sky130_fd_sc_hd__mux2_1
XFILLER_150_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11157_ _20429_/Q vssd1 vssd1 vccd1 vccd1 _13527_/A sky130_fd_sc_hd__inv_2
XFILLER_68_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10108_ _21395_/Q _10106_/Y _10156_/A _20792_/Q _10107_/X vssd1 vssd1 vccd1 vccd1
+ _10112_/C sky130_fd_sc_hd__o221a_1
X_18753_ _17539_/Y _20336_/Q _18909_/S vssd1 vssd1 vccd1 vccd1 _18753_/X sky130_fd_sc_hd__mux2_2
X_11088_ _11088_/A vssd1 vssd1 vccd1 vccd1 _21234_/D sky130_fd_sc_hd__inv_2
X_15965_ _19551_/Q _15961_/X _15949_/X _15962_/X vssd1 vssd1 vccd1 vccd1 _19551_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_191_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18719__S _18896_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17704_ _18704_/X _17775_/B vssd1 vssd1 vccd1 vccd1 _17704_/Y sky130_fd_sc_hd__nand2_1
XFILLER_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14916_ _20596_/Q _14885_/Y _20588_/Q _14963_/C vssd1 vssd1 vccd1 vccd1 _14916_/X
+ sky130_fd_sc_hd__o22a_1
X_10039_ _21377_/Q vssd1 vssd1 vccd1 vccd1 _10040_/A sky130_fd_sc_hd__inv_2
XFILLER_236_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18684_ _18683_/X _10081_/Y _18885_/S vssd1 vssd1 vccd1 vccd1 _18684_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13690__A1 _20346_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15896_ _15896_/A vssd1 vssd1 vccd1 vccd1 _15896_/X sky130_fd_sc_hd__buf_1
XANTENNA__09930__A input38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17635_ _20816_/Q vssd1 vssd1 vccd1 vccd1 _17635_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14847_ _20088_/Q vssd1 vssd1 vccd1 vccd1 _14960_/D sky130_fd_sc_hd__inv_2
XFILLER_224_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13452__A _15429_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17566_ _17564_/Y _17639_/A _17565_/Y _17381_/X vssd1 vssd1 vccd1 vccd1 _17566_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__19253__S0 _19275_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14778_ _14779_/A _14318_/X _14777_/X vssd1 vssd1 vccd1 vccd1 _20127_/D sky130_fd_sc_hd__o21ba_1
XANTENNA__20284__RESET_B repeater263/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19305_ _20172_/CLK _19305_/D vssd1 vssd1 vccd1 vccd1 _19305_/Q sky130_fd_sc_hd__dfxtp_1
X_16517_ _19997_/Q vssd1 vssd1 vccd1 vccd1 _16576_/B sky130_fd_sc_hd__inv_2
XFILLER_232_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20213__RESET_B repeater203/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13729_ _20326_/Q vssd1 vssd1 vccd1 vccd1 _15772_/A sky130_fd_sc_hd__buf_1
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17497_ _19778_/Q vssd1 vssd1 vccd1 vccd1 _17497_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18454__S _18617_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19236_ _19232_/X _19233_/X _19234_/X _19235_/X _21005_/Q _21006_/Q vssd1 vssd1 vccd1
+ vccd1 _19236_/X sky130_fd_sc_hd__mux4_2
XFILLER_220_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16448_ _17054_/B vssd1 vssd1 vccd1 vccd1 _17055_/B sky130_fd_sc_hd__inv_2
XFILLER_158_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15379__A _15389_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19167_ _19703_/Q _19567_/Q _19559_/Q _19551_/Q _19280_/S0 _20122_/Q vssd1 vssd1
+ vccd1 vccd1 _19167_/X sky130_fd_sc_hd__mux4_2
XFILLER_192_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16379_ _16385_/A vssd1 vssd1 vccd1 vccd1 _16386_/A sky130_fd_sc_hd__inv_2
XANTENNA__14283__A _20123_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18118_ vssd1 vssd1 vccd1 vccd1 _18118_/HI _18118_/LO sky130_fd_sc_hd__conb_1
XFILLER_129_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19098_ _16672_/X _21080_/Q _19870_/D vssd1 vssd1 vccd1 vccd1 _19098_/X sky130_fd_sc_hd__mux2_1
XFILLER_145_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18049_ _18308_/X _18048_/X _18333_/X _17996_/X vssd1 vssd1 vccd1 vccd1 _18049_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_145_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12705__B1 _12550_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21060_ _21087_/CLK _21060_/D repeater228/X vssd1 vssd1 vccd1 vccd1 _21060_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_160_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09822_ _15871_/A _09813_/X _09821_/X _09815_/X vssd1 vssd1 vccd1 vccd1 _21451_/D
+ sky130_fd_sc_hd__a22o_1
X_20011_ _21438_/CLK _20011_/D repeater237/X vssd1 vssd1 vccd1 vccd1 _20011_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__21001__RESET_B repeater190/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09753_ _21232_/Q vssd1 vssd1 vccd1 vccd1 _11093_/A sky130_fd_sc_hd__inv_2
XFILLER_39_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18629__S _18909_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13130__B1 _12920_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09684_ input64/X vssd1 vssd1 vccd1 vccd1 _10892_/A sky130_fd_sc_hd__buf_2
XFILLER_243_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20913_ _20915_/CLK _20913_/D repeater218/X vssd1 vssd1 vccd1 vccd1 _20913_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__15958__B1 _15891_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20844_ _20857_/CLK _20844_/D repeater243/X vssd1 vssd1 vccd1 vccd1 _20844_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_81_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09637__B1 _09636_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19244__S0 _19275_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18364__S _18891_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20775_ _21379_/CLK _20775_/D repeater213/X vssd1 vssd1 vccd1 vccd1 _20775_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_11_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_6_HCLK clkbuf_opt_2_HCLK/A vssd1 vssd1 vccd1 vccd1 _20326_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__13197__B1 _12989_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12944__B1 _12860_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10390_ _10277_/A _10277_/B _10388_/Y _10383_/X vssd1 vssd1 vccd1 vccd1 _21362_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_136_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21327_ _21477_/CLK _21327_/D repeater201/X vssd1 vssd1 vccd1 vccd1 _21327_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_163_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12060_ _12060_/A _12060_/B _12060_/C _12060_/D vssd1 vssd1 vccd1 vccd1 _12060_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_150_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21258_ _21390_/CLK _21258_/D repeater239/X vssd1 vssd1 vccd1 vccd1 _21258_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_104_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11011_ _21017_/Q _11010_/Y _21017_/Q _11010_/Y vssd1 vssd1 vccd1 vccd1 _11983_/C
+ sky130_fd_sc_hd__a2bb2o_1
X_20209_ _20220_/CLK _20209_/D repeater203/X vssd1 vssd1 vccd1 vccd1 _20209_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__13537__A _13566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21189_ _21191_/CLK _21189_/D repeater224/X vssd1 vssd1 vccd1 vccd1 _21189_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_38_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_142_HCLK_A clkbuf_4_3_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18539__S _18835_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20795__RESET_B repeater252/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15750_ _15750_/A vssd1 vssd1 vccd1 vccd1 _15750_/X sky130_fd_sc_hd__buf_1
X_12962_ _20706_/Q _12960_/X _12875_/X _12961_/X vssd1 vssd1 vccd1 vccd1 _20706_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_246_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20724__RESET_B repeater264/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input10_A HADDR[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14701_ _14730_/B vssd1 vssd1 vccd1 vccd1 _16433_/A sky130_fd_sc_hd__buf_1
X_11913_ _11913_/A _15396_/B vssd1 vssd1 vccd1 vccd1 _11913_/Y sky130_fd_sc_hd__nor2_1
XFILLER_246_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15681_ _15681_/A vssd1 vssd1 vccd1 vccd1 _15681_/X sky130_fd_sc_hd__buf_1
X_12893_ _17087_/A _12899_/A vssd1 vssd1 vccd1 vccd1 _12894_/S sky130_fd_sc_hd__or2_1
XPHY_4430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17420_ _19777_/Q vssd1 vssd1 vccd1 vccd1 _17420_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13272__A input59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14632_ _14577_/A _14577_/B _14621_/X _14630_/Y vssd1 vssd1 vccd1 vccd1 _20188_/D
+ sky130_fd_sc_hd__a211oi_2
X_11844_ _11844_/A vssd1 vssd1 vccd1 vccd1 _21033_/D sky130_fd_sc_hd__inv_2
XFILLER_221_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19235__S0 _19275_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17351_ _19448_/Q vssd1 vssd1 vccd1 vccd1 _17351_/Y sky130_fd_sc_hd__inv_2
X_14563_ _20133_/Q _14562_/X _20133_/Q _14562_/X vssd1 vssd1 vccd1 vccd1 _14563_/X
+ sky130_fd_sc_hd__a2bb2o_1
XPHY_3773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11775_ _19090_/X _11770_/X _21044_/Q _11771_/X vssd1 vssd1 vccd1 vccd1 _21044_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18274__S _18907_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16302_ _19388_/Q _16298_/X _16281_/X _16300_/X vssd1 vssd1 vccd1 vccd1 _19388_/D
+ sky130_fd_sc_hd__a22o_1
X_10726_ _10726_/A vssd1 vssd1 vccd1 vccd1 _10729_/A sky130_fd_sc_hd__inv_2
X_13514_ _13514_/A vssd1 vssd1 vccd1 vccd1 _13514_/X sky130_fd_sc_hd__buf_1
X_14494_ _20222_/Q _14493_/Y _14472_/X _14366_/B vssd1 vssd1 vccd1 vccd1 _20222_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_202_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17282_ _20774_/Q vssd1 vssd1 vccd1 vccd1 _17282_/Y sky130_fd_sc_hd__inv_2
X_19021_ _16907_/X _20402_/Q _19026_/S vssd1 vssd1 vccd1 vccd1 _19955_/D sky130_fd_sc_hd__mux2_1
XFILLER_146_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16233_ _16241_/A vssd1 vssd1 vccd1 vccd1 _16233_/X sky130_fd_sc_hd__buf_1
X_13445_ input63/X vssd1 vssd1 vccd1 vccd1 _15424_/A sky130_fd_sc_hd__clkbuf_2
X_10657_ _10657_/A _10657_/B vssd1 vssd1 vccd1 vccd1 _10687_/A sky130_fd_sc_hd__or2_1
XANTENNA__18115__A1 _21486_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11738__A1 _21059_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater247_A repeater248/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11520__A _15354_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16164_ _19454_/Q _16158_/X _16163_/X _16159_/X vssd1 vssd1 vccd1 vccd1 _19454_/D
+ sky130_fd_sc_hd__a22o_1
X_13376_ _20502_/Q _13371_/X _13163_/X _13372_/X vssd1 vssd1 vccd1 vccd1 _20502_/D
+ sky130_fd_sc_hd__a22o_1
X_10588_ _20759_/Q vssd1 vssd1 vccd1 vccd1 _10588_/Y sky130_fd_sc_hd__inv_2
X_15115_ _20435_/Q vssd1 vssd1 vccd1 vccd1 _15115_/Y sky130_fd_sc_hd__inv_2
X_12327_ _12327_/A _12327_/B vssd1 vssd1 vccd1 vccd1 _12347_/A sky130_fd_sc_hd__or2_1
XANTENNA__19978__RESET_B repeater270/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16095_ _16101_/A vssd1 vssd1 vccd1 vccd1 _16102_/A sky130_fd_sc_hd__inv_2
XANTENNA__15927__A _15927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19907__RESET_B repeater202/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19923_ _21319_/CLK _19923_/D repeater191/X vssd1 vssd1 vccd1 vccd1 _19923_/Q sky130_fd_sc_hd__dfrtp_1
X_15046_ _20056_/Q vssd1 vssd1 vccd1 vccd1 _15070_/A sky130_fd_sc_hd__inv_2
X_12258_ _12258_/A vssd1 vssd1 vccd1 vccd1 _12427_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_79_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13447__A _13447_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11209_ _21212_/Q _11206_/X _09641_/X _11208_/X vssd1 vssd1 vccd1 vccd1 _21212_/D
+ sky130_fd_sc_hd__a22o_1
X_19854_ _21429_/CLK _19854_/D repeater228/X vssd1 vssd1 vccd1 vccd1 _19854_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_123_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12189_ _20959_/Q _12186_/Y _12326_/A _20355_/Q _12188_/X vssd1 vssd1 vccd1 vccd1
+ _12190_/D sky130_fd_sc_hd__o221a_1
XFILLER_69_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18805_ _18845_/A0 _10308_/Y _18884_/S vssd1 vssd1 vccd1 vccd1 _18805_/X sky130_fd_sc_hd__mux2_1
X_19785_ _19835_/CLK _19785_/D vssd1 vssd1 vccd1 vccd1 _19785_/Q sky130_fd_sc_hd__dfxtp_1
X_16997_ _19976_/Q _16997_/B vssd1 vssd1 vccd1 vccd1 _16998_/A sky130_fd_sc_hd__or2_1
XFILLER_84_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18449__S _18884_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16758__A _16758_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18736_ _17631_/X _19338_/Q _18926_/S vssd1 vssd1 vccd1 vccd1 _18736_/X sky130_fd_sc_hd__mux2_1
X_15948_ _19560_/Q _15943_/X _15947_/X _15945_/X vssd1 vssd1 vccd1 vccd1 _19560_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_225_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17929__B2 _17214_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_64_HCLK_A clkbuf_4_11_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18667_ _18666_/X _10287_/A _18667_/S vssd1 vssd1 vccd1 vccd1 _18667_/X sky130_fd_sc_hd__mux2_1
X_15879_ _15879_/A vssd1 vssd1 vccd1 vccd1 _15879_/X sky130_fd_sc_hd__buf_1
XFILLER_236_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17618_ _19579_/Q vssd1 vssd1 vccd1 vccd1 _17618_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12218__A2 _20499_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13415__A1 _20481_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19226__S0 _21005_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18598_ _18597_/X _10103_/Y _18644_/S vssd1 vssd1 vccd1 vccd1 _18598_/X sky130_fd_sc_hd__mux2_1
XFILLER_211_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17549_ _17549_/A vssd1 vssd1 vccd1 vccd1 _17550_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_211_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18184__S _18903_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20560_ _20592_/CLK _20560_/D repeater260/X vssd1 vssd1 vccd1 vccd1 _20560_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_138_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19219_ _17619_/Y _17620_/Y _17621_/Y _17622_/Y _20130_/Q _20131_/Q vssd1 vssd1 vccd1
+ vccd1 _19219_/X sky130_fd_sc_hd__mux4_1
XFILLER_149_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20491_ _20944_/CLK _20491_/D repeater274/X vssd1 vssd1 vccd1 vccd1 _20491_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_118_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21112_ _21417_/CLK _21112_/D repeater234/X vssd1 vssd1 vccd1 vccd1 _21112_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_133_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21043_ _21183_/CLK _21043_/D repeater219/X vssd1 vssd1 vccd1 vccd1 _21043_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA__13357__A _13357_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09805_ _09793_/C _09804_/X _09800_/Y vssd1 vssd1 vccd1 vccd1 _21456_/D sky130_fd_sc_hd__a21oi_1
XANTENNA_input2_A HADDR[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18359__S _18875_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13103__B1 _12884_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09736_ _21231_/Q vssd1 vssd1 vccd1 vccd1 _11096_/A sky130_fd_sc_hd__buf_1
XFILLER_86_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09667_ _21471_/Q _09657_/X _09666_/X _09660_/X vssd1 vssd1 vccd1 vccd1 _21471_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__20135__RESET_B repeater248/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_243_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19217__S0 _20130_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09598_ _20887_/Q vssd1 vssd1 vccd1 vccd1 _09937_/B sky130_fd_sc_hd__inv_2
XPHY_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20827_ _20841_/CLK _20827_/D repeater251/X vssd1 vssd1 vccd1 vccd1 _20827_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11560_ _13163_/A vssd1 vssd1 vccd1 vccd1 _11560_/X sky130_fd_sc_hd__buf_1
XFILLER_51_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20758_ _21477_/CLK _20758_/D repeater201/X vssd1 vssd1 vccd1 vccd1 _20758_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_168_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10511_ _21293_/Q vssd1 vssd1 vccd1 vccd1 _10769_/A sky130_fd_sc_hd__inv_2
XPHY_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11491_ _20889_/Q vssd1 vssd1 vccd1 vccd1 _12713_/B sky130_fd_sc_hd__inv_2
X_20689_ _21302_/CLK _20689_/D repeater209/X vssd1 vssd1 vccd1 vccd1 _20689_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18822__S _18910_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13230_ _20579_/Q _13226_/X _13144_/X _13228_/X vssd1 vssd1 vccd1 vccd1 _20579_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12917__B1 _12673_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10442_ _21306_/Q vssd1 vssd1 vccd1 vccd1 _10782_/A sky130_fd_sc_hd__inv_2
XFILLER_40_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_107_HCLK clkbuf_opt_3_HCLK/A vssd1 vssd1 vccd1 vccd1 _20495_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__17946__B _18007_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13161_ _20605_/Q _13158_/X _12954_/X _13159_/X vssd1 vssd1 vccd1 vccd1 _20605_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13590__B1 _13506_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10373_ _10381_/A vssd1 vssd1 vccd1 vccd1 _10373_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_123_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12112_ _20961_/Q vssd1 vssd1 vccd1 vccd1 _12314_/A sky130_fd_sc_hd__inv_2
XANTENNA_input58_A HWDATA[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13092_ _13098_/A vssd1 vssd1 vccd1 vccd1 _13092_/X sky130_fd_sc_hd__buf_1
XANTENNA__20976__RESET_B repeater278/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13342__B1 _13280_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16920_ _16956_/A _16920_/B vssd1 vssd1 vccd1 vccd1 _16920_/Y sky130_fd_sc_hd__nor2_1
X_12043_ _20978_/Q vssd1 vssd1 vccd1 vccd1 _12331_/A sky130_fd_sc_hd__inv_2
XFILLER_78_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20905__RESET_B repeater217/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16851_ _19942_/Q _16853_/B vssd1 vssd1 vccd1 vccd1 _16856_/B sky130_fd_sc_hd__or2_1
XFILLER_66_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18269__S _18850_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15802_ _15808_/A vssd1 vssd1 vccd1 vccd1 _15802_/X sky130_fd_sc_hd__clkbuf_2
X_19570_ _19812_/CLK _19570_/D vssd1 vssd1 vccd1 vccd1 _19570_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16782_ _16835_/A vssd1 vssd1 vccd1 vccd1 _16820_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_207_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13994_ _20312_/Q _13993_/Y _13969_/X _13889_/B vssd1 vssd1 vccd1 vccd1 _20312_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_74_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18521_ _17946_/Y _16954_/Y _18680_/S vssd1 vssd1 vccd1 vccd1 _18521_/X sky130_fd_sc_hd__mux2_2
X_15733_ _16237_/A vssd1 vssd1 vccd1 vccd1 _15733_/X sky130_fd_sc_hd__buf_1
X_12945_ _20713_/Q _12942_/X _12863_/X _12943_/X vssd1 vssd1 vccd1 vccd1 _20713_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_218_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11515__A input49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18452_ _18845_/A0 _10450_/Y _18884_/S vssd1 vssd1 vccd1 vccd1 _18452_/X sky130_fd_sc_hd__mux2_1
XFILLER_233_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19208__S0 _20130_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15664_ _19691_/Q _15656_/X _15663_/X _15659_/X vssd1 vssd1 vccd1 vccd1 _19691_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12876_ _12876_/A vssd1 vssd1 vccd1 vccd1 _12876_/X sky130_fd_sc_hd__buf_1
XFILLER_60_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17403_ _18816_/X _17211_/A _18819_/X _17319_/X _17402_/X vssd1 vssd1 vccd1 vccd1
+ _17403_/X sky130_fd_sc_hd__o221a_2
XFILLER_233_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14615_ _14587_/A _14587_/B _14607_/X _14613_/Y vssd1 vssd1 vccd1 vccd1 _20198_/D
+ sky130_fd_sc_hd__a211oi_2
XPHY_4293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18383_ _18382_/X _12273_/Y _18910_/S vssd1 vssd1 vccd1 vccd1 _18383_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11827_ _11827_/A vssd1 vssd1 vccd1 vccd1 _11827_/X sky130_fd_sc_hd__buf_1
X_15595_ _15610_/A _15756_/B _16261_/C vssd1 vssd1 vccd1 vccd1 _15603_/A sky130_fd_sc_hd__or3_4
XFILLER_199_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17334_ _19360_/Q vssd1 vssd1 vccd1 vccd1 _17334_/Y sky130_fd_sc_hd__inv_2
X_11758_ _11770_/A vssd1 vssd1 vccd1 vccd1 _11771_/A sky130_fd_sc_hd__inv_2
X_14546_ _15832_/B vssd1 vssd1 vccd1 vccd1 _14747_/B sky130_fd_sc_hd__buf_1
XFILLER_186_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10709_ _21321_/Q _10708_/Y _10712_/A _10651_/B vssd1 vssd1 vccd1 vccd1 _21321_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17265_ _19487_/Q vssd1 vssd1 vccd1 vccd1 _17265_/Y sky130_fd_sc_hd__inv_2
X_14477_ _14477_/A vssd1 vssd1 vccd1 vccd1 _14477_/X sky130_fd_sc_hd__clkbuf_2
X_11689_ _11689_/A vssd1 vssd1 vccd1 vccd1 _11689_/X sky130_fd_sc_hd__buf_1
X_19004_ _16982_/X _20419_/Q _19019_/S vssd1 vssd1 vccd1 vccd1 _19972_/D sky130_fd_sc_hd__mux2_1
XANTENNA__12908__B1 _12660_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16216_ _16223_/A vssd1 vssd1 vccd1 vccd1 _16216_/X sky130_fd_sc_hd__clkbuf_2
X_13428_ _13444_/A vssd1 vssd1 vccd1 vccd1 _13428_/X sky130_fd_sc_hd__buf_1
X_17196_ _17472_/A vssd1 vssd1 vccd1 vccd1 _17196_/X sky130_fd_sc_hd__buf_1
XFILLER_161_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16147_ _21447_/Q vssd1 vssd1 vccd1 vccd1 _16147_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15657__A _15657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13359_ _13359_/A vssd1 vssd1 vccd1 vccd1 _13378_/A sky130_fd_sc_hd__buf_1
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09655__A _12860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16078_ _16405_/A vssd1 vssd1 vccd1 vccd1 _16179_/A sky130_fd_sc_hd__buf_1
XFILLER_170_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19906_ _19907_/CLK input78/X repeater202/X vssd1 vssd1 vccd1 vccd1 _19907_/D sky130_fd_sc_hd__dfrtp_1
X_15029_ _15029_/A vssd1 vssd1 vccd1 vccd1 _15087_/A sky130_fd_sc_hd__inv_2
XFILLER_229_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19997__SET_B repeater220/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18272__A0 _17079_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_229_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19837_ _20172_/CLK _19837_/D vssd1 vssd1 vccd1 vccd1 _19837_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18179__S _18902_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput2 HADDR[10] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_1
X_19768_ _19784_/CLK _19768_/D vssd1 vssd1 vccd1 vccd1 _19768_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_232_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18719_ _18845_/A0 _13793_/Y _18896_/S vssd1 vssd1 vccd1 vccd1 _18719_/X sky130_fd_sc_hd__mux2_1
X_19699_ _21009_/CLK _19699_/D vssd1 vssd1 vccd1 vccd1 _19699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_232_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18907__S _18907_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_225_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20612_ _20657_/CLK _20612_/D repeater195/X vssd1 vssd1 vccd1 vccd1 _20612_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_178_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20543_ _20724_/CLK _20543_/D repeater264/X vssd1 vssd1 vccd1 vccd1 _20543_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18642__S _18907_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20474_ _20476_/CLK _20474_/D repeater280/X vssd1 vssd1 vccd1 vccd1 _20474_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_133_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13324__B1 _13169_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21282__CLK _21342_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21026_ _21255_/CLK _21026_/D repeater241/X vssd1 vssd1 vccd1 vccd1 _21026_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_101_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20316__RESET_B repeater262/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09719_ _20157_/Q vssd1 vssd1 vccd1 vccd1 _09719_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10991_ _10991_/A _10991_/B vssd1 vssd1 vccd1 vccd1 _10995_/B sky130_fd_sc_hd__nor2_1
XFILLER_215_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18817__S _18908_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10877__C _12605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12730_ _20702_/Q vssd1 vssd1 vccd1 vccd1 _14686_/A sky130_fd_sc_hd__buf_1
XFILLER_243_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_230_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12661_ _20839_/Q _12650_/X _12660_/X _12654_/X vssd1 vssd1 vccd1 vccd1 _20839_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14400_ _21469_/Q _14500_/A _21483_/Q _14460_/B vssd1 vssd1 vccd1 vccd1 _14400_/X
+ sky130_fd_sc_hd__o22a_1
X_11612_ _20015_/Q vssd1 vssd1 vccd1 vccd1 _11613_/A sky130_fd_sc_hd__buf_1
XPHY_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13550__A input57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21175__RESET_B repeater216/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12592_ _20878_/Q _12588_/X _18230_/X _12589_/X vssd1 vssd1 vccd1 vccd1 _20878_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_42_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16329__B1 _16231_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15380_ _15390_/A vssd1 vssd1 vccd1 vccd1 _15380_/X sky130_fd_sc_hd__buf_1
XPHY_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12602__A2 _12600_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11543_ _11543_/A _20902_/Q _11543_/C _11307_/C vssd1 vssd1 vccd1 vccd1 _11544_/B
+ sky130_fd_sc_hd__or4b_4
X_14331_ _20232_/Q vssd1 vssd1 vccd1 vccd1 _14463_/C sky130_fd_sc_hd__inv_2
XPHY_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18552__S _18841_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17050_ _20039_/Q _20037_/Q _20038_/Q _17049_/X vssd1 vssd1 vccd1 vccd1 _19848_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14262_ _14262_/A vssd1 vssd1 vccd1 vccd1 _14262_/X sky130_fd_sc_hd__clkbuf_4
X_11474_ _11480_/A vssd1 vssd1 vccd1 vccd1 _11474_/X sky130_fd_sc_hd__buf_1
XFILLER_183_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16001_ _16008_/A vssd1 vssd1 vccd1 vccd1 _16010_/A sky130_fd_sc_hd__inv_2
X_13213_ input50/X vssd1 vssd1 vccd1 vccd1 _13213_/X sky130_fd_sc_hd__clkbuf_2
X_10425_ _21294_/Q vssd1 vssd1 vccd1 vccd1 _10770_/A sky130_fd_sc_hd__inv_2
XANTENNA__15477__A _15766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14193_ _14207_/A vssd1 vssd1 vccd1 vccd1 _14193_/X sky130_fd_sc_hd__buf_2
XFILLER_152_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13144_ input43/X vssd1 vssd1 vccd1 vccd1 _13144_/X sky130_fd_sc_hd__clkbuf_4
X_10356_ _20734_/Q vssd1 vssd1 vccd1 vccd1 _10356_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15304__B2 _18962_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14512__C1 _14469_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17952_ _17952_/A vssd1 vssd1 vccd1 vccd1 _17952_/X sky130_fd_sc_hd__buf_1
XFILLER_97_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13075_ _20652_/Q _13072_/X _12928_/X _13073_/X vssd1 vssd1 vccd1 vccd1 _20652_/D
+ sky130_fd_sc_hd__a22o_1
X_10287_ _10287_/A _10287_/B vssd1 vssd1 vccd1 vccd1 _10369_/A sky130_fd_sc_hd__or2_1
XFILLER_78_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12026_ _19076_/X _12023_/X _20989_/Q _12024_/X vssd1 vssd1 vccd1 vccd1 _20989_/D
+ sky130_fd_sc_hd__a22o_1
X_16903_ _16906_/B _16902_/Y _16898_/X vssd1 vssd1 vccd1 vccd1 _16903_/X sky130_fd_sc_hd__o21a_1
XFILLER_239_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20057__RESET_B repeater281/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17883_ _17852_/X _17878_/X _17880_/X _17882_/X vssd1 vssd1 vccd1 vccd1 _17883_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_239_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19622_ _21449_/CLK _19622_/D vssd1 vssd1 vccd1 vccd1 _19622_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16834_ _16834_/A vssd1 vssd1 vccd1 vccd1 _16834_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19553_ _19706_/CLK _19553_/D vssd1 vssd1 vccd1 vccd1 _19553_/Q sky130_fd_sc_hd__dfxtp_1
X_16765_ _16765_/A vssd1 vssd1 vccd1 vccd1 _16770_/B sky130_fd_sc_hd__inv_2
XANTENNA__18727__S _18907_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13977_ _20318_/Q _20317_/Q _13977_/C vssd1 vssd1 vccd1 vccd1 _13977_/X sky130_fd_sc_hd__and3_1
XFILLER_207_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18504_ _18503_/X _10769_/A _18617_/S vssd1 vssd1 vccd1 vccd1 _18504_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15716_ _15716_/A vssd1 vssd1 vccd1 vccd1 _15716_/X sky130_fd_sc_hd__buf_1
X_19484_ _19626_/CLK _19484_/D vssd1 vssd1 vccd1 vccd1 _19484_/Q sky130_fd_sc_hd__dfxtp_1
X_12928_ input47/X vssd1 vssd1 vccd1 vccd1 _12928_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__21005__CLK _21009_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16696_ _16700_/A _18944_/X vssd1 vssd1 vccd1 vccd1 _19892_/D sky130_fd_sc_hd__and2_1
XFILLER_61_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18435_ _18845_/A0 _10309_/Y _18884_/S vssd1 vssd1 vccd1 vccd1 _18435_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15647_ _15647_/A vssd1 vssd1 vccd1 vccd1 _15647_/X sky130_fd_sc_hd__buf_1
XPHY_4090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12859_ _12874_/A vssd1 vssd1 vccd1 vccd1 _12859_/X sky130_fd_sc_hd__buf_1
XFILLER_33_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18366_ _17983_/Y _16834_/Y _18875_/S vssd1 vssd1 vccd1 vccd1 _18366_/X sky130_fd_sc_hd__mux2_1
XFILLER_159_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15578_ _15586_/A vssd1 vssd1 vccd1 vccd1 _15578_/X sky130_fd_sc_hd__buf_1
XFILLER_30_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17317_ _18870_/X _17315_/X _18836_/X _17844_/A vssd1 vssd1 vccd1 vccd1 _17317_/X
+ sky130_fd_sc_hd__o22a_2
X_14529_ _16617_/B _14529_/B vssd1 vssd1 vccd1 vccd1 _16618_/A sky130_fd_sc_hd__nand2_1
XFILLER_174_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18462__S _18775_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18297_ _18296_/X _10093_/Y _18644_/S vssd1 vssd1 vccd1 vccd1 _18297_/X sky130_fd_sc_hd__mux2_1
XFILLER_175_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19922__RESET_B repeater212/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17248_ _19711_/Q vssd1 vssd1 vccd1 vccd1 _17248_/Y sky130_fd_sc_hd__inv_2
XFILLER_147_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13554__B1 _13553_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17179_ _17193_/B vssd1 vssd1 vccd1 vccd1 _17187_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__20827__RESET_B repeater251/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12804__A _12804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18493__A0 _17079_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20190_ _20626_/CLK _20190_/D repeater200/X vssd1 vssd1 vccd1 vccd1 _20190_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_143_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13306__B1 _13148_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13609__A1 _20395_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10978__B _15884_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18637__S _18902_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17220__A1 _18930_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18372__S _18910_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16681__A _21088_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20526_ _20946_/CLK _20526_/D repeater274/X vssd1 vssd1 vccd1 vccd1 _20526_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_153_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20457_ _20495_/CLK _20457_/D repeater276/X vssd1 vssd1 vccd1 vccd1 _20457_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__18484__A0 _17079_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10210_ _10210_/A vssd1 vssd1 vccd1 vccd1 _10210_/Y sky130_fd_sc_hd__inv_2
XFILLER_180_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11190_ _11190_/A _16487_/A vssd1 vssd1 vccd1 vccd1 _11192_/A sky130_fd_sc_hd__or2_2
X_20388_ _20980_/CLK _20388_/D repeater278/X vssd1 vssd1 vccd1 vccd1 _20388_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_79_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10141_ _21407_/Q _10147_/A _10079_/Y _10078_/A _10140_/X vssd1 vssd1 vccd1 vccd1
+ _21407_/D sky130_fd_sc_hd__o221a_1
XFILLER_88_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10072_ _21401_/Q vssd1 vssd1 vccd1 vccd1 _10162_/A sky130_fd_sc_hd__inv_2
XANTENNA__20150__RESET_B repeater250/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13545__A input59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21009_ _21009_/CLK _21009_/D repeater235/X vssd1 vssd1 vccd1 vccd1 _21009_/Q sky130_fd_sc_hd__dfrtp_1
X_13900_ _20659_/Q vssd1 vssd1 vccd1 vccd1 _13900_/Y sky130_fd_sc_hd__inv_2
XFILLER_208_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14880_ _14880_/A _14880_/B vssd1 vssd1 vccd1 vccd1 _14968_/A sky130_fd_sc_hd__or2_1
XFILLER_87_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13831_ _20192_/Q vssd1 vssd1 vccd1 vccd1 _14581_/A sky130_fd_sc_hd__inv_2
XFILLER_46_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18547__S _18902_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_216_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16550_ _21148_/Q vssd1 vssd1 vccd1 vccd1 _16550_/Y sky130_fd_sc_hd__inv_2
XFILLER_189_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13762_ _20178_/Q vssd1 vssd1 vccd1 vccd1 _14568_/A sky130_fd_sc_hd__inv_2
X_10974_ _20890_/Q _20889_/Q _13047_/C vssd1 vssd1 vccd1 vccd1 _17315_/A sky130_fd_sc_hd__or3_4
XANTENNA__21356__RESET_B repeater254/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15501_ _19769_/Q _15499_/X _15424_/X _15500_/X vssd1 vssd1 vccd1 vccd1 _19769_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_189_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12713_ _12753_/A _12713_/B _14303_/C vssd1 vssd1 vccd1 vccd1 _17316_/A sky130_fd_sc_hd__or3_1
X_16481_ _16481_/A _16481_/B vssd1 vssd1 vccd1 vccd1 _16481_/Y sky130_fd_sc_hd__nor2_1
XFILLER_188_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13693_ _13706_/A vssd1 vssd1 vccd1 vccd1 _13693_/X sky130_fd_sc_hd__buf_1
XFILLER_204_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18220_ _20844_/Q input12/X _18236_/S vssd1 vssd1 vccd1 vccd1 _18220_/X sky130_fd_sc_hd__mux2_2
XANTENNA__13280__A input56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15432_ _19798_/Q _15423_/X _15431_/X _15425_/X vssd1 vssd1 vccd1 vccd1 _19798_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12644_ _13046_/A vssd1 vssd1 vccd1 vccd1 _17083_/A sky130_fd_sc_hd__buf_2
XPHY_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18151_ _18150_/X _16975_/Y _18680_/S vssd1 vssd1 vccd1 vccd1 _18151_/X sky130_fd_sc_hd__mux2_1
XPHY_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12575_ _12575_/A vssd1 vssd1 vccd1 vccd1 _12575_/X sky130_fd_sc_hd__buf_1
X_15363_ _19828_/Q _15359_/X _14262_/X _15361_/X vssd1 vssd1 vccd1 vccd1 _19828_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18282__S _18884_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17102_ _19382_/Q vssd1 vssd1 vccd1 vccd1 _17102_/Y sky130_fd_sc_hd__inv_2
XFILLER_184_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14314_ _15335_/B _20121_/Q _14779_/B _14288_/X _19120_/X vssd1 vssd1 vccd1 vccd1
+ _14324_/B sky130_fd_sc_hd__o221ai_1
X_11526_ _11678_/A _14273_/D vssd1 vssd1 vccd1 vccd1 _11534_/A sky130_fd_sc_hd__or2_2
X_18082_ _18082_/A _18083_/B vssd1 vssd1 vccd1 vccd1 _18082_/Y sky130_fd_sc_hd__nor2_1
XPHY_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15294_ _19860_/Q _15294_/B vssd1 vssd1 vccd1 vccd1 _15295_/B sky130_fd_sc_hd__or2_1
XPHY_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17033_ _17033_/A _17035_/B vssd1 vssd1 vccd1 vccd1 _20017_/D sky130_fd_sc_hd__nor2_1
X_14245_ _14249_/A vssd1 vssd1 vccd1 vccd1 _18946_/S sky130_fd_sc_hd__buf_8
X_11457_ _11457_/A _19850_/D _11457_/C vssd1 vssd1 vccd1 vccd1 _11457_/X sky130_fd_sc_hd__or3_4
XFILLER_183_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10408_ _10268_/A _10268_/B _10406_/Y _10397_/X vssd1 vssd1 vccd1 vccd1 _21352_/D
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__18475__A0 _18848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14176_ _14176_/A vssd1 vssd1 vccd1 vccd1 _14207_/A sky130_fd_sc_hd__buf_1
X_11388_ _11388_/A _11388_/B _11386_/B vssd1 vssd1 vccd1 vccd1 _11389_/C sky130_fd_sc_hd__nor3b_4
XANTENNA_output89_A _17973_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20238__RESET_B repeater205/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13127_ _13133_/A vssd1 vssd1 vccd1 vccd1 _13127_/X sky130_fd_sc_hd__buf_1
XANTENNA__15935__A _15943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10339_ _21354_/Q _10336_/Y _10264_/A _20707_/Q _10338_/X vssd1 vssd1 vccd1 vccd1
+ _10340_/D sky130_fd_sc_hd__o221a_1
X_18984_ _21412_/Q _17039_/Y _18984_/S vssd1 vssd1 vccd1 vccd1 _18984_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17935_ _18444_/X _17931_/X _18540_/X _17932_/X _17934_/X vssd1 vssd1 vccd1 vccd1
+ _17936_/C sky130_fd_sc_hd__o221a_1
X_13058_ _20663_/Q _13052_/X _12991_/X _13055_/X vssd1 vssd1 vccd1 vccd1 _20663_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09933__A _14304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18030__B _18032_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12009_ _12011_/A vssd1 vssd1 vccd1 vccd1 _12029_/A sky130_fd_sc_hd__buf_1
XFILLER_38_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17866_ _20822_/Q vssd1 vssd1 vccd1 vccd1 _17866_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater149 _17281_/X vssd1 vssd1 vccd1 vccd1 _18848_/A0 sky130_fd_sc_hd__clkbuf_16
XFILLER_226_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16817_ _19935_/Q vssd1 vssd1 vccd1 vccd1 _16822_/A sky130_fd_sc_hd__buf_1
X_19605_ _20142_/CLK _19605_/D vssd1 vssd1 vccd1 vccd1 _19605_/Q sky130_fd_sc_hd__dfxtp_1
X_17797_ _16566_/A _17550_/X _17791_/X _17796_/X vssd1 vssd1 vccd1 vccd1 _17797_/X
+ sky130_fd_sc_hd__o211a_2
XANTENNA__18457__S _18928_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15461__B1 _15424_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19536_ _19784_/CLK _19536_/D vssd1 vssd1 vccd1 vccd1 _19536_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_207_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16748_ _16758_/A _19918_/Q vssd1 vssd1 vccd1 vccd1 _16748_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__19568__CLK _19706_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19467_ _19834_/CLK _19467_/D vssd1 vssd1 vccd1 vccd1 _19467_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16679_ _21167_/Q _11454_/X _21167_/Q _11454_/X vssd1 vssd1 vccd1 vccd1 _16679_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_61_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18950__A1 _21086_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13190__A _13329_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18418_ _18417_/X _16808_/Y _18875_/S vssd1 vssd1 vccd1 vccd1 _18418_/X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_119_HCLK_A clkbuf_opt_3_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19398_ _19812_/CLK _19398_/D vssd1 vssd1 vccd1 vccd1 _19398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18349_ _18348_/X _10133_/Y _18885_/S vssd1 vssd1 vccd1 vccd1 _18349_/X sky130_fd_sc_hd__mux2_1
XANTENNA__18192__S _18884_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21360_ _21367_/CLK _21360_/D repeater254/X vssd1 vssd1 vccd1 vccd1 _21360_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_147_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20311_ _20316_/CLK _20311_/D repeater197/X vssd1 vssd1 vccd1 vccd1 _20311_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_238_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput60 HWDATA[2] vssd1 vssd1 vccd1 vccd1 input60/X sky130_fd_sc_hd__clkbuf_4
XFILLER_116_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21291_ _21357_/CLK _21291_/D repeater199/X vssd1 vssd1 vccd1 vccd1 _21291_/Q sky130_fd_sc_hd__dfrtp_4
Xinput71 MSI_S2 vssd1 vssd1 vccd1 vccd1 input71/X sky130_fd_sc_hd__buf_2
XANTENNA__16006__A _16332_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20242_ _21452_/CLK _20242_/D repeater247/X vssd1 vssd1 vccd1 vccd1 _20242_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_116_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20173_ _20241_/CLK _20173_/D repeater248/X vssd1 vssd1 vccd1 vccd1 _20173_/Q sky130_fd_sc_hd__dfrtp_1
X_09984_ _20020_/Q _10013_/A vssd1 vssd1 vccd1 vccd1 _09985_/A sky130_fd_sc_hd__nand2_1
XFILLER_107_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18218__A0 _12566_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_1_0_HCLK clkbuf_3_1_0_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_3_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10989__A _21017_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18367__S _18775_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18941__A1 _20900_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10690_ _10690_/A vssd1 vssd1 vccd1 vccd1 _10690_/Y sky130_fd_sc_hd__inv_2
XFILLER_197_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20749__RESET_B repeater207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12360_ _20969_/Q _12358_/Y _12359_/X _12323_/B vssd1 vssd1 vccd1 vccd1 _20969_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_120_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11311_ _11311_/A _11311_/B _11306_/B vssd1 vssd1 vccd1 vccd1 _16568_/B sky130_fd_sc_hd__nor3b_4
XFILLER_165_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13518__B1 _13452_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20509_ _20947_/CLK _20509_/D repeater266/X vssd1 vssd1 vccd1 vccd1 _20509_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_148_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12291_ _20526_/Q vssd1 vssd1 vccd1 vccd1 _12291_/Y sky130_fd_sc_hd__inv_2
XFILLER_180_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18830__S _18926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14030_ _14030_/A vssd1 vssd1 vccd1 vccd1 _14031_/A sky130_fd_sc_hd__clkbuf_2
X_11242_ _11241_/A _19911_/Q _11241_/Y _11233_/C vssd1 vssd1 vccd1 vccd1 _11243_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_180_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20331__RESET_B repeater190/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11173_ _11176_/A _11173_/B vssd1 vssd1 vccd1 vccd1 _11173_/X sky130_fd_sc_hd__or2_1
XANTENNA_input40_A HWDATA[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10124_ _10154_/A _20790_/Q _10202_/A _20778_/Q vssd1 vssd1 vccd1 vccd1 _10124_/X
+ sky130_fd_sc_hd__a22o_1
X_15981_ _19544_/Q _15978_/X _15947_/X _15979_/X vssd1 vssd1 vccd1 vccd1 _19544_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17720_ _21133_/Q vssd1 vssd1 vccd1 vccd1 _17720_/Y sky130_fd_sc_hd__inv_2
X_14932_ _14929_/Y _20093_/Q _14930_/Y _20088_/Q _14931_/X vssd1 vssd1 vccd1 vccd1
+ _14933_/D sky130_fd_sc_hd__o221a_1
X_10055_ _21390_/Q vssd1 vssd1 vccd1 vccd1 _10056_/A sky130_fd_sc_hd__inv_2
XFILLER_248_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17651_ _20249_/Q vssd1 vssd1 vccd1 vccd1 _17651_/Y sky130_fd_sc_hd__inv_2
XFILLER_236_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14863_ _15005_/A _15004_/A _14863_/C _15006_/A vssd1 vssd1 vccd1 vccd1 _14864_/D
+ sky130_fd_sc_hd__or4_4
XANTENNA_output127_A _17090_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15443__B1 _15424_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_224_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16602_ _16602_/A _16603_/C vssd1 vssd1 vccd1 vccd1 _16602_/Y sky130_fd_sc_hd__nand2_1
X_13814_ _20188_/Q vssd1 vssd1 vccd1 vccd1 _14577_/A sky130_fd_sc_hd__inv_2
X_17582_ _18750_/X _17823_/A _18754_/X _17820_/A vssd1 vssd1 vccd1 vccd1 _17582_/Y
+ sky130_fd_sc_hd__a22oi_4
XFILLER_223_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14794_ _14794_/A vssd1 vssd1 vccd1 vccd1 _14807_/B sky130_fd_sc_hd__inv_2
XFILLER_44_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19321_ _19626_/CLK _19321_/D vssd1 vssd1 vccd1 vccd1 _19321_/Q sky130_fd_sc_hd__dfxtp_1
X_16533_ _16602_/A vssd1 vssd1 vccd1 vccd1 _16556_/A sky130_fd_sc_hd__buf_1
X_13745_ _20195_/Q vssd1 vssd1 vccd1 vccd1 _14584_/A sky130_fd_sc_hd__inv_2
XFILLER_232_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10957_ _21034_/Q vssd1 vssd1 vccd1 vccd1 _11811_/A sky130_fd_sc_hd__inv_2
XANTENNA__17735__A2 _17856_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_repeater277_A repeater278/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19280__S1 _20122_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18932__A1 _21144_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19252_ _17330_/Y _17331_/Y _17332_/Y _17333_/Y _19275_/S0 _21004_/Q vssd1 vssd1
+ vccd1 vccd1 _19252_/X sky130_fd_sc_hd__mux4_2
XFILLER_232_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14549__A2 _20130_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16464_ _19300_/Q _16459_/X _16342_/X _16460_/X vssd1 vssd1 vccd1 vccd1 _19300_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_189_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13676_ _20354_/Q _13673_/X _13475_/X _13674_/X vssd1 vssd1 vccd1 vccd1 _20354_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_189_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10888_ _10888_/A vssd1 vssd1 vccd1 vccd1 _10888_/X sky130_fd_sc_hd__buf_1
X_18203_ _18202_/X _10106_/Y _18644_/S vssd1 vssd1 vccd1 vccd1 _18203_/X sky130_fd_sc_hd__mux2_1
X_15415_ _15423_/A vssd1 vssd1 vccd1 vccd1 _15415_/X sky130_fd_sc_hd__buf_1
XPHY_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12627_ input4/X _12625_/X _20855_/Q _12626_/X vssd1 vssd1 vccd1 vccd1 _20855_/D
+ sky130_fd_sc_hd__o22a_1
X_19183_ _19546_/Q _19538_/Q _19530_/Q _19514_/Q _19280_/S0 _20122_/Q vssd1 vssd1
+ vccd1 vccd1 _19183_/X sky130_fd_sc_hd__mux4_2
XPHY_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16395_ _19340_/Q _16392_/X _16231_/X _16394_/X vssd1 vssd1 vccd1 vccd1 _19340_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18134_ _18848_/A0 _18060_/Y _18666_/S vssd1 vssd1 vccd1 vccd1 _18134_/X sky130_fd_sc_hd__mux2_1
XFILLER_200_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15346_ _15424_/A vssd1 vssd1 vccd1 vccd1 _15346_/X sky130_fd_sc_hd__clkbuf_2
X_12558_ _20893_/Q _12553_/X _11743_/X _12554_/X vssd1 vssd1 vccd1 vccd1 _20893_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20419__RESET_B repeater187/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11509_ _16338_/A vssd1 vssd1 vccd1 vccd1 _11509_/Y sky130_fd_sc_hd__inv_2
X_18065_ _18065_/A vssd1 vssd1 vccd1 vccd1 _18065_/X sky130_fd_sc_hd__buf_1
X_15277_ _20495_/Q vssd1 vssd1 vccd1 vccd1 _15277_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18740__S _18926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12489_ _20922_/Q _12492_/A _12486_/A _12480_/X vssd1 vssd1 vccd1 vccd1 _20922_/D
+ sky130_fd_sc_hd__o211a_1
X_17016_ _11045_/B _17015_/X _16984_/X vssd1 vssd1 vccd1 vccd1 _17016_/X sky130_fd_sc_hd__o21a_1
XFILLER_144_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14228_ _14228_/A vssd1 vssd1 vccd1 vccd1 _14228_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20072__RESET_B repeater276/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14159_ _20551_/Q vssd1 vssd1 vccd1 vccd1 _14159_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20001__RESET_B repeater225/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18967_ _11341_/B _11375_/B _21184_/Q vssd1 vssd1 vccd1 vccd1 _18967_/X sky130_fd_sc_hd__mux2_1
XFILLER_112_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21278__RESET_B repeater207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17918_ _18448_/X _17214_/X _18431_/X _17203_/X _17917_/X vssd1 vssd1 vccd1 vccd1
+ _17918_/X sky130_fd_sc_hd__o221a_2
XFILLER_224_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18898_ _18897_/X _14566_/A _18898_/S vssd1 vssd1 vccd1 vccd1 _18898_/X sky130_fd_sc_hd__mux2_2
XFILLER_67_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19390__CLK _19813_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18620__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17849_ _20644_/Q vssd1 vssd1 vccd1 vccd1 _17849_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18187__S _18891_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20860_ _21444_/CLK _20860_/D repeater243/X vssd1 vssd1 vccd1 vccd1 _20860_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_241_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19519_ _19521_/CLK _19519_/D vssd1 vssd1 vccd1 vccd1 _19519_/Q sky130_fd_sc_hd__dfxtp_1
X_20791_ _21374_/CLK _20791_/D repeater255/X vssd1 vssd1 vccd1 vccd1 _20791_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_240_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19271__S1 _20133_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20842__RESET_B repeater255/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21412_ _21417_/CLK _21412_/D repeater232/X vssd1 vssd1 vccd1 vccd1 _21412_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_136_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21343_ _21481_/CLK _21343_/D repeater205/X vssd1 vssd1 vccd1 vccd1 _21343_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_162_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18650__S _18666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21274_ _21462_/CLK _21274_/D repeater245/X vssd1 vssd1 vccd1 vccd1 _21274_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_118_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_140_HCLK clkbuf_4_3_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _21207_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_190_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20225_ _21484_/CLK _20225_/D repeater202/X vssd1 vssd1 vccd1 vccd1 _20225_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__13920__B1 _13919_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20156_ _20159_/CLK _20156_/D repeater189/X vssd1 vssd1 vccd1 vccd1 _20156_/Q sky130_fd_sc_hd__dfrtp_1
X_09967_ _09969_/A vssd1 vssd1 vccd1 vccd1 _09975_/A sky130_fd_sc_hd__buf_1
XANTENNA__17790__A _20900_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20087_ _20496_/CLK _20087_/D repeater273/X vssd1 vssd1 vccd1 vccd1 _20087_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09898_ _20006_/Q vssd1 vssd1 vccd1 vccd1 _09898_/X sky130_fd_sc_hd__buf_1
XANTENNA__18611__A0 _17281_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11860_ _21028_/Q _11860_/B vssd1 vssd1 vccd1 vccd1 _11860_/Y sky130_fd_sc_hd__nor2_1
XPHY_4634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10811_ _10811_/A vssd1 vssd1 vccd1 vccd1 _10811_/Y sky130_fd_sc_hd__inv_2
X_11791_ _11794_/A vssd1 vssd1 vccd1 vccd1 _12637_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_214_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20989_ _21191_/CLK _20989_/D repeater222/X vssd1 vssd1 vccd1 vccd1 _20989_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18825__S _18926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19262__S1 _21004_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13530_ _13530_/A _13530_/B vssd1 vssd1 vccd1 vccd1 _13530_/Y sky130_fd_sc_hd__nor2_1
XPHY_3977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10742_ _19931_/Q _19930_/Q _16794_/A vssd1 vssd1 vccd1 vccd1 _16801_/A sky130_fd_sc_hd__or3_4
XFILLER_213_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10673_ _21337_/Q _10672_/Y _10534_/B _10672_/A _10642_/X vssd1 vssd1 vccd1 vccd1
+ _21337_/D sky130_fd_sc_hd__o221a_1
X_13461_ _13483_/A vssd1 vssd1 vccd1 vccd1 _13461_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_40_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_102_HCLK_A clkbuf_4_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15200_ _15068_/B _15202_/A _15068_/A vssd1 vssd1 vccd1 vccd1 _15201_/C sky130_fd_sc_hd__o21a_1
X_12412_ _20949_/Q _12417_/B _12298_/Y _12409_/A _12411_/X vssd1 vssd1 vccd1 vccd1
+ _20949_/D sky130_fd_sc_hd__o221a_1
XFILLER_173_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_165_HCLK_A clkbuf_opt_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16180_ _16187_/A vssd1 vssd1 vccd1 vccd1 _16180_/X sky130_fd_sc_hd__buf_1
X_13392_ _13419_/A vssd1 vssd1 vccd1 vccd1 _13411_/A sky130_fd_sc_hd__buf_1
XANTENNA__20512__RESET_B repeater267/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15131_ _15127_/Y _20054_/Q _20437_/Q _15128_/X _15130_/X vssd1 vssd1 vccd1 vccd1
+ _15131_/X sky130_fd_sc_hd__a221o_1
XFILLER_166_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12343_ _12373_/A vssd1 vssd1 vccd1 vccd1 _12359_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_126_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18560__S _18896_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15062_ _15062_/A _15211_/A vssd1 vssd1 vccd1 vccd1 _15063_/B sky130_fd_sc_hd__or2_2
X_12274_ _20512_/Q vssd1 vssd1 vccd1 vccd1 _12274_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11517__A2 _11497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11225_ _11225_/A vssd1 vssd1 vccd1 vccd1 _11225_/X sky130_fd_sc_hd__buf_1
X_14013_ _14013_/A _14013_/B vssd1 vssd1 vccd1 vccd1 _14023_/A sky130_fd_sc_hd__or2_1
XFILLER_135_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19870_ _21167_/CLK _19870_/D repeater225/X vssd1 vssd1 vccd1 vccd1 _19870_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_150_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18821_ _18820_/X _12195_/Y _18909_/S vssd1 vssd1 vccd1 vccd1 _18821_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11156_ _20430_/Q vssd1 vssd1 vccd1 vccd1 _13180_/A sky130_fd_sc_hd__inv_2
XFILLER_191_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10107_ _10205_/A _20781_/Q _10049_/A _20781_/Q vssd1 vssd1 vccd1 vccd1 _10107_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_68_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18752_ _18751_/X _20569_/Q _18907_/S vssd1 vssd1 vccd1 vccd1 _18752_/X sky130_fd_sc_hd__mux2_1
X_11087_ _11081_/B _11079_/X _11086_/Y _11082_/X _11059_/A vssd1 vssd1 vccd1 vccd1
+ _11088_/A sky130_fd_sc_hd__o32a_1
X_15964_ _19552_/Q _15961_/X _15947_/X _15962_/X vssd1 vssd1 vccd1 vccd1 _19552_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__21371__RESET_B repeater255/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17703_ _18705_/X _17703_/B vssd1 vssd1 vccd1 vccd1 _17703_/X sky130_fd_sc_hd__and2_1
XANTENNA__17405__A1 _17060_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14915_ _20580_/Q vssd1 vssd1 vccd1 vccd1 _14915_/Y sky130_fd_sc_hd__inv_2
X_10038_ _21378_/Q vssd1 vssd1 vccd1 vccd1 _10041_/B sky130_fd_sc_hd__inv_2
XANTENNA__11237__B _19910_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18683_ _18845_/A0 _10320_/Y _18884_/S vssd1 vssd1 vccd1 vccd1 _18683_/X sky130_fd_sc_hd__mux2_1
X_15895_ _19586_/Q _15886_/X _15785_/X _15889_/X vssd1 vssd1 vccd1 vccd1 _19586_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11150__B1 _21004_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17634_ _17777_/A _20114_/Q vssd1 vssd1 vccd1 vccd1 _17634_/Y sky130_fd_sc_hd__nand2_1
X_14846_ _20089_/Q vssd1 vssd1 vccd1 vccd1 _14960_/C sky130_fd_sc_hd__inv_2
XFILLER_223_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_21_HCLK clkbuf_4_3_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _21223_/CLK sky130_fd_sc_hd__clkbuf_16
X_17565_ _21190_/Q vssd1 vssd1 vccd1 vccd1 _17565_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14777_ _14775_/A _14315_/A _15967_/B vssd1 vssd1 vccd1 vccd1 _14777_/X sky130_fd_sc_hd__o21a_1
X_11989_ _19909_/Q vssd1 vssd1 vccd1 vccd1 _12008_/A sky130_fd_sc_hd__inv_2
XANTENNA__18735__S _18930_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19253__S1 _21004_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19304_ _20172_/CLK _19304_/D vssd1 vssd1 vccd1 vccd1 _19304_/Q sky130_fd_sc_hd__dfxtp_1
X_16516_ _16516_/A vssd1 vssd1 vccd1 vccd1 _16632_/B sky130_fd_sc_hd__buf_1
XFILLER_44_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13728_ _15766_/A _15769_/A _13734_/S vssd1 vssd1 vccd1 vccd1 _20327_/D sky130_fd_sc_hd__mux2_1
X_17496_ _19714_/Q vssd1 vssd1 vccd1 vccd1 _17496_/Y sky130_fd_sc_hd__inv_2
XFILLER_232_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19235_ _17496_/Y _17497_/Y _17498_/Y _17499_/Y _19275_/S0 _21004_/Q vssd1 vssd1
+ vccd1 vccd1 _19235_/X sky130_fd_sc_hd__mux4_1
X_16447_ _19850_/D vssd1 vssd1 vccd1 vccd1 _17054_/B sky130_fd_sc_hd__buf_1
XFILLER_176_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13659_ _13679_/A vssd1 vssd1 vccd1 vccd1 _13659_/X sky130_fd_sc_hd__buf_1
XFILLER_31_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19166_ _19162_/X _19163_/X _19164_/X _19165_/X _20123_/Q _20124_/Q vssd1 vssd1 vccd1
+ vccd1 _19166_/X sky130_fd_sc_hd__mux4_2
XANTENNA__09658__A input39/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16378_ _16385_/A vssd1 vssd1 vccd1 vccd1 _16378_/X sky130_fd_sc_hd__buf_1
Xclkbuf_leaf_163_HCLK clkbuf_opt_0_HCLK/A vssd1 vssd1 vccd1 vccd1 _21273_/CLK sky130_fd_sc_hd__clkbuf_16
X_18117_ vssd1 vssd1 vccd1 vccd1 _18117_/HI _18117_/LO sky130_fd_sc_hd__conb_1
XANTENNA__10413__C1 _10381_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17875__A _20344_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15329_ _15329_/A vssd1 vssd1 vccd1 vccd1 _15329_/X sky130_fd_sc_hd__buf_1
X_19097_ _16673_/X _21081_/Q _19870_/D vssd1 vssd1 vccd1 vccd1 _19097_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18470__S _18835_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_24_HCLK_A clkbuf_4_9_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18048_ _18048_/A vssd1 vssd1 vccd1 vccd1 _18048_/X sky130_fd_sc_hd__buf_1
XANTENNA__19756__CLK _19813_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_87_HCLK_A clkbuf_4_12_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21459__RESET_B repeater245/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20010_ _21438_/CLK _20010_/D repeater238/X vssd1 vssd1 vccd1 vccd1 _20010_/Q sky130_fd_sc_hd__dfrtp_1
X_09821_ _15869_/A vssd1 vssd1 vccd1 vccd1 _09821_/X sky130_fd_sc_hd__buf_1
XFILLER_99_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19999_ _21167_/CLK _19999_/D repeater225/X vssd1 vssd1 vccd1 vccd1 _19999_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09752_ _20147_/Q vssd1 vssd1 vccd1 vccd1 _09752_/Y sky130_fd_sc_hd__inv_2
XFILLER_228_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09683_ _21468_/Q _09673_/X _09682_/X _09678_/X vssd1 vssd1 vccd1 vccd1 _21468_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__15407__B1 _15346_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20912_ _20915_/CLK _20912_/D repeater217/X vssd1 vssd1 vccd1 vccd1 _20912_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__11692__A1 _21082_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20843_ _21444_/CLK _20843_/D repeater246/X vssd1 vssd1 vccd1 vccd1 _20843_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__09637__A1 _21480_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18645__S _18886_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19244__S1 _21004_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20774_ _21379_/CLK _20774_/D repeater213/X vssd1 vssd1 vccd1 vccd1 _20774_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10507__A _20693_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18380__S _18680_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21326_ _21341_/CLK _21326_/D repeater201/X vssd1 vssd1 vccd1 vccd1 _21326_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_163_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15894__B1 _15893_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21257_ _21390_/CLK _21257_/D repeater239/X vssd1 vssd1 vccd1 vccd1 _21257_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12722__A _17177_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11010_ _15505_/A _15505_/B _15374_/B vssd1 vssd1 vccd1 vccd1 _11010_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_132_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19180__S0 _19280_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20208_ _20241_/CLK _20208_/D repeater248/X vssd1 vssd1 vccd1 vccd1 _20208_/Q sky130_fd_sc_hd__dfrtp_2
X_21188_ _21191_/CLK _21188_/D repeater224/X vssd1 vssd1 vccd1 vccd1 _21188_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_49_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20139_ _21218_/CLK _20139_/D repeater250/X vssd1 vssd1 vccd1 vccd1 _20139_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_237_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_44_HCLK clkbuf_4_11_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _21185_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_58_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12961_ _12961_/A vssd1 vssd1 vccd1 vccd1 _12961_/X sky130_fd_sc_hd__buf_1
XANTENNA__17399__B1 _18802_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13553__A input56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14700_ _20160_/Q _14696_/X _18243_/X _14688_/X vssd1 vssd1 vccd1 vccd1 _20160_/D
+ sky130_fd_sc_hd__a22o_1
X_11912_ _11003_/X _11906_/Y _11910_/X vssd1 vssd1 vccd1 vccd1 _21014_/D sky130_fd_sc_hd__o21a_1
XANTENNA__11683__A1 _21087_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15680_ _19682_/Q _15674_/X _15582_/X _15676_/X vssd1 vssd1 vccd1 vccd1 _19682_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12880__B1 _12879_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12892_ _13106_/B vssd1 vssd1 vccd1 vccd1 _17087_/A sky130_fd_sc_hd__clkbuf_4
XPHY_4431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14631_ _20189_/Q _14630_/Y _14624_/X _14579_/B vssd1 vssd1 vccd1 vccd1 _20189_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_54_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11843_ _11838_/B _11827_/X _11842_/Y _11834_/X _11810_/A vssd1 vssd1 vccd1 vccd1
+ _11844_/A sky130_fd_sc_hd__o32a_1
XPHY_4464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18555__S _18910_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20764__RESET_B repeater211/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19235__S1 _21004_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_221_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17350_ _19480_/Q vssd1 vssd1 vccd1 vccd1 _17350_/Y sky130_fd_sc_hd__inv_2
XFILLER_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14562_ _15799_/A _15833_/B _14541_/A _15816_/A _14561_/Y vssd1 vssd1 vccd1 vccd1
+ _14562_/X sky130_fd_sc_hd__o32a_1
XPHY_3763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11774_ _19089_/X _11770_/X _21045_/Q _11771_/X vssd1 vssd1 vccd1 vccd1 _21045_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_214_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16301_ _19389_/Q _16298_/X _16277_/X _16300_/X vssd1 vssd1 vccd1 vccd1 _19389_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13513_ _20437_/Q _13505_/X _13442_/X _13507_/X vssd1 vssd1 vccd1 vccd1 _20437_/D
+ sky130_fd_sc_hd__a22o_1
X_10725_ _10725_/A _10725_/B _10729_/C vssd1 vssd1 vccd1 vccd1 _21313_/D sky130_fd_sc_hd__nor3_1
XFILLER_158_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17281_ _18901_/S _18899_/S _18910_/S _17193_/B vssd1 vssd1 vccd1 vccd1 _17281_/X
+ sky130_fd_sc_hd__or4b_4
X_14493_ _14493_/A vssd1 vssd1 vccd1 vccd1 _14493_/Y sky130_fd_sc_hd__inv_2
XFILLER_201_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19020_ _16911_/X _20403_/Q _19026_/S vssd1 vssd1 vccd1 vccd1 _19956_/D sky130_fd_sc_hd__mux2_1
X_16232_ _16240_/A vssd1 vssd1 vccd1 vccd1 _16241_/A sky130_fd_sc_hd__inv_2
X_13444_ _13444_/A vssd1 vssd1 vccd1 vccd1 _13444_/X sky130_fd_sc_hd__buf_1
XANTENNA__19779__CLK _21009_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10656_ _10656_/A _10690_/A vssd1 vssd1 vccd1 vccd1 _10657_/B sky130_fd_sc_hd__or2_2
X_16163_ _16163_/A vssd1 vssd1 vccd1 vccd1 _16163_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_127_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10587_ _10705_/A _20745_/Q _21317_/Q _10583_/Y _10586_/X vssd1 vssd1 vccd1 vccd1
+ _10591_/C sky130_fd_sc_hd__o221a_1
XANTENNA__18290__S _18928_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13375_ _20503_/Q _13371_/X _13245_/X _13372_/X vssd1 vssd1 vccd1 vccd1 _20503_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_6_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15114_ _20451_/Q _15076_/A _15111_/Y _20050_/Q _15113_/X vssd1 vssd1 vccd1 vccd1
+ _15126_/A sky130_fd_sc_hd__a221o_1
XFILLER_126_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12326_ _12326_/A _12352_/A vssd1 vssd1 vccd1 vccd1 _12327_/B sky130_fd_sc_hd__or2_2
X_16094_ _16101_/A vssd1 vssd1 vccd1 vccd1 _16094_/X sky130_fd_sc_hd__buf_1
XFILLER_108_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19922_ _21141_/CLK _19922_/D repeater212/X vssd1 vssd1 vccd1 vccd1 _19922_/Q sky130_fd_sc_hd__dfrtp_1
X_15045_ _20057_/Q vssd1 vssd1 vccd1 vccd1 _15071_/A sky130_fd_sc_hd__inv_2
X_12257_ _20938_/Q vssd1 vssd1 vccd1 vccd1 _12258_/A sky130_fd_sc_hd__inv_2
XFILLER_123_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19171__S0 _20123_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11208_ _11226_/A vssd1 vssd1 vccd1 vccd1 _11208_/X sky130_fd_sc_hd__buf_1
X_19853_ _21429_/CLK _19853_/D repeater229/X vssd1 vssd1 vccd1 vccd1 _19853_/Q sky130_fd_sc_hd__dfrtp_1
X_12188_ _12064_/Y _20363_/Q _20973_/Q _12187_/Y vssd1 vssd1 vccd1 vccd1 _12188_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_150_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18804_ _18803_/X _16755_/Y _18880_/S vssd1 vssd1 vccd1 vccd1 _18804_/X sky130_fd_sc_hd__mux2_1
XANTENNA__15943__A _15943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19947__RESET_B repeater251/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15101__A2 _20062_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11139_ _11176_/B _11136_/X _15609_/B _21003_/Q _11138_/Y vssd1 vssd1 vccd1 vccd1
+ _11151_/B sky130_fd_sc_hd__a221o_1
XFILLER_205_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16996_ _19976_/Q vssd1 vssd1 vccd1 vccd1 _16999_/A sky130_fd_sc_hd__inv_2
X_19784_ _19784_/CLK _19784_/D vssd1 vssd1 vccd1 vccd1 _19784_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15947_ _16012_/A vssd1 vssd1 vccd1 vccd1 _15947_/X sky130_fd_sc_hd__clkbuf_2
X_18735_ _18734_/X _19221_/X _18930_/S vssd1 vssd1 vccd1 vccd1 _18735_/X sky130_fd_sc_hd__mux2_2
XFILLER_110_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11674__A1 _16654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18666_ _18665_/X _18069_/Y _18666_/S vssd1 vssd1 vccd1 vccd1 _18666_/X sky130_fd_sc_hd__mux2_1
XFILLER_224_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12871__B1 _12550_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15878_ _19593_/Q _15875_/X _15876_/X _15877_/X vssd1 vssd1 vccd1 vccd1 _19593_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_64_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17617_ _19595_/Q vssd1 vssd1 vccd1 vccd1 _17617_/Y sky130_fd_sc_hd__inv_2
X_14829_ _20103_/Q vssd1 vssd1 vccd1 vccd1 _14881_/B sky130_fd_sc_hd__inv_2
X_18597_ _18848_/A0 _10292_/Y _18884_/S vssd1 vssd1 vccd1 vccd1 _18597_/X sky130_fd_sc_hd__mux2_1
XANTENNA__19226__S1 _21006_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18465__S _18617_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17548_ _17548_/A vssd1 vssd1 vccd1 vccd1 _17548_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__20434__RESET_B repeater278/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17479_ _18782_/X _17211_/A _18785_/X _17319_/X _17478_/X vssd1 vssd1 vccd1 vccd1
+ _17479_/X sky130_fd_sc_hd__o221a_2
XANTENNA__11711__A _17553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19218_ _17615_/Y _17616_/Y _17617_/Y _17618_/Y _20130_/Q _20131_/Q vssd1 vssd1 vccd1
+ vccd1 _19218_/X sky130_fd_sc_hd__mux4_2
X_20490_ _20944_/CLK _20490_/D repeater274/X vssd1 vssd1 vccd1 vccd1 _20490_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_146_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19149_ _19690_/Q _19378_/Q _19674_/Q _19666_/Q _19285_/S0 _21017_/Q vssd1 vssd1
+ vccd1 vccd1 _19149_/X sky130_fd_sc_hd__mux4_2
XFILLER_118_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21111_ _21417_/CLK _21111_/D repeater234/X vssd1 vssd1 vccd1 vccd1 _21111_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_117_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_246_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21293__RESET_B repeater211/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16014__A _16340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19162__S0 _19280_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21042_ _21183_/CLK _21042_/D repeater219/X vssd1 vssd1 vccd1 vccd1 _21042_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA__18814__A0 _18848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_67_HCLK clkbuf_4_11_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20256_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_99_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21222__RESET_B repeater235/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15628__B1 _15544_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09804_ _09804_/A _09806_/A _09804_/C vssd1 vssd1 vccd1 vccd1 _09804_/X sky130_fd_sc_hd__or3_1
XFILLER_140_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_247_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09735_ _11054_/A _09734_/Y _21229_/Q _20149_/Q vssd1 vssd1 vccd1 vccd1 _09742_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_74_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12862__B1 _12860_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09666_ _13313_/A vssd1 vssd1 vccd1 vccd1 _09666_/X sky130_fd_sc_hd__buf_6
XFILLER_243_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18375__S _18669_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19217__S1 _20131_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09597_ _13047_/B vssd1 vssd1 vccd1 vccd1 _10859_/B sky130_fd_sc_hd__buf_2
XPHY_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20826_ _20841_/CLK _20826_/D repeater251/X vssd1 vssd1 vccd1 vccd1 _20826_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20175__RESET_B repeater249/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20757_ _21477_/CLK _20757_/D repeater201/X vssd1 vssd1 vccd1 vccd1 _20757_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_24_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20104__RESET_B repeater259/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10510_ _21283_/Q vssd1 vssd1 vccd1 vccd1 _10760_/A sky130_fd_sc_hd__inv_2
XPHY_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11490_ _15847_/B vssd1 vssd1 vccd1 vccd1 _17549_/A sky130_fd_sc_hd__clkbuf_2
XPHY_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20688_ _21486_/CLK _20688_/D repeater199/X vssd1 vssd1 vccd1 vccd1 _20688_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10441_ _20671_/Q vssd1 vssd1 vccd1 vccd1 _10441_/Y sky130_fd_sc_hd__inv_2
XFILLER_136_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13160_ _20606_/Q _13158_/X _12950_/X _13159_/X vssd1 vssd1 vccd1 vccd1 _20606_/D
+ sky130_fd_sc_hd__a22o_1
X_10372_ _10372_/A vssd1 vssd1 vccd1 vccd1 _10372_/Y sky130_fd_sc_hd__inv_2
XFILLER_200_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12111_ _12105_/X _20384_/Q _12330_/A _20391_/Q _12110_/X vssd1 vssd1 vccd1 vccd1
+ _12145_/B sky130_fd_sc_hd__o221a_1
X_21309_ _21406_/CLK _21309_/D repeater211/X vssd1 vssd1 vccd1 vccd1 _21309_/Q sky130_fd_sc_hd__dfrtp_1
X_13091_ _20642_/Q _13086_/X _13032_/X _13087_/X vssd1 vssd1 vccd1 vccd1 _20642_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_70_HCLK_A clkbuf_opt_7_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12042_ _20394_/Q vssd1 vssd1 vccd1 vccd1 _12042_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19153__S0 _19285_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18805__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16850_ _19942_/Q vssd1 vssd1 vccd1 vccd1 _16850_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_238_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15801_ _15807_/A vssd1 vssd1 vccd1 vccd1 _15808_/A sky130_fd_sc_hd__inv_2
XFILLER_65_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16781_ _19926_/Q vssd1 vssd1 vccd1 vccd1 _16781_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13993_ _13993_/A vssd1 vssd1 vccd1 vccd1 _13993_/Y sky130_fd_sc_hd__inv_2
X_18520_ _18519_/X _14087_/A _18850_/S vssd1 vssd1 vccd1 vccd1 _18520_/X sky130_fd_sc_hd__mux2_1
XFILLER_207_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15732_ input65/X vssd1 vssd1 vccd1 vccd1 _16237_/A sky130_fd_sc_hd__buf_2
X_12944_ _20714_/Q _12942_/X _12860_/X _12943_/X vssd1 vssd1 vccd1 vccd1 _20714_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16044__B1 _16009_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18451_ _18450_/X _10271_/A _18841_/S vssd1 vssd1 vccd1 vccd1 _18451_/X sky130_fd_sc_hd__mux2_1
X_15663_ _15663_/A vssd1 vssd1 vccd1 vccd1 _15663_/X sky130_fd_sc_hd__buf_1
XPHY_4250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18285__S _18896_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12875_ _13166_/A vssd1 vssd1 vccd1 vccd1 _12875_/X sky130_fd_sc_hd__buf_2
XANTENNA__19208__S1 _20131_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17402_ _18822_/X _17401_/X _18829_/X _17320_/X vssd1 vssd1 vccd1 vccd1 _17402_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_4272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14614_ _20199_/Q _14613_/Y _14610_/X _14589_/B vssd1 vssd1 vccd1 vccd1 _20199_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_45_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18382_ _18381_/X _12172_/Y _18909_/S vssd1 vssd1 vccd1 vccd1 _18382_/X sky130_fd_sc_hd__mux2_1
X_11826_ _11822_/A _11816_/Y _11825_/X _11817_/X _21037_/Q vssd1 vssd1 vccd1 vccd1
+ _21037_/D sky130_fd_sc_hd__a32o_1
XPHY_4294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15594_ _15594_/A _16616_/B vssd1 vssd1 vccd1 vccd1 _16261_/C sky130_fd_sc_hd__or2_2
XPHY_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17333_ _19472_/Q vssd1 vssd1 vccd1 vccd1 _17333_/Y sky130_fd_sc_hd__inv_2
XFILLER_230_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14545_ _20134_/Q vssd1 vssd1 vccd1 vccd1 _15798_/B sky130_fd_sc_hd__buf_1
X_11757_ _19873_/Q _19872_/Q vssd1 vssd1 vccd1 vccd1 _11770_/A sky130_fd_sc_hd__or2_1
XPHY_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10708_ _10708_/A _10708_/B vssd1 vssd1 vccd1 vccd1 _10708_/Y sky130_fd_sc_hd__nor2_2
X_17264_ _19575_/Q vssd1 vssd1 vccd1 vccd1 _17264_/Y sky130_fd_sc_hd__inv_2
X_14476_ _14476_/A vssd1 vssd1 vccd1 vccd1 _14476_/Y sky130_fd_sc_hd__inv_2
XPHY_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11688_ _21084_/Q _11679_/X _11560_/X _11682_/X vssd1 vssd1 vccd1 vccd1 _21084_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_197_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19003_ _16985_/X _20420_/Q _19019_/S vssd1 vssd1 vccd1 vccd1 _19973_/D sky130_fd_sc_hd__mux2_1
XFILLER_128_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16215_ _16247_/A _16215_/B _16297_/C vssd1 vssd1 vccd1 vccd1 _16223_/A sky130_fd_sc_hd__or3_4
X_13427_ _20477_/Q _13417_/X _13426_/X _13420_/X vssd1 vssd1 vccd1 vccd1 _20477_/D
+ sky130_fd_sc_hd__a22o_1
X_10639_ _10639_/A _10639_/B _10639_/C _10639_/D vssd1 vssd1 vccd1 vccd1 _10685_/A
+ sky130_fd_sc_hd__and4_1
X_17195_ _17195_/A vssd1 vssd1 vccd1 vccd1 _17472_/A sky130_fd_sc_hd__buf_1
XFILLER_127_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16146_ _19464_/Q _16141_/X _16145_/X _16143_/X vssd1 vssd1 vccd1 vccd1 _19464_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09936__A _20888_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13358_ _13377_/A vssd1 vssd1 vccd1 vccd1 _13358_/X sky130_fd_sc_hd__buf_1
XFILLER_182_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15858__B1 _15788_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12309_ _12309_/A _12383_/A vssd1 vssd1 vccd1 vccd1 _12310_/B sky130_fd_sc_hd__or2_1
XANTENNA__13458__A _13481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16077_ _16077_/A vssd1 vssd1 vccd1 vccd1 _16405_/A sky130_fd_sc_hd__buf_1
X_13289_ _20553_/Q _13286_/X _13287_/X _13288_/X vssd1 vssd1 vccd1 vccd1 _20553_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19144__S0 _19285_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19905_ _20256_/CLK _19905_/D repeater217/X vssd1 vssd1 vccd1 vccd1 _19905_/Q sky130_fd_sc_hd__dfrtp_1
X_15028_ _20073_/Q vssd1 vssd1 vccd1 vccd1 _15029_/A sky130_fd_sc_hd__clkbuf_2
X_19836_ _20172_/CLK _19836_/D vssd1 vssd1 vccd1 vccd1 _19836_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19767_ _19828_/CLK _19767_/D vssd1 vssd1 vccd1 vccd1 _19767_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13097__B1 _12872_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16979_ _16979_/A _16979_/B vssd1 vssd1 vccd1 vccd1 _16980_/A sky130_fd_sc_hd__or2_1
Xinput3 HADDR[11] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_1
XFILLER_237_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18718_ _18717_/X _10759_/A _18880_/S vssd1 vssd1 vccd1 vccd1 _18718_/X sky130_fd_sc_hd__mux2_1
XFILLER_232_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12844__B1 _09633_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_225_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19698_ _21222_/CLK _19698_/D vssd1 vssd1 vccd1 vccd1 _19698_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_225_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18649_ _18648_/X _14945_/Y _18907_/S vssd1 vssd1 vccd1 vccd1 _18649_/X sky130_fd_sc_hd__mux2_2
XANTENNA__18195__S _18896_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_240_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20921__CLK _20930_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20611_ _20657_/CLK _20611_/D repeater198/X vssd1 vssd1 vccd1 vccd1 _20611_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_32_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12072__B2 _20393_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18923__S _18928_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20542_ _20724_/CLK _20542_/D repeater264/X vssd1 vssd1 vccd1 vccd1 _20542_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20473_ _20476_/CLK _20473_/D repeater280/X vssd1 vssd1 vccd1 vccd1 _20473_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21474__RESET_B repeater204/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14752__A _20132_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21403__RESET_B repeater255/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19869__RESET_B repeater216/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19135__S0 _19285_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21025_ _21401_/CLK _21025_/D repeater241/X vssd1 vssd1 vccd1 vccd1 _21025_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_102_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_3_1_0_HCLK_A clkbuf_3_1_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13088__B1 _12860_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09718_ _21225_/Q vssd1 vssd1 vccd1 vccd1 _11112_/A sky130_fd_sc_hd__inv_2
XFILLER_27_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10990_ _21016_/Q vssd1 vssd1 vccd1 vccd1 _10991_/B sky130_fd_sc_hd__inv_2
XFILLER_71_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09649_ _12855_/A vssd1 vssd1 vccd1 vccd1 _09649_/X sky130_fd_sc_hd__buf_4
XFILLER_27_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_215_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17303__A _21137_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_230_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12660_ input58/X vssd1 vssd1 vccd1 vccd1 _12660_/X sky130_fd_sc_hd__clkbuf_4
XPHY_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11611_ _11636_/A _21112_/Q _21111_/Q vssd1 vssd1 vccd1 vccd1 _21112_/D sky130_fd_sc_hd__a21o_1
XPHY_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20809_ _20809_/CLK _20809_/D repeater189/X vssd1 vssd1 vccd1 vccd1 _20809_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13260__A0 _13254_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12591_ _20879_/Q _12588_/X _18231_/X _12589_/X vssd1 vssd1 vccd1 vccd1 _20879_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18833__S _18929_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14330_ _20233_/Q vssd1 vssd1 vccd1 vccd1 _14465_/B sky130_fd_sc_hd__inv_2
XPHY_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11542_ _11542_/A vssd1 vssd1 vccd1 vccd1 _11542_/Y sky130_fd_sc_hd__inv_2
XANTENNA__10613__A2 _10609_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17957__B _17957_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14261_ _16720_/A _14257_/X _14258_/X _14260_/X vssd1 vssd1 vccd1 vccd1 _20251_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11473_ _19098_/X _11468_/X _21160_/Q _11469_/X vssd1 vssd1 vccd1 vccd1 _21160_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_7_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16000_ _16008_/A vssd1 vssd1 vccd1 vccd1 _16000_/X sky130_fd_sc_hd__buf_1
XFILLER_7_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input70_A HWRITE vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13212_ _20586_/Q _13206_/X _13211_/X _13207_/X vssd1 vssd1 vccd1 vccd1 _20586_/D
+ sky130_fd_sc_hd__a22o_1
X_10424_ _21285_/Q vssd1 vssd1 vccd1 vccd1 _10762_/A sky130_fd_sc_hd__inv_2
XFILLER_125_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14192_ _20282_/Q _14190_/Y _14093_/B _14191_/X vssd1 vssd1 vccd1 vccd1 _20282_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_151_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13143_ _20614_/Q _13139_/X _13140_/X _13142_/X vssd1 vssd1 vccd1 vccd1 _20614_/D
+ sky130_fd_sc_hd__a22o_1
X_10355_ _20719_/Q vssd1 vssd1 vccd1 vccd1 _10355_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17951_ _17951_/A vssd1 vssd1 vccd1 vccd1 _17951_/X sky130_fd_sc_hd__buf_1
X_10286_ _10286_/A _10372_/A vssd1 vssd1 vccd1 vccd1 _10287_/B sky130_fd_sc_hd__or2_2
X_13074_ _20653_/Q _13072_/X _12925_/X _13073_/X vssd1 vssd1 vccd1 vccd1 _20653_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_105_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12025_ _19075_/X _12023_/X _20990_/Q _12024_/X vssd1 vssd1 vccd1 vccd1 _20990_/D
+ sky130_fd_sc_hd__a22o_1
X_16902_ _16902_/A _16902_/B vssd1 vssd1 vccd1 vccd1 _16902_/Y sky130_fd_sc_hd__nor2_1
XFILLER_78_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17882_ _18463_/X _17861_/X _18451_/X _17862_/X _17881_/X vssd1 vssd1 vccd1 vccd1
+ _17882_/X sky130_fd_sc_hd__o221a_2
XFILLER_38_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19621_ _21452_/CLK _19621_/D vssd1 vssd1 vccd1 vccd1 _19621_/Q sky130_fd_sc_hd__dfxtp_1
X_16833_ _19938_/Q vssd1 vssd1 vccd1 vccd1 _16834_/A sky130_fd_sc_hd__buf_1
XFILLER_238_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16764_ _19922_/Q vssd1 vssd1 vccd1 vccd1 _16766_/A sky130_fd_sc_hd__inv_2
X_19552_ _19706_/CLK _19552_/D vssd1 vssd1 vccd1 vccd1 _19552_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12826__B1 _12656_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13976_ _13974_/X _20315_/Q _20316_/Q _13976_/D vssd1 vssd1 vccd1 vccd1 _13977_/C
+ sky130_fd_sc_hd__and4b_1
XFILLER_202_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16017__B1 _16016_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20097__RESET_B repeater259/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18503_ _18502_/X _10609_/Y _18775_/S vssd1 vssd1 vccd1 vccd1 _18503_/X sky130_fd_sc_hd__mux2_1
X_15715_ _19666_/Q _15709_/X _15694_/X _15711_/X vssd1 vssd1 vccd1 vccd1 _19666_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_207_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12927_ _20722_/Q _12924_/X _12925_/X _12926_/X vssd1 vssd1 vccd1 vccd1 _20722_/D
+ sky130_fd_sc_hd__a22o_1
X_16695_ _19892_/Q _14232_/B _14233_/B vssd1 vssd1 vccd1 vccd1 _16695_/X sky130_fd_sc_hd__a21bo_1
X_19483_ _19626_/CLK _19483_/D vssd1 vssd1 vccd1 vccd1 _19483_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10301__A1 _21373_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18434_ _17903_/Y _16941_/Y _18680_/S vssd1 vssd1 vccd1 vccd1 _18434_/X sky130_fd_sc_hd__mux2_2
X_15646_ _19698_/Q _15640_/X _15477_/X _15642_/X vssd1 vssd1 vccd1 vccd1 _19698_/D
+ sky130_fd_sc_hd__a22o_1
X_12858_ _20750_/Q _12848_/X _12857_/X _12851_/X vssd1 vssd1 vccd1 vccd1 _20750_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15240__B2 _20062_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18365_ _18364_/X _21301_/Q _18617_/S vssd1 vssd1 vccd1 vccd1 _18365_/X sky130_fd_sc_hd__mux2_2
XFILLER_33_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11809_ _11845_/A _11845_/B vssd1 vssd1 vccd1 vccd1 _11841_/A sky130_fd_sc_hd__or2_1
XFILLER_21_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15577_ _15584_/A vssd1 vssd1 vccd1 vccd1 _15586_/A sky130_fd_sc_hd__inv_2
XANTENNA__13251__B1 _13169_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12789_ _20786_/Q _12784_/X _09649_/X _12786_/X vssd1 vssd1 vccd1 vccd1 _20786_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18743__S _18885_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17316_ _17316_/A vssd1 vssd1 vccd1 vccd1 _17844_/A sky130_fd_sc_hd__buf_1
X_14528_ _14528_/A _21458_/Q vssd1 vssd1 vccd1 vccd1 _14529_/B sky130_fd_sc_hd__nor2_1
XFILLER_202_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18296_ _18848_/A0 _10333_/Y _18884_/S vssd1 vssd1 vccd1 vccd1 _18296_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17247_ _19719_/Q vssd1 vssd1 vccd1 vccd1 _17247_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14459_ _20238_/Q _14467_/A _14458_/X _14382_/B vssd1 vssd1 vccd1 vccd1 _20238_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_175_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17178_ _17178_/A vssd1 vssd1 vccd1 vccd1 _17193_/B sky130_fd_sc_hd__buf_2
X_16129_ _16179_/A _16150_/B _16377_/C vssd1 vssd1 vccd1 vccd1 _16141_/A sky130_fd_sc_hd__or3_4
XANTENNA__13188__A _13188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17296__A2 _17141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19962__RESET_B repeater185/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20867__RESET_B repeater247/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19819_ _19821_/CLK _19819_/D vssd1 vssd1 vccd1 vccd1 _19819_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_217_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13490__B1 _13489_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13949__A1_N _20648_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17220__A2 _17854_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_212_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18653__S _18875_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13242__B1 _13240_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20525_ _20944_/CLK _20525_/D repeater275/X vssd1 vssd1 vccd1 vccd1 _20525_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_20_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20456_ _20476_/CLK _20456_/D repeater279/X vssd1 vssd1 vccd1 vccd1 _20456_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_4_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11556__B1 _10886_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20387_ _20972_/CLK _20387_/D repeater280/X vssd1 vssd1 vccd1 vccd1 _20387_/Q sky130_fd_sc_hd__dfrtp_1
X_10140_ _10183_/A vssd1 vssd1 vccd1 vccd1 _10140_/X sky130_fd_sc_hd__buf_1
XFILLER_133_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10071_ _10071_/A vssd1 vssd1 vccd1 vccd1 _10159_/A sky130_fd_sc_hd__buf_1
XANTENNA__20537__RESET_B repeater267/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21008_ _21009_/CLK _21008_/D repeater235/X vssd1 vssd1 vccd1 vccd1 _21008_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_101_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_236_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18828__S _18929_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13830_ _20600_/Q vssd1 vssd1 vccd1 vccd1 _13830_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12808__B1 _11743_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20190__RESET_B repeater200/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13761_ _13761_/A _13761_/B _13761_/C _13761_/D vssd1 vssd1 vccd1 vccd1 _13837_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_28_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10973_ _20888_/Q _20887_/Q _10973_/C vssd1 vssd1 vccd1 vccd1 _13047_/C sky130_fd_sc_hd__or3_4
X_15500_ _15500_/A vssd1 vssd1 vccd1 vccd1 _15500_/X sky130_fd_sc_hd__buf_1
XFILLER_243_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12712_ _20811_/Q _12707_/X _11743_/X _12708_/X vssd1 vssd1 vccd1 vccd1 _20811_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13561__A _13567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16480_ _16480_/A vssd1 vssd1 vccd1 vccd1 _19126_/S sky130_fd_sc_hd__inv_2
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13692_ _20344_/Q _13686_/X _12857_/A _13688_/X vssd1 vssd1 vccd1 vccd1 _20344_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_15_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20256__SET_B repeater217/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15431_ _15592_/A vssd1 vssd1 vccd1 vccd1 _15431_/X sky130_fd_sc_hd__clkbuf_2
X_12643_ input1/X _12619_/A _20843_/Q _12620_/A vssd1 vssd1 vccd1 vccd1 _20843_/D
+ sky130_fd_sc_hd__o22a_1
XPHY_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18563__S _18835_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18150_ _17281_/X _17992_/Y _18787_/S vssd1 vssd1 vccd1 vccd1 _18150_/X sky130_fd_sc_hd__mux2_1
XPHY_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15362_ _19829_/Q _15359_/X _14258_/X _15361_/X vssd1 vssd1 vccd1 vccd1 _19829_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__21325__RESET_B repeater204/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12574_ _12574_/A vssd1 vssd1 vccd1 vccd1 _12574_/X sky130_fd_sc_hd__buf_1
XPHY_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18172__A0 _18848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17101_ _19518_/Q vssd1 vssd1 vccd1 vccd1 _17101_/Y sky130_fd_sc_hd__inv_2
XPHY_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14313_ _20241_/Q vssd1 vssd1 vccd1 vccd1 _14313_/Y sky130_fd_sc_hd__inv_2
XFILLER_184_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18081_ _18081_/A _18083_/B vssd1 vssd1 vccd1 vccd1 _18081_/Y sky130_fd_sc_hd__nor2_1
XPHY_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11525_ _14256_/B vssd1 vssd1 vccd1 vccd1 _14273_/D sky130_fd_sc_hd__clkbuf_2
X_15293_ _19859_/Q _15293_/B vssd1 vssd1 vccd1 vccd1 _15294_/B sky130_fd_sc_hd__or2_1
XFILLER_157_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14392__A _20026_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17032_ _17032_/A _17035_/B vssd1 vssd1 vccd1 vccd1 _20016_/D sky130_fd_sc_hd__nor2_1
X_14244_ _14246_/A vssd1 vssd1 vccd1 vccd1 _14249_/A sky130_fd_sc_hd__inv_2
XFILLER_7_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11456_ _19850_/Q vssd1 vssd1 vccd1 vccd1 _11457_/C sky130_fd_sc_hd__inv_2
X_10407_ _10346_/X _10406_/A _21353_/Q _10406_/Y _10364_/X vssd1 vssd1 vccd1 vccd1
+ _21353_/D sky130_fd_sc_hd__o221a_1
XANTENNA__18014__D _18014_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14175_ _20290_/Q _14100_/Y _14101_/Y _14100_/A _14174_/X vssd1 vssd1 vccd1 vccd1
+ _20290_/D sky130_fd_sc_hd__o221a_1
X_11387_ _11387_/A _11387_/B _11379_/B vssd1 vssd1 vccd1 vccd1 _11389_/B sky130_fd_sc_hd__nor3b_4
X_13126_ _13132_/A vssd1 vssd1 vccd1 vccd1 _13126_/X sky130_fd_sc_hd__buf_1
X_10338_ _21366_/Q _18006_/A _10281_/A _20725_/Q vssd1 vssd1 vccd1 vccd1 _10338_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_112_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18983_ _21423_/Q _21096_/Q _18983_/S vssd1 vssd1 vccd1 vccd1 _18983_/X sky130_fd_sc_hd__mux2_1
XFILLER_113_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20960__RESET_B repeater186/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17934_ _18507_/X _17203_/X _18536_/X _17947_/A vssd1 vssd1 vccd1 vccd1 _17934_/X
+ sky130_fd_sc_hd__o22a_1
X_13057_ _20664_/Q _13052_/X _12989_/X _13055_/X vssd1 vssd1 vccd1 vccd1 _20664_/D
+ sky130_fd_sc_hd__a22o_1
X_10269_ _10269_/A _10346_/A _10406_/A vssd1 vssd1 vccd1 vccd1 _10402_/A sky130_fd_sc_hd__or3_1
XANTENNA__20278__RESET_B repeater262/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16238__B1 _16237_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12008_ _12008_/A _19908_/D vssd1 vssd1 vccd1 vccd1 _12011_/A sky130_fd_sc_hd__or2_1
X_17865_ _17852_/X _17855_/X _17860_/X _17864_/X vssd1 vssd1 vccd1 vccd1 _17865_/Y
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__18738__S _18929_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15951__A _16016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19604_ _20142_/CLK _19604_/D vssd1 vssd1 vccd1 vccd1 _19604_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_226_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16816_ _16814_/Y _16815_/Y _16803_/X vssd1 vssd1 vccd1 vccd1 _16816_/X sky130_fd_sc_hd__o21a_1
XFILLER_213_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17796_ _17792_/Y _17290_/X _16691_/A _17292_/X _17795_/X vssd1 vssd1 vccd1 vccd1
+ _17796_/X sky130_fd_sc_hd__o221a_1
X_19535_ _21462_/CLK _19535_/D vssd1 vssd1 vccd1 vccd1 _19535_/Q sky130_fd_sc_hd__dfxtp_1
X_16747_ _16835_/A vssd1 vssd1 vccd1 vccd1 _16758_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_19_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13959_ _13958_/Y _20314_/Q _20657_/Q _13974_/C vssd1 vssd1 vccd1 vccd1 _13959_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_222_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_234_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16678_ _21166_/Q _11454_/B _11454_/X vssd1 vssd1 vccd1 vccd1 _16678_/X sky130_fd_sc_hd__a21bo_1
X_19466_ _20136_/CLK _19466_/D vssd1 vssd1 vccd1 vccd1 _19466_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18417_ _18848_/A0 _17912_/Y _18874_/S vssd1 vssd1 vccd1 vccd1 _18417_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13190__B _13456_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15629_ _19708_/Q _15625_/X _15548_/X _15627_/X vssd1 vssd1 vccd1 vccd1 _19708_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18473__S _18897_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16782__A _16835_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19397_ _21001_/CLK _19397_/D vssd1 vssd1 vccd1 vccd1 _19397_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09979__B1 _09688_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18163__A0 _18848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18348_ _18845_/A0 _10330_/Y _18884_/S vssd1 vssd1 vccd1 vccd1 _18348_/X sky130_fd_sc_hd__mux2_1
XFILLER_187_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10589__B2 _10588_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18279_ _19186_/X _21274_/Q _18281_/S vssd1 vssd1 vccd1 vccd1 _18279_/X sky130_fd_sc_hd__mux2_1
XFILLER_135_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12815__A _12815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20310_ _20316_/CLK _20310_/D repeater197/X vssd1 vssd1 vccd1 vccd1 _20310_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_238_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput50 HWDATA[20] vssd1 vssd1 vccd1 vccd1 input50/X sky130_fd_sc_hd__buf_2
X_21290_ _21349_/CLK _21290_/D repeater210/X vssd1 vssd1 vccd1 vccd1 _21290_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_163_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput61 HWDATA[30] vssd1 vssd1 vccd1 vccd1 input61/X sky130_fd_sc_hd__buf_4
Xinput72 MSI_S3 vssd1 vssd1 vccd1 vccd1 input72/X sky130_fd_sc_hd__buf_2
XANTENNA__11538__B1 _10898_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_238_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20241_ _20241_/CLK _20241_/D repeater248/X vssd1 vssd1 vccd1 vccd1 _20241_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_143_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20172_ _20172_/CLK _20172_/D repeater248/X vssd1 vssd1 vccd1 vccd1 _20172_/Q sky130_fd_sc_hd__dfrtp_1
X_09983_ _20016_/Q _20017_/Q _20018_/Q _20019_/Q vssd1 vssd1 vccd1 vccd1 _10013_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_115_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12550__A _12550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18648__S _18906_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13463__B1 _13270_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18383__S _18910_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13766__A1 _20612_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18154__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11310_ _11543_/A _11310_/B _11310_/C _11310_/D vssd1 vssd1 vccd1 vccd1 _12503_/B
+ sky130_fd_sc_hd__nor4_2
XFILLER_148_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14715__B1 _13584_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20508_ _20947_/CLK _20508_/D repeater266/X vssd1 vssd1 vccd1 vccd1 _20508_/Q sky130_fd_sc_hd__dfrtp_4
X_12290_ _20500_/Q vssd1 vssd1 vccd1 vccd1 _12290_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11241_ _11241_/A vssd1 vssd1 vccd1 vccd1 _11241_/Y sky130_fd_sc_hd__inv_2
X_20439_ _20476_/CLK _20439_/D repeater279/X vssd1 vssd1 vccd1 vccd1 _20439_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_107_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20718__RESET_B repeater254/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11172_ _16465_/B _11172_/B vssd1 vssd1 vccd1 vccd1 _11173_/B sky130_fd_sc_hd__or2_1
XFILLER_164_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17028__A _21248_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10123_ _20778_/Q vssd1 vssd1 vccd1 vccd1 _10123_/Y sky130_fd_sc_hd__inv_2
XFILLER_164_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15980_ _19545_/Q _15978_/X _15944_/X _15979_/X vssd1 vssd1 vccd1 vccd1 _19545_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_input33_A HREADY vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14931_ _20587_/Q _14835_/A _20586_/Q _14960_/A vssd1 vssd1 vccd1 vccd1 _14931_/X
+ sky130_fd_sc_hd__o22a_1
X_10054_ _21391_/Q vssd1 vssd1 vccd1 vccd1 _10152_/A sky130_fd_sc_hd__inv_2
XANTENNA__18558__S _18835_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_125_HCLK_A clkbuf_4_4_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_236_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17650_ _21141_/Q vssd1 vssd1 vccd1 vccd1 _17650_/Y sky130_fd_sc_hd__inv_2
X_14862_ _20086_/Q vssd1 vssd1 vccd1 vccd1 _15006_/A sky130_fd_sc_hd__inv_2
XFILLER_91_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16601_ _19993_/Q _19995_/Q _19996_/Q _19992_/Q vssd1 vssd1 vccd1 vccd1 _16603_/C
+ sky130_fd_sc_hd__or4_4
X_13813_ _20602_/Q vssd1 vssd1 vccd1 vccd1 _13813_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17581_ _17581_/A vssd1 vssd1 vccd1 vccd1 _17820_/A sky130_fd_sc_hd__inv_2
X_14793_ _20242_/Q _16480_/A vssd1 vssd1 vccd1 vccd1 _14794_/A sky130_fd_sc_hd__or2_2
XANTENNA__14387__A _20030_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16532_ _19881_/Q vssd1 vssd1 vccd1 vccd1 _16602_/A sky130_fd_sc_hd__inv_2
X_19320_ _21449_/CLK _19320_/D vssd1 vssd1 vccd1 vccd1 _19320_/Q sky130_fd_sc_hd__dfxtp_1
X_13744_ _20622_/Q vssd1 vssd1 vccd1 vccd1 _13744_/Y sky130_fd_sc_hd__inv_2
XFILLER_188_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10956_ _21210_/Q vssd1 vssd1 vccd1 vccd1 _10956_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18393__A0 _18848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_216_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19251_ _19247_/X _19248_/X _19249_/X _19250_/X _20132_/Q _20133_/Q vssd1 vssd1 vccd1
+ vccd1 _19251_/X sky130_fd_sc_hd__mux4_2
X_16463_ _19301_/Q _16459_/X _16340_/X _16460_/X vssd1 vssd1 vccd1 vccd1 _19301_/D
+ sky130_fd_sc_hd__a22o_1
X_13675_ _20355_/Q _13673_/X _13560_/X _13674_/X vssd1 vssd1 vccd1 vccd1 _20355_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18293__S _18903_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_232_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_repeater172_A _18775_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10887_ _21256_/Q _10879_/X _10886_/X _10881_/X vssd1 vssd1 vccd1 vccd1 _21256_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_231_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15414_ _15528_/A _15655_/B _15778_/C vssd1 vssd1 vccd1 vccd1 _15423_/A sky130_fd_sc_hd__or3_4
X_18202_ _18848_/A0 _10296_/Y _18884_/S vssd1 vssd1 vccd1 vccd1 _18202_/X sky130_fd_sc_hd__mux2_1
XPHY_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12626_ _12638_/A vssd1 vssd1 vccd1 vccd1 _12626_/X sky130_fd_sc_hd__buf_1
X_19182_ _19706_/Q _19570_/Q _19562_/Q _19554_/Q _19280_/S0 _20122_/Q vssd1 vssd1
+ vccd1 vccd1 _19182_/X sky130_fd_sc_hd__mux4_2
XPHY_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16394_ _16400_/A vssd1 vssd1 vccd1 vccd1 _16394_/X sky130_fd_sc_hd__buf_1
XANTENNA__18145__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18133_ _18132_/X _14591_/A _18748_/S vssd1 vssd1 vccd1 vccd1 _18133_/X sky130_fd_sc_hd__mux2_1
X_15345_ _15345_/A vssd1 vssd1 vccd1 vccd1 _15345_/X sky130_fd_sc_hd__buf_1
X_12557_ _20894_/Q _12553_/X _11741_/X _12554_/X vssd1 vssd1 vccd1 vccd1 _20894_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_8_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11508_ _21147_/Q vssd1 vssd1 vccd1 vccd1 _11508_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18064_ _18064_/A vssd1 vssd1 vccd1 vccd1 _18064_/X sky130_fd_sc_hd__buf_1
XFILLER_145_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15276_ _20469_/Q vssd1 vssd1 vccd1 vccd1 _17540_/A sky130_fd_sc_hd__inv_2
X_12488_ _12488_/A vssd1 vssd1 vccd1 vccd1 _12492_/A sky130_fd_sc_hd__inv_2
X_17015_ _19980_/Q _17008_/A _19981_/Q vssd1 vssd1 vccd1 vccd1 _17015_/X sky130_fd_sc_hd__o21a_1
XFILLER_172_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14227_ _14072_/A _14072_/B _14225_/Y _14185_/X vssd1 vssd1 vccd1 vccd1 _20261_/D
+ sky130_fd_sc_hd__a211oi_2
X_11439_ _11439_/A vssd1 vssd1 vccd1 vccd1 _21168_/D sky130_fd_sc_hd__inv_2
XFILLER_160_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20459__RESET_B repeater276/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14158_ _20534_/Q _14074_/A _14156_/Y _20262_/Q _14157_/X vssd1 vssd1 vccd1 vccd1
+ _14170_/A sky130_fd_sc_hd__o221a_1
XFILLER_112_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13109_ _12978_/X _20631_/Q _13109_/S vssd1 vssd1 vccd1 vccd1 _20631_/D sky130_fd_sc_hd__mux2_1
XANTENNA__13466__A _13481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18966_ _14309_/B _14307_/C _18976_/S vssd1 vssd1 vccd1 vccd1 _18966_/X sky130_fd_sc_hd__mux2_1
X_14089_ _14089_/A _14089_/B vssd1 vssd1 vccd1 vccd1 _14195_/A sky130_fd_sc_hd__or2_1
XFILLER_239_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17917_ _18477_/X _18020_/A _18460_/X _17326_/X vssd1 vssd1 vccd1 vccd1 _17917_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__18468__S _18897_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18897_ _18896_/X _14414_/Y _18897_/S vssd1 vssd1 vccd1 vccd1 _18897_/X sky130_fd_sc_hd__mux2_1
XANTENNA__16777__A _16777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17848_ _20342_/Q vssd1 vssd1 vccd1 vccd1 _17848_/Y sky130_fd_sc_hd__inv_2
XFILLER_94_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17779_ _20404_/Q vssd1 vssd1 vccd1 vccd1 _17779_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19685__CLK _19813_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_47_HCLK_A _20004_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_241_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19518_ _19521_/CLK _19518_/D vssd1 vssd1 vccd1 vccd1 _19518_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_240_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18384__A0 _17079_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20790_ _21374_/CLK _20790_/D repeater255/X vssd1 vssd1 vccd1 vccd1 _20790_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__21247__RESET_B repeater233/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19449_ _20137_/CLK _19449_/D vssd1 vssd1 vccd1 vccd1 _19449_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__18136__A0 _17079_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21411_ _21417_/CLK _21411_/D repeater234/X vssd1 vssd1 vccd1 vccd1 _21411_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_148_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21342_ _21342_/CLK _21342_/D repeater211/X vssd1 vssd1 vccd1 vccd1 _21342_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_162_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15370__B1 _15352_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21273_ _21273_/CLK _21273_/D repeater245/X vssd1 vssd1 vccd1 vccd1 _21273_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_162_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20224_ _21484_/CLK _20224_/D repeater202/X vssd1 vssd1 vccd1 vccd1 _20224_/Q sky130_fd_sc_hd__dfrtp_4
X_20155_ _21242_/CLK _20155_/D repeater189/X vssd1 vssd1 vccd1 vccd1 _20155_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_89_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09966_ _10877_/A _15312_/A _12605_/A _10026_/B vssd1 vssd1 vccd1 vccd1 _09969_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_58_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20086_ _20495_/CLK _20086_/D repeater273/X vssd1 vssd1 vccd1 vccd1 _20086_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__18378__S _18880_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13684__B1 _13489_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09897_ _17024_/A vssd1 vssd1 vccd1 vccd1 _09897_/Y sky130_fd_sc_hd__inv_2
XFILLER_245_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_4_15_0_HCLK_A clkbuf_3_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10810_ _10771_/A _10771_/B _10809_/X _10807_/Y vssd1 vssd1 vccd1 vccd1 _21295_/D
+ sky130_fd_sc_hd__a211oi_2
XPHY_3912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11790_ input33/X hold9/A vssd1 vssd1 vccd1 vccd1 _11794_/A sky130_fd_sc_hd__nand2_4
XPHY_3934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20988_ _21319_/CLK _20988_/D repeater191/X vssd1 vssd1 vccd1 vccd1 _20988_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_214_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10741_ _19929_/Q _16790_/A vssd1 vssd1 vccd1 vccd1 _16794_/A sky130_fd_sc_hd__or2_2
XPHY_3967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19002__S _19019_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13460_ _13493_/A vssd1 vssd1 vccd1 vccd1 _13483_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_41_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_230_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10672_ _10672_/A vssd1 vssd1 vccd1 vccd1 _10672_/Y sky130_fd_sc_hd__inv_2
X_12411_ _12462_/A vssd1 vssd1 vccd1 vccd1 _12411_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__19408__CLK _19813_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13391_ _13416_/A vssd1 vssd1 vccd1 vccd1 _13419_/A sky130_fd_sc_hd__inv_2
XANTENNA__18841__S _18841_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15130_ _20455_/Q _15129_/X _20455_/Q _15129_/X vssd1 vssd1 vccd1 vccd1 _15130_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_12342_ _12342_/A vssd1 vssd1 vccd1 vccd1 _12342_/Y sky130_fd_sc_hd__inv_2
XFILLER_182_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_opt_2_HCLK clkbuf_opt_2_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_opt_2_HCLK/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_126_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15061_ _15061_/A _15061_/B vssd1 vssd1 vccd1 vccd1 _15211_/A sky130_fd_sc_hd__or2_1
XANTENNA__15766__A _15766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12273_ _20523_/Q vssd1 vssd1 vccd1 vccd1 _12273_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19558__CLK _19706_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14012_ _14012_/A _14026_/A vssd1 vssd1 vccd1 vccd1 _14013_/B sky130_fd_sc_hd__or2_1
XFILLER_141_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11224_ _21201_/Q _11219_/X _10892_/X _11220_/X vssd1 vssd1 vccd1 vccd1 _21201_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_108_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18820_ _17079_/Y _12137_/Y _18908_/S vssd1 vssd1 vccd1 vccd1 _18820_/X sky130_fd_sc_hd__mux2_1
XFILLER_122_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11155_ _20598_/Q vssd1 vssd1 vccd1 vccd1 _13182_/A sky130_fd_sc_hd__inv_2
XFILLER_150_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10106_ _20792_/Q vssd1 vssd1 vccd1 vccd1 _10106_/Y sky130_fd_sc_hd__inv_2
X_18751_ _17540_/Y _20437_/Q _18909_/S vssd1 vssd1 vccd1 vccd1 _18751_/X sky130_fd_sc_hd__mux2_2
XFILLER_48_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11086_ _21234_/Q _11086_/B vssd1 vssd1 vccd1 vccd1 _11086_/Y sky130_fd_sc_hd__nor2_1
X_15963_ _19553_/Q _15961_/X _15944_/X _15962_/X vssd1 vssd1 vccd1 vccd1 _19553_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_110_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13675__B1 _13560_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18288__S _18667_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17702_ _19315_/Q _17829_/B vssd1 vssd1 vccd1 vccd1 _17702_/X sky130_fd_sc_hd__and2_1
XANTENNA__18063__C1 _18062_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14914_ _20565_/Q vssd1 vssd1 vccd1 vccd1 _14914_/Y sky130_fd_sc_hd__inv_2
X_10037_ _21379_/Q vssd1 vssd1 vccd1 vccd1 _10041_/A sky130_fd_sc_hd__inv_2
X_18682_ _18681_/X _16774_/A _18880_/S vssd1 vssd1 vccd1 vccd1 _18682_/X sky130_fd_sc_hd__mux2_1
X_15894_ _19587_/Q _15886_/X _15893_/X _15889_/X vssd1 vssd1 vccd1 vccd1 _19587_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_208_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17633_ _21436_/Q _17776_/B vssd1 vssd1 vccd1 vccd1 _17633_/Y sky130_fd_sc_hd__nand2_1
XFILLER_208_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13427__B1 _13426_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14845_ _14845_/A vssd1 vssd1 vccd1 vccd1 _14962_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_63_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17564_ _20897_/Q vssd1 vssd1 vccd1 vccd1 _17564_/Y sky130_fd_sc_hd__inv_2
X_14776_ _16451_/B vssd1 vssd1 vccd1 vccd1 _15967_/B sky130_fd_sc_hd__buf_1
XFILLER_210_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11988_ _11988_/A vssd1 vssd1 vccd1 vccd1 _20999_/D sky130_fd_sc_hd__inv_2
X_19303_ _20172_/CLK _19303_/D vssd1 vssd1 vccd1 vccd1 _19303_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13727_ _13727_/A vssd1 vssd1 vccd1 vccd1 _13734_/S sky130_fd_sc_hd__clkbuf_2
X_16515_ _16515_/A _16525_/B vssd1 vssd1 vccd1 vccd1 _16515_/Y sky130_fd_sc_hd__nor2_1
X_10939_ _21037_/Q vssd1 vssd1 vccd1 vccd1 _11814_/A sky130_fd_sc_hd__inv_2
X_17495_ _19722_/Q vssd1 vssd1 vccd1 vccd1 _17495_/Y sky130_fd_sc_hd__inv_2
XFILLER_71_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19234_ _17492_/Y _17493_/Y _17494_/Y _17495_/Y _19275_/S0 _21004_/Q vssd1 vssd1
+ vccd1 vccd1 _19234_/X sky130_fd_sc_hd__mux4_2
X_13658_ _13685_/A vssd1 vssd1 vccd1 vccd1 _13679_/A sky130_fd_sc_hd__clkbuf_2
X_16446_ _19309_/Q _16441_/X _16342_/X _16442_/X vssd1 vssd1 vccd1 vccd1 _19309_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_176_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18036__B _18084_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12609_ _20867_/Q _12574_/A _18219_/X _12575_/A vssd1 vssd1 vccd1 vccd1 _20867_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18669__A1 _14442_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19165_ _19300_/Q _19822_/Q _19830_/Q _19414_/Q _19280_/S0 _20122_/Q vssd1 vssd1
+ vccd1 vccd1 _19165_/X sky130_fd_sc_hd__mux4_2
XFILLER_31_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16377_ _16419_/A _16419_/B _16377_/C vssd1 vssd1 vccd1 vccd1 _16385_/A sky130_fd_sc_hd__or3_4
X_13589_ _13595_/A vssd1 vssd1 vccd1 vccd1 _13589_/X sky130_fd_sc_hd__buf_1
XANTENNA__18751__S _18909_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18116_ vssd1 vssd1 vccd1 vccd1 _18218_/A1 _18116_/LO sky130_fd_sc_hd__conb_1
X_15328_ _20028_/Q _15323_/X _13550_/X _15324_/X vssd1 vssd1 vccd1 vccd1 _20028_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_191_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19096_ _16674_/X _21082_/Q _19870_/D vssd1 vssd1 vccd1 vccd1 _19096_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15259_ _15259_/A _15259_/B _15259_/C _15258_/X vssd1 vssd1 vccd1 vccd1 _15259_/X
+ sky130_fd_sc_hd__or4b_4
X_18047_ _18326_/X _18019_/X _18264_/X _18020_/X _18046_/X vssd1 vssd1 vccd1 vccd1
+ _18051_/B sky130_fd_sc_hd__o221a_2
XFILLER_144_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20293__RESET_B repeater263/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09674__A input66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19094__A1 _21084_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20222__RESET_B repeater202/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09820_ _21451_/Q vssd1 vssd1 vccd1 vccd1 _15871_/A sky130_fd_sc_hd__buf_1
X_19998_ _20042_/CLK _19998_/D repeater219/X vssd1 vssd1 vccd1 vccd1 _19998_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_247_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09751_ _21237_/Q vssd1 vssd1 vccd1 vccd1 _11062_/A sky130_fd_sc_hd__inv_2
X_18949_ _16662_/X _21087_/Q _18962_/S vssd1 vssd1 vccd1 vccd1 _18949_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13666__B1 _13547_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18198__S _18666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09682_ _12550_/A vssd1 vssd1 vccd1 vccd1 _09682_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_104_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20911_ _20915_/CLK _20911_/D repeater218/X vssd1 vssd1 vccd1 vccd1 _20911_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_243_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18926__S _18926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_242_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20842_ _21374_/CLK _20842_/D repeater255/X vssd1 vssd1 vccd1 vccd1 _20842_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_35_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21010__RESET_B repeater238/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20773_ _21379_/CLK _20773_/D repeater213/X vssd1 vssd1 vccd1 vccd1 _20773_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_211_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14755__A _20133_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15591__B1 _15590_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18661__S _18909_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21325_ _21476_/CLK _21325_/D repeater204/X vssd1 vssd1 vccd1 vccd1 _21325_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_2_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20558__CLK _20592_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21256_ _21390_/CLK _21256_/D repeater239/X vssd1 vssd1 vccd1 vccd1 _21256_/Q sky130_fd_sc_hd__dfrtp_1
X_20207_ _20622_/CLK _20207_/D repeater195/X vssd1 vssd1 vccd1 vccd1 _20207_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__19180__S1 _20122_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21187_ _21193_/CLK _21187_/D repeater224/X vssd1 vssd1 vccd1 vccd1 _21187_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_132_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20138_ _21218_/CLK _20138_/D repeater242/X vssd1 vssd1 vccd1 vccd1 _20138_/Q sky130_fd_sc_hd__dfrtp_1
X_09949_ _10026_/B _13384_/C vssd1 vssd1 vccd1 vccd1 _09957_/A sky130_fd_sc_hd__or2_2
XFILLER_86_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20069_ _20070_/CLK _20069_/D repeater276/X vssd1 vssd1 vccd1 vccd1 _20069_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_58_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12960_ _12960_/A vssd1 vssd1 vccd1 vccd1 _12960_/X sky130_fd_sc_hd__buf_1
XANTENNA__21169__RESET_B repeater220/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11132__A1 _21005_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11911_ _15375_/A _11003_/X _11906_/Y _15397_/A _11910_/X vssd1 vssd1 vccd1 vccd1
+ _21015_/D sky130_fd_sc_hd__a32o_1
X_12891_ _13600_/A vssd1 vssd1 vccd1 vccd1 _12891_/X sky130_fd_sc_hd__buf_1
XPHY_4410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18836__S _18875_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14630_ _14630_/A vssd1 vssd1 vccd1 vccd1 _14630_/Y sky130_fd_sc_hd__inv_2
XPHY_4443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11842_ _21033_/Q _11842_/B vssd1 vssd1 vccd1 vccd1 _11842_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10891__B1 _10889_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18348__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_30_HCLK_A clkbuf_opt_4_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14561_ _14561_/A vssd1 vssd1 vccd1 vccd1 _14561_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11773_ _19088_/X _11770_/X _21046_/Q _11771_/X vssd1 vssd1 vccd1 vccd1 _21046_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_60_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_93_HCLK_A clkbuf_4_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13512_ _20438_/Q _13505_/X _13511_/X _13507_/X vssd1 vssd1 vccd1 vccd1 _20438_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_41_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16300_ _16306_/A vssd1 vssd1 vccd1 vccd1 _16300_/X sky130_fd_sc_hd__buf_1
XPHY_3786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10724_ _10540_/B _10726_/A _10540_/A vssd1 vssd1 vccd1 vccd1 _10725_/B sky130_fd_sc_hd__o21a_1
XFILLER_159_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17280_ _17449_/A _20110_/Q vssd1 vssd1 vccd1 vccd1 _17280_/X sky130_fd_sc_hd__and2_1
X_14492_ _14462_/B _14366_/B _14490_/Y _14488_/X vssd1 vssd1 vccd1 vccd1 _20223_/D
+ sky130_fd_sc_hd__a211oi_2
XPHY_3797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16231_ _16231_/A vssd1 vssd1 vccd1 vccd1 _16231_/X sky130_fd_sc_hd__buf_2
X_13443_ _20469_/Q _13436_/X _13442_/X _13437_/X vssd1 vssd1 vccd1 vccd1 _20469_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11801__B _12968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10655_ _10655_/A _10655_/B vssd1 vssd1 vccd1 vccd1 _10690_/A sky130_fd_sc_hd__or2_1
XANTENNA__18571__S _18666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20733__RESET_B repeater257/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16162_ _19455_/Q _16158_/X _16147_/X _16159_/X vssd1 vssd1 vccd1 vccd1 _19455_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_6_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13374_ _20504_/Q _13371_/X _13243_/X _13372_/X vssd1 vssd1 vccd1 vccd1 _20504_/D
+ sky130_fd_sc_hd__a22o_1
X_10586_ _21322_/Q _10584_/Y _21315_/Q _10585_/Y vssd1 vssd1 vccd1 vccd1 _10586_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_154_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15113_ _20443_/Q _15068_/A _20453_/Q _15112_/X vssd1 vssd1 vccd1 vccd1 _15113_/X
+ sky130_fd_sc_hd__a22o_1
X_12325_ _12325_/A _12325_/B vssd1 vssd1 vccd1 vccd1 _12352_/A sky130_fd_sc_hd__or2_1
X_16093_ _16093_/A _16165_/B _16405_/C vssd1 vssd1 vccd1 vccd1 _16101_/A sky130_fd_sc_hd__or3_4
XFILLER_115_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19921_ _21379_/CLK _19921_/D repeater211/X vssd1 vssd1 vccd1 vccd1 _19921_/Q sky130_fd_sc_hd__dfrtp_1
X_15044_ _20058_/Q vssd1 vssd1 vccd1 vccd1 _15099_/A sky130_fd_sc_hd__inv_2
XFILLER_108_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12256_ _12256_/A vssd1 vssd1 vccd1 vccd1 _12472_/A sky130_fd_sc_hd__clkbuf_2
X_11207_ _11207_/A vssd1 vssd1 vccd1 vccd1 _11226_/A sky130_fd_sc_hd__inv_2
X_19852_ _21424_/CLK _19852_/D repeater229/X vssd1 vssd1 vccd1 vccd1 _19852_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__19171__S1 _20124_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12187_ _20355_/Q vssd1 vssd1 vccd1 vccd1 _12187_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18803_ _18845_/A0 _17373_/Y _18879_/S vssd1 vssd1 vccd1 vccd1 _18803_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11138_ _19116_/X vssd1 vssd1 vccd1 vccd1 _11138_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13648__B1 _13509_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19783_ _19828_/CLK _19783_/D vssd1 vssd1 vccd1 vccd1 _19783_/Q sky130_fd_sc_hd__dfxtp_1
X_16995_ _16999_/B _16994_/Y _16967_/X vssd1 vssd1 vccd1 vccd1 _16995_/X sky130_fd_sc_hd__o21a_1
XFILLER_96_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18734_ _18733_/X _17630_/Y _18929_/S vssd1 vssd1 vccd1 vccd1 _18734_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15946_ _19561_/Q _15943_/X _15944_/X _15945_/X vssd1 vssd1 vccd1 vccd1 _19561_/D
+ sky130_fd_sc_hd__a22o_1
X_11069_ _11069_/A vssd1 vssd1 vccd1 vccd1 _21239_/D sky130_fd_sc_hd__inv_2
XFILLER_64_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18587__A0 _18586_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_225_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19987__RESET_B repeater218/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18665_ _18848_/A0 _10317_/Y _18884_/S vssd1 vssd1 vccd1 vccd1 _18665_/X sky130_fd_sc_hd__mux2_1
XFILLER_92_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11674__A2 _11657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18746__S _18880_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15877_ _15877_/A vssd1 vssd1 vccd1 vccd1 _15877_/X sky130_fd_sc_hd__buf_1
XFILLER_224_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17616_ _19611_/Q vssd1 vssd1 vccd1 vccd1 _17616_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10882__B1 _09663_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_221_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19916__RESET_B repeater220/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14828_ _20104_/Q vssd1 vssd1 vccd1 vccd1 _14881_/A sky130_fd_sc_hd__inv_2
XFILLER_17_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18596_ _18595_/X _12264_/Y _18910_/S vssd1 vssd1 vccd1 vccd1 _18596_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_130_HCLK clkbuf_4_4_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20428_/CLK sky130_fd_sc_hd__clkbuf_16
X_17547_ _20401_/Q _18835_/S vssd1 vssd1 vccd1 vccd1 _17547_/Y sky130_fd_sc_hd__nand2_1
XFILLER_63_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14759_ _14535_/Y _14758_/Y _14754_/Y vssd1 vssd1 vccd1 vccd1 _20132_/D sky130_fd_sc_hd__a21oi_1
XFILLER_232_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17478_ _18788_/X _17401_/X _18795_/X _17320_/X vssd1 vssd1 vccd1 vccd1 _17478_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_20_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19217_ _17611_/Y _17612_/Y _17613_/Y _17614_/Y _20130_/Q _20131_/Q vssd1 vssd1 vccd1
+ vccd1 _19217_/X sky130_fd_sc_hd__mux4_1
X_16429_ _19320_/Q _16427_/X _15876_/A _16428_/X vssd1 vssd1 vccd1 vccd1 _19320_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18481__S _18884_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19148_ _19762_/Q _19754_/Q _19746_/Q _19738_/Q _19285_/S0 _21017_/Q vssd1 vssd1
+ vccd1 vccd1 _19148_/X sky130_fd_sc_hd__mux4_2
XANTENNA__18511__A0 _17281_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15325__B1 _13543_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19079_ _16724_/X _20896_/Q _19908_/D vssd1 vssd1 vccd1 vccd1 _19079_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21110_ _21417_/CLK _21110_/D repeater231/X vssd1 vssd1 vccd1 vccd1 _21110_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_117_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19067__A1 _21143_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12542__B _14273_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21041_ _21183_/CLK _21041_/D repeater219/X vssd1 vssd1 vccd1 vccd1 _21041_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__19162__S1 _20122_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09803_ _09803_/A vssd1 vssd1 vccd1 vccd1 _09806_/A sky130_fd_sc_hd__buf_1
XFILLER_219_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09734_ _20149_/Q vssd1 vssd1 vccd1 vccd1 _09734_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09665_ input68/X vssd1 vssd1 vccd1 vccd1 _13313_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_39_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18656__S _18910_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_199_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10873__B1 _09688_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09596_ _20889_/Q vssd1 vssd1 vccd1 vccd1 _13047_/B sky130_fd_sc_hd__buf_1
XPHY_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20825_ _20841_/CLK _20825_/D repeater256/X vssd1 vssd1 vccd1 vccd1 _20825_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20756_ _21481_/CLK _20756_/D repeater205/X vssd1 vssd1 vccd1 vccd1 _20756_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12717__B _13104_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18391__S _18784_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15564__B1 _15544_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10518__A _20697_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20687_ _21302_/CLK _20687_/D repeater209/X vssd1 vssd1 vccd1 vccd1 _20687_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10440_ _21284_/Q vssd1 vssd1 vccd1 vccd1 _10761_/A sky130_fd_sc_hd__inv_2
XFILLER_155_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18502__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20144__RESET_B repeater250/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10371_ _10287_/A _10287_/B _10369_/Y _10405_/B vssd1 vssd1 vccd1 vccd1 _21372_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_109_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12110_ _20956_/Q _12107_/Y _12109_/X _20368_/Q vssd1 vssd1 vccd1 vccd1 _12110_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_124_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21308_ _21481_/CLK _21308_/D repeater206/X vssd1 vssd1 vccd1 vccd1 _21308_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_156_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13090_ _20643_/Q _13086_/X _13030_/X _13087_/X vssd1 vssd1 vccd1 vccd1 _20643_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_3_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_11_HCLK clkbuf_opt_2_HCLK/A vssd1 vssd1 vccd1 vccd1 _21009_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_156_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12041_ _12036_/X _20378_/Q _20968_/Q _12037_/Y _12040_/X vssd1 vssd1 vccd1 vccd1
+ _12060_/A sky130_fd_sc_hd__o221a_1
XANTENNA__19153__S1 _21017_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21239_ _21239_/CLK _21239_/D repeater251/X vssd1 vssd1 vccd1 vccd1 _21239_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_2_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15800_ _15807_/A vssd1 vssd1 vccd1 vccd1 _15800_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_172_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16780_ _16777_/Y _16778_/Y _16779_/X vssd1 vssd1 vccd1 vccd1 _16780_/X sky130_fd_sc_hd__o21a_1
X_13992_ _13974_/B _13889_/B _13986_/Y _13991_/X vssd1 vssd1 vccd1 vccd1 _20313_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_207_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_153_HCLK clkbuf_opt_1_HCLK/A vssd1 vssd1 vccd1 vccd1 _21449_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_58_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15731_ _19660_/Q _15723_/X _15730_/X _15727_/X vssd1 vssd1 vccd1 vccd1 _19660_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_74_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12943_ _12961_/A vssd1 vssd1 vccd1 vccd1 _12943_/X sky130_fd_sc_hd__buf_1
XFILLER_207_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18566__S _18906_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18450_ _18449_/X _10126_/Y _18885_/S vssd1 vssd1 vccd1 vccd1 _18450_/X sky130_fd_sc_hd__mux2_1
X_12874_ _12874_/A vssd1 vssd1 vccd1 vccd1 _12874_/X sky130_fd_sc_hd__buf_1
XFILLER_34_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15662_ _19692_/Q _15656_/X _15661_/X _15659_/X vssd1 vssd1 vccd1 vccd1 _19692_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19746__CLK _19765_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17401_ _17581_/A vssd1 vssd1 vccd1 vccd1 _17401_/X sky130_fd_sc_hd__buf_1
XPHY_4273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14613_ _14613_/A vssd1 vssd1 vccd1 vccd1 _14613_/Y sky130_fd_sc_hd__inv_2
X_11825_ _21037_/Q _11825_/B vssd1 vssd1 vccd1 vccd1 _11825_/X sky130_fd_sc_hd__or2_1
XFILLER_233_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output102_A _18097_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18381_ _17079_/Y _12131_/Y _18908_/S vssd1 vssd1 vccd1 vccd1 _18381_/X sky130_fd_sc_hd__mux2_1
X_15593_ _19726_/Q _15584_/X _15592_/X _15586_/X vssd1 vssd1 vccd1 vccd1 _19726_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20914__RESET_B repeater218/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14544_ _14536_/X _14541_/Y _14561_/A vssd1 vssd1 vccd1 vccd1 _14544_/X sky130_fd_sc_hd__o21a_1
X_17332_ _19696_/Q vssd1 vssd1 vccd1 vccd1 _17332_/Y sky130_fd_sc_hd__inv_2
X_11756_ _21054_/Q _11755_/A _11754_/Y _11755_/Y _19872_/Q vssd1 vssd1 vccd1 vccd1
+ _21054_/D sky130_fd_sc_hd__a221o_1
XPHY_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10707_ _10707_/A _10711_/A vssd1 vssd1 vccd1 vccd1 _10708_/B sky130_fd_sc_hd__or2_2
XPHY_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14475_ _14465_/B _14376_/B _14471_/Y _14474_/X vssd1 vssd1 vccd1 vccd1 _20233_/D
+ sky130_fd_sc_hd__a211oi_2
XPHY_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17263_ _19591_/Q vssd1 vssd1 vccd1 vccd1 _17263_/Y sky130_fd_sc_hd__inv_2
XFILLER_186_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11687_ _21085_/Q _11679_/X _11686_/X _11682_/X vssd1 vssd1 vccd1 vccd1 _21085_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_repeater252_A repeater255/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19002_ _16990_/X _20421_/Q _19019_/S vssd1 vssd1 vccd1 vccd1 _19974_/D sky130_fd_sc_hd__mux2_1
XFILLER_201_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16214_ _19430_/Q _16206_/X _16163_/X _16208_/X vssd1 vssd1 vccd1 vccd1 _19430_/D
+ sky130_fd_sc_hd__a22o_1
X_13426_ input41/X vssd1 vssd1 vccd1 vccd1 _13426_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_128_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10638_ _10625_/X _10638_/B _10638_/C _10638_/D vssd1 vssd1 vccd1 vccd1 _10639_/D
+ sky130_fd_sc_hd__and4b_1
X_17194_ _18920_/X vssd1 vssd1 vccd1 vccd1 _17194_/Y sky130_fd_sc_hd__inv_2
X_16145_ _21448_/Q vssd1 vssd1 vccd1 vccd1 _16145_/X sky130_fd_sc_hd__clkbuf_2
X_13357_ _13357_/A vssd1 vssd1 vccd1 vccd1 _13377_/A sky130_fd_sc_hd__buf_1
X_10569_ _10569_/A vssd1 vssd1 vccd1 vccd1 _10661_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_182_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12308_ _12308_/A _12308_/B vssd1 vssd1 vccd1 vccd1 _12383_/A sky130_fd_sc_hd__or2_1
X_16076_ _19494_/Q _16071_/X _15776_/X _16072_/X vssd1 vssd1 vccd1 vccd1 _19494_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_170_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13288_ _13294_/A vssd1 vssd1 vccd1 vccd1 _13288_/X sky130_fd_sc_hd__buf_1
XFILLER_108_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19904_ _19904_/CLK input76/X repeater202/X vssd1 vssd1 vccd1 vccd1 _19905_/D sky130_fd_sc_hd__dfrtp_1
X_15027_ _20074_/Q vssd1 vssd1 vccd1 vccd1 _15088_/A sky130_fd_sc_hd__inv_2
XANTENNA__15954__A _15961_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12239_ _20506_/Q vssd1 vssd1 vccd1 vccd1 _12239_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19144__S1 _21017_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19835_ _19835_/CLK _19835_/D vssd1 vssd1 vccd1 vccd1 _19835_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19766_ _19828_/CLK _19766_/D vssd1 vssd1 vccd1 vccd1 _19766_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13097__A1 _20638_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16978_ _19972_/Q vssd1 vssd1 vccd1 vccd1 _16978_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput4 HADDR[12] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_1
X_18717_ _18716_/X _10585_/Y _18879_/S vssd1 vssd1 vccd1 vccd1 _18717_/X sky130_fd_sc_hd__mux2_1
X_15929_ _19569_/Q _15927_/X _15788_/X _15928_/X vssd1 vssd1 vccd1 vccd1 _19569_/D
+ sky130_fd_sc_hd__a22o_1
X_19697_ _20326_/CLK _19697_/D vssd1 vssd1 vccd1 vccd1 _19697_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__18476__S _18903_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_237_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18648_ _18647_/X _18098_/Y _18906_/S vssd1 vssd1 vccd1 vccd1 _18648_/X sky130_fd_sc_hd__mux2_1
XFILLER_91_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_225_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18579_ _18845_/A0 _13802_/Y _18896_/S vssd1 vssd1 vccd1 vccd1 _18579_/X sky130_fd_sc_hd__mux2_1
XANTENNA__15794__B1 _15793_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_212_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20610_ _20657_/CLK _20610_/D repeater198/X vssd1 vssd1 vccd1 vccd1 _20610_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_177_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20541_ _20592_/CLK _20541_/D repeater265/X vssd1 vssd1 vccd1 vccd1 _20541_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_220_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19100__S _19870_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20472_ _20937_/CLK _20472_/D repeater279/X vssd1 vssd1 vccd1 vccd1 _20472_/Q sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_34_HCLK clkbuf_opt_4_HCLK/X vssd1 vssd1 vccd1 vccd1 _20331_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__12780__B1 _09633_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19135__S1 _21017_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21024_ _21255_/CLK _21024_/D repeater241/X vssd1 vssd1 vccd1 vccd1 _21024_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_248_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13384__A _17177_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09717_ _09787_/B vssd1 vssd1 vccd1 vccd1 _16617_/B sky130_fd_sc_hd__inv_2
XFILLER_56_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18386__S _18910_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09648_ input42/X vssd1 vssd1 vccd1 vccd1 _12855_/A sky130_fd_sc_hd__buf_4
XANTENNA__20746__CLK _21342_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11610_ _21408_/Q vssd1 vssd1 vccd1 vccd1 _11636_/A sky130_fd_sc_hd__inv_2
XPHY_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20808_ _21242_/CLK _20808_/D repeater189/X vssd1 vssd1 vccd1 vccd1 _20808_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_168_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12590_ _20880_/Q _12588_/X _18232_/X _12589_/X vssd1 vssd1 vccd1 vccd1 _20880_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20325__RESET_B repeater250/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11541_ _11541_/A _11541_/B _11541_/C vssd1 vssd1 vccd1 vccd1 _11542_/A sky130_fd_sc_hd__or3_1
XFILLER_184_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20739_ _21321_/CLK _20739_/D repeater205/X vssd1 vssd1 vccd1 vccd1 _20739_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_168_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19010__S _19019_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14260_ _14268_/A vssd1 vssd1 vccd1 vccd1 _14260_/X sky130_fd_sc_hd__buf_1
X_11472_ _19097_/X _11468_/X _21161_/Q _11469_/X vssd1 vssd1 vccd1 vccd1 _21161_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13211_ input51/X vssd1 vssd1 vccd1 vccd1 _13211_/X sky130_fd_sc_hd__clkbuf_2
X_10423_ _20675_/Q vssd1 vssd1 vccd1 vccd1 _10423_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13559__A _13566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14191_ _14191_/A vssd1 vssd1 vccd1 vccd1 _14191_/X sky130_fd_sc_hd__buf_1
XFILLER_152_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11574__A1 _21127_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20126__CLK _21452_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13142_ _13167_/A vssd1 vssd1 vccd1 vccd1 _13142_/X sky130_fd_sc_hd__buf_1
XANTENNA_input63_A HWDATA[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10354_ _10266_/A _20709_/Q _10275_/A _20719_/Q _10353_/X vssd1 vssd1 vccd1 vccd1
+ _10360_/C sky130_fd_sc_hd__o221a_1
XANTENNA__17973__B _17973_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17950_ _18517_/X _17907_/X _18531_/X _17908_/X vssd1 vssd1 vccd1 vccd1 _17957_/B
+ sky130_fd_sc_hd__a22o_1
X_13073_ _13073_/A vssd1 vssd1 vccd1 vccd1 _13073_/X sky130_fd_sc_hd__buf_1
XANTENNA__21184__RESET_B repeater220/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10285_ _10285_/A _10285_/B vssd1 vssd1 vccd1 vccd1 _10372_/A sky130_fd_sc_hd__or2_1
X_12024_ _12030_/A vssd1 vssd1 vccd1 vccd1 _12024_/X sky130_fd_sc_hd__buf_1
XFILLER_151_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16901_ _16901_/A vssd1 vssd1 vccd1 vccd1 _16906_/B sky130_fd_sc_hd__inv_2
XFILLER_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17881_ _18483_/X _17839_/X _18474_/X _17840_/X vssd1 vssd1 vccd1 vccd1 _17881_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__21113__RESET_B repeater233/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19620_ _21452_/CLK _19620_/D vssd1 vssd1 vccd1 vccd1 _19620_/Q sky130_fd_sc_hd__dfxtp_1
X_16832_ _16829_/Y _16830_/Y _16831_/X vssd1 vssd1 vccd1 vccd1 _16832_/X sky130_fd_sc_hd__o21a_1
XFILLER_93_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11526__B _14273_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19551_ _19706_/CLK _19551_/D vssd1 vssd1 vccd1 vccd1 _19551_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_207_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16763_ _16766_/B _16761_/X _16762_/X vssd1 vssd1 vccd1 vccd1 _16763_/X sky130_fd_sc_hd__o21a_1
XFILLER_93_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18296__S _18884_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13975_ _20563_/Q _13990_/A vssd1 vssd1 vccd1 vccd1 _13976_/D sky130_fd_sc_hd__or2_1
X_18502_ _18845_/A0 _10517_/Y _18896_/S vssd1 vssd1 vccd1 vccd1 _18502_/X sky130_fd_sc_hd__mux2_1
XFILLER_202_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15714_ _19667_/Q _15709_/X _15663_/X _15711_/X vssd1 vssd1 vccd1 vccd1 _19667_/D
+ sky130_fd_sc_hd__a22o_1
X_19482_ _19626_/CLK _19482_/D vssd1 vssd1 vccd1 vccd1 _19482_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12926_ _12926_/A vssd1 vssd1 vccd1 vccd1 _12926_/X sky130_fd_sc_hd__buf_1
X_16694_ _16700_/A _18945_/X vssd1 vssd1 vccd1 vccd1 _19891_/D sky130_fd_sc_hd__and2_1
XFILLER_207_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18433_ _18432_/X _20579_/Q _18907_/S vssd1 vssd1 vccd1 vccd1 _18433_/X sky130_fd_sc_hd__mux2_2
XFILLER_222_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15645_ _19699_/Q _15640_/X _15475_/X _15642_/X vssd1 vssd1 vccd1 vccd1 _19699_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12857_ _12857_/A vssd1 vssd1 vccd1 vccd1 _12857_/X sky130_fd_sc_hd__buf_2
XPHY_4081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18364_ _18034_/Y _20762_/Q _18891_/S vssd1 vssd1 vccd1 vccd1 _18364_/X sky130_fd_sc_hd__mux2_1
X_11808_ _11848_/A _11848_/B vssd1 vssd1 vccd1 vccd1 _11845_/B sky130_fd_sc_hd__nand2_1
X_15576_ _15584_/A vssd1 vssd1 vccd1 vccd1 _15576_/X sky130_fd_sc_hd__buf_1
X_12788_ _20787_/Q _12784_/X _09645_/X _12786_/X vssd1 vssd1 vccd1 vccd1 _20787_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_57_HCLK clkbuf_4_14_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _21319_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17315_ _17315_/A vssd1 vssd1 vccd1 vccd1 _17315_/X sky130_fd_sc_hd__clkbuf_2
X_11739_ _11739_/A vssd1 vssd1 vccd1 vccd1 _11739_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__15949__A _16340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14527_ _17169_/A _17169_/B _16479_/A _17320_/A vssd1 vssd1 vccd1 vccd1 _16484_/A
+ sky130_fd_sc_hd__or4_4
X_18295_ _18009_/Y _16978_/Y _18680_/S vssd1 vssd1 vccd1 vccd1 _18295_/X sky130_fd_sc_hd__mux2_2
XPHY_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17246_ _19503_/Q vssd1 vssd1 vccd1 vccd1 _17246_/Y sky130_fd_sc_hd__inv_2
X_14458_ _14477_/A vssd1 vssd1 vccd1 vccd1 _14458_/X sky130_fd_sc_hd__buf_1
XFILLER_30_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13409_ _20485_/Q _13404_/X _13213_/X _13405_/X vssd1 vssd1 vccd1 vccd1 _20485_/D
+ sky130_fd_sc_hd__a22o_1
X_14389_ _14328_/A _20027_/Q _21467_/Q _14498_/A vssd1 vssd1 vccd1 vccd1 _14394_/B
+ sky130_fd_sc_hd__a22o_1
X_17177_ _17177_/A _17177_/B vssd1 vssd1 vccd1 vccd1 _18901_/S sky130_fd_sc_hd__nor2_8
XFILLER_183_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12762__B1 _12656_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16128_ _19470_/Q _16119_/X _16127_/X _16121_/X vssd1 vssd1 vccd1 vccd1 _19470_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_115_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16059_ _19504_/Q _16056_/X _15772_/X _16057_/X vssd1 vssd1 vccd1 vccd1 _19504_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_143_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09682__A _12550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19818_ _19820_/CLK _19818_/D vssd1 vssd1 vccd1 vccd1 _19818_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__19931__RESET_B repeater251/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19749_ _19811_/CLK _19749_/D vssd1 vssd1 vccd1 vccd1 _19749_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_244_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20836__RESET_B repeater257/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15216__C1 _15160_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_240_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18934__S _18946_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12548__A _12548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20524_ _20944_/CLK _20524_/D repeater274/X vssd1 vssd1 vccd1 vccd1 _20524_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_165_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20455_ _20476_/CLK _20455_/D repeater280/X vssd1 vssd1 vccd1 vccd1 _20455_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_107_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20386_ _20971_/CLK _20386_/D repeater280/X vssd1 vssd1 vccd1 vccd1 _20386_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_88_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10070_ _21398_/Q vssd1 vssd1 vccd1 vccd1 _10071_/A sky130_fd_sc_hd__inv_2
XFILLER_130_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21007_ _21011_/CLK _21007_/D repeater235/X vssd1 vssd1 vccd1 vccd1 _21007_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_75_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_236_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19005__S _19019_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13760_ _13755_/Y _20183_/Q _20604_/Q _14571_/A _13759_/X vssd1 vssd1 vccd1 vccd1
+ _13761_/D sky130_fd_sc_hd__o221a_1
XFILLER_62_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10972_ _12742_/A _12735_/A _11964_/A vssd1 vssd1 vccd1 vccd1 _16594_/A sky130_fd_sc_hd__or3_4
XFILLER_46_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12711_ _20812_/Q _12707_/X _11741_/X _12708_/X vssd1 vssd1 vccd1 vccd1 _20812_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_231_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13691_ _20345_/Q _13686_/X _12855_/A _13688_/X vssd1 vssd1 vccd1 vccd1 _20345_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18844__S _18898_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12642_ input12/X _12637_/X _20844_/Q _12638_/X vssd1 vssd1 vccd1 vccd1 _20844_/D
+ sky130_fd_sc_hd__o22a_1
XPHY_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15430_ _19799_/Q _15423_/X _15429_/X _15425_/X vssd1 vssd1 vccd1 vccd1 _19799_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_70_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15361_ _15367_/A vssd1 vssd1 vccd1 vccd1 _15361_/X sky130_fd_sc_hd__buf_1
XFILLER_200_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12573_ _10859_/B _12566_/X _18241_/X _18242_/S vssd1 vssd1 vccd1 vccd1 _20889_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17100_ _19406_/Q vssd1 vssd1 vccd1 vccd1 _17100_/Y sky130_fd_sc_hd__inv_2
X_11524_ _17290_/A vssd1 vssd1 vccd1 vccd1 _11678_/A sky130_fd_sc_hd__buf_1
XFILLER_157_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12992__B1 _12991_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14312_ _14275_/Y _14302_/X _14290_/Y _14311_/X vssd1 vssd1 vccd1 vccd1 _20242_/D
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15292_ _19858_/Q _15292_/B vssd1 vssd1 vccd1 vccd1 _15293_/B sky130_fd_sc_hd__or2_1
XFILLER_12_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18080_ _18080_/A _18083_/B vssd1 vssd1 vccd1 vccd1 _18080_/Y sky130_fd_sc_hd__nor2_1
XFILLER_129_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14243_ _19903_/Q _14243_/B vssd1 vssd1 vccd1 vccd1 _14246_/A sky130_fd_sc_hd__or2_4
X_17031_ _17031_/A vssd1 vssd1 vccd1 vccd1 _17035_/B sky130_fd_sc_hd__buf_1
XFILLER_144_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_148_HCLK_A clkbuf_opt_1_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11455_ _21043_/Q vssd1 vssd1 vccd1 vccd1 _11457_/A sky130_fd_sc_hd__inv_2
XFILLER_172_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15930__B1 _15791_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__21365__RESET_B repeater254/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10406_ _10406_/A vssd1 vssd1 vccd1 vccd1 _10406_/Y sky130_fd_sc_hd__inv_2
X_14174_ _14191_/A vssd1 vssd1 vccd1 vccd1 _14174_/X sky130_fd_sc_hd__clkbuf_2
X_11386_ _11388_/B _11386_/B _11388_/A vssd1 vssd1 vccd1 vccd1 _11389_/A sky130_fd_sc_hd__nor3b_4
X_13125_ _20623_/Q _13120_/X _13003_/X _13121_/X vssd1 vssd1 vccd1 vccd1 _20623_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_98_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10337_ _20725_/Q vssd1 vssd1 vccd1 vccd1 _18006_/A sky130_fd_sc_hd__inv_2
X_18982_ _21424_/Q _21097_/Q _18983_/S vssd1 vssd1 vccd1 vccd1 _18982_/X sky130_fd_sc_hd__mux2_1
XFILLER_152_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17933_ _17933_/A vssd1 vssd1 vccd1 vccd1 _17947_/A sky130_fd_sc_hd__clkbuf_2
X_13056_ _20665_/Q _13052_/X _12984_/X _13055_/X vssd1 vssd1 vccd1 vccd1 _20665_/D
+ sky130_fd_sc_hd__a22o_1
X_10268_ _10268_/A _10268_/B vssd1 vssd1 vccd1 vccd1 _10406_/A sky130_fd_sc_hd__or2_2
XFILLER_238_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12007_ _20998_/Q _12003_/X _20251_/Q _12006_/X vssd1 vssd1 vccd1 vccd1 _19908_/D
+ sky130_fd_sc_hd__o211ai_4
XFILLER_94_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17864_ _18546_/X _17861_/X _18584_/X _17862_/X _17863_/X vssd1 vssd1 vccd1 vccd1
+ _17864_/X sky130_fd_sc_hd__o221a_2
XFILLER_238_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10199_ _10199_/A vssd1 vssd1 vccd1 vccd1 _10221_/A sky130_fd_sc_hd__buf_1
XFILLER_213_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19603_ _20142_/CLK _19603_/D vssd1 vssd1 vccd1 vccd1 _19603_/Q sky130_fd_sc_hd__dfxtp_1
X_16815_ _16815_/A _16815_/B vssd1 vssd1 vccd1 vccd1 _16815_/Y sky130_fd_sc_hd__nor2_1
X_17795_ _17793_/Y _17141_/A _17794_/Y _17295_/X vssd1 vssd1 vccd1 vccd1 _17795_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__15997__B1 _15949_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14848__A _20497_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19534_ _19784_/CLK _19534_/D vssd1 vssd1 vccd1 vccd1 _19534_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16746_ _16848_/A vssd1 vssd1 vccd1 vccd1 _16835_/A sky130_fd_sc_hd__inv_2
XANTENNA__19283__S0 _19285_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13958_ _20657_/Q vssd1 vssd1 vccd1 vccd1 _13958_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19465_ _20137_/CLK _19465_/D vssd1 vssd1 vccd1 vccd1 _19465_/Q sky130_fd_sc_hd__dfxtp_1
X_12909_ _12924_/A vssd1 vssd1 vccd1 vccd1 _12909_/X sky130_fd_sc_hd__buf_1
X_16677_ _21165_/Q _11453_/B _11454_/B vssd1 vssd1 vccd1 vccd1 _16677_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__18754__S _18910_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13889_ _13974_/B _13889_/B vssd1 vssd1 vccd1 vccd1 _13986_/A sky130_fd_sc_hd__or2_1
X_18416_ _17830_/X _09725_/Y _18928_/S vssd1 vssd1 vccd1 vccd1 _18416_/X sky130_fd_sc_hd__mux2_1
X_15628_ _19709_/Q _15625_/X _15544_/X _15627_/X vssd1 vssd1 vccd1 vccd1 _19709_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_222_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19396_ _21001_/CLK _19396_/D vssd1 vssd1 vccd1 vccd1 _19396_/Q sky130_fd_sc_hd__dfxtp_1
X_18347_ _18346_/X _12229_/Y _18910_/S vssd1 vssd1 vccd1 vccd1 _18347_/X sky130_fd_sc_hd__mux2_1
XFILLER_159_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15559_ _15559_/A vssd1 vssd1 vccd1 vccd1 _15778_/B sky130_fd_sc_hd__buf_1
XFILLER_159_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18278_ _19181_/X _21273_/Q _18281_/S vssd1 vssd1 vccd1 vccd1 _18278_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12815__B _13108_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput40 HWDATA[11] vssd1 vssd1 vccd1 vccd1 input40/X sky130_fd_sc_hd__clkbuf_2
X_17229_ _17732_/A vssd1 vssd1 vccd1 vccd1 _18019_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_238_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19112__A0 _17046_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11538__A1 _21137_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput51 HWDATA[21] vssd1 vssd1 vccd1 vccd1 input51/X sky130_fd_sc_hd__buf_2
Xinput62 HWDATA[31] vssd1 vssd1 vccd1 vccd1 input62/X sky130_fd_sc_hd__buf_4
Xinput73 RsRx_S0 vssd1 vssd1 vccd1 vccd1 input73/X sky130_fd_sc_hd__clkbuf_4
XFILLER_128_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20240_ _21481_/CLK _20240_/D repeater206/X vssd1 vssd1 vccd1 vccd1 _20240_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__21035__RESET_B repeater242/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09982_ _21412_/Q _09975_/A _09702_/X _09976_/A vssd1 vssd1 vccd1 vccd1 _21412_/D
+ sky130_fd_sc_hd__a22o_1
X_20171_ _21125_/CLK _20171_/D repeater190/X vssd1 vssd1 vccd1 vccd1 _20171_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__20591__CLK _20592_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18929__S _18929_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13160__B1 _12950_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20670__RESET_B repeater211/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13662__A _13680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09667__B1 _09666_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19274__S0 _19275_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18664__S _18907_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_9_HCLK clkbuf_opt_2_HCLK/A vssd1 vssd1 vccd1 vccd1 _20327_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_40_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20507_ _20929_/CLK _20507_/D repeater266/X vssd1 vssd1 vccd1 vccd1 _20507_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_138_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11240_ _21195_/Q _11239_/X _19910_/Q _11235_/Y vssd1 vssd1 vccd1 vccd1 _21195_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_180_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20438_ _20470_/CLK _20438_/D repeater279/X vssd1 vssd1 vccd1 vccd1 _20438_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_106_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11171_ _21221_/Q vssd1 vssd1 vccd1 vccd1 _16465_/B sky130_fd_sc_hd__inv_2
X_20369_ _20957_/CLK _20369_/D repeater187/X vssd1 vssd1 vccd1 vccd1 _20369_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_164_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10122_ _10114_/X _10122_/B _10122_/C _10122_/D vssd1 vssd1 vccd1 vccd1 _10137_/C
+ sky130_fd_sc_hd__and4b_1
XFILLER_121_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18839__S _18884_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14930_ _20577_/Q vssd1 vssd1 vccd1 vccd1 _14930_/Y sky130_fd_sc_hd__inv_2
X_10053_ _10201_/A _10200_/C _10053_/C _10053_/D vssd1 vssd1 vccd1 vccd1 _10148_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_208_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input26_A HADDR[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14861_ _20087_/Q vssd1 vssd1 vccd1 vccd1 _14863_/C sky130_fd_sc_hd__inv_2
XFILLER_208_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16600_ _19989_/Q vssd1 vssd1 vccd1 vccd1 _16600_/Y sky130_fd_sc_hd__inv_2
XFILLER_180_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13812_ _20180_/Q vssd1 vssd1 vccd1 vccd1 _14570_/A sky130_fd_sc_hd__inv_2
Xclkbuf_4_3_0_HCLK clkbuf_4_3_0_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_3_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_17580_ _17889_/A vssd1 vssd1 vccd1 vccd1 _17823_/A sky130_fd_sc_hd__inv_2
XFILLER_29_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14792_ _14792_/A _16481_/B vssd1 vssd1 vccd1 vccd1 _16480_/A sky130_fd_sc_hd__or2_1
XANTENNA__19265__S0 _19275_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16531_ _16681_/B _16530_/Y _19997_/Q _16521_/B _16632_/B vssd1 vssd1 vccd1 vccd1
+ _19997_/D sky130_fd_sc_hd__a221o_1
XFILLER_216_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13743_ _20194_/Q vssd1 vssd1 vccd1 vccd1 _14583_/A sky130_fd_sc_hd__inv_2
X_10955_ _10951_/Y _21030_/Q _21203_/Q _11807_/A _10954_/X vssd1 vssd1 vccd1 vccd1
+ _10969_/B sky130_fd_sc_hd__o221a_1
XANTENNA__18574__S _18902_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19250_ _17362_/Y _17363_/Y _17364_/Y _17365_/Y _20130_/Q _20131_/Q vssd1 vssd1 vccd1
+ vccd1 _19250_/X sky130_fd_sc_hd__mux4_2
X_16462_ _19302_/Q _16459_/X _16338_/X _16460_/X vssd1 vssd1 vccd1 vccd1 _19302_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_73_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13674_ _13680_/A vssd1 vssd1 vccd1 vccd1 _13674_/X sky130_fd_sc_hd__buf_1
X_10886_ _12548_/A vssd1 vssd1 vccd1 vccd1 _10886_/X sky130_fd_sc_hd__buf_2
X_18201_ _18200_/X _16957_/Y _18680_/S vssd1 vssd1 vccd1 vccd1 _18201_/X sky130_fd_sc_hd__mux2_2
XFILLER_92_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11217__B1 _09663_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15413_ _15413_/A _15505_/B _16594_/B vssd1 vssd1 vccd1 vccd1 _15778_/C sky130_fd_sc_hd__or3_4
XPHY_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19181_ _19177_/X _19178_/X _19179_/X _19180_/X _20123_/Q _20124_/Q vssd1 vssd1 vccd1
+ vccd1 _19181_/X sky130_fd_sc_hd__mux4_2
X_12625_ _12637_/A vssd1 vssd1 vccd1 vccd1 _12625_/X sky130_fd_sc_hd__buf_1
XPHY_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16393_ _16399_/A vssd1 vssd1 vccd1 vccd1 _16400_/A sky130_fd_sc_hd__inv_2
XPHY_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_repeater165_A _18874_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18132_ _18131_/X _18052_/Y _18669_/S vssd1 vssd1 vccd1 vccd1 _18132_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12965__B1 _12884_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12556_ _20895_/Q _12553_/X _11739_/X _12554_/X vssd1 vssd1 vccd1 vccd1 _20895_/D
+ sky130_fd_sc_hd__a22o_1
X_15344_ _19834_/Q _15337_/X _15343_/X _15339_/X vssd1 vssd1 vccd1 vccd1 _19834_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_157_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11507_ _20251_/Q vssd1 vssd1 vccd1 vccd1 _16711_/A sky130_fd_sc_hd__buf_1
XFILLER_129_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18063_ _18274_/X _18019_/X _18127_/X _18020_/X _18062_/X vssd1 vssd1 vccd1 vccd1
+ _18068_/B sky130_fd_sc_hd__o221a_2
XANTENNA__10436__A _20695_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15275_ _20485_/Q _15112_/X _20476_/Q _15069_/A _15274_/X vssd1 vssd1 vccd1 vccd1
+ _15284_/B sky130_fd_sc_hd__o221a_1
X_12487_ _20923_/Q _12486_/Y _12472_/B _12480_/X vssd1 vssd1 vccd1 vccd1 _20923_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_7_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17014_ _19981_/Q vssd1 vssd1 vccd1 vccd1 _17014_/Y sky130_fd_sc_hd__inv_2
X_11438_ _11437_/Y _11408_/X _11413_/X _11384_/B _11414_/X vssd1 vssd1 vccd1 vccd1
+ _11439_/A sky130_fd_sc_hd__o32a_1
XFILLER_144_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output94_A _18027_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14226_ _20262_/Q _14225_/Y _14191_/A _14074_/B vssd1 vssd1 vccd1 vccd1 _20262_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_99_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14157_ _20542_/Q _14081_/A _20550_/Q _14089_/A vssd1 vssd1 vccd1 vccd1 _14157_/X
+ sky130_fd_sc_hd__o22a_1
X_11369_ _21175_/Q vssd1 vssd1 vccd1 vccd1 _11387_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_99_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12651__A input62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13108_ _13108_/A _13108_/B vssd1 vssd1 vccd1 vccd1 _13109_/S sky130_fd_sc_hd__or2_1
X_18965_ _16617_/X _16617_/A _18976_/S vssd1 vssd1 vccd1 vccd1 _18965_/X sky130_fd_sc_hd__mux2_1
X_14088_ _14088_/A _14198_/A vssd1 vssd1 vccd1 vccd1 _14089_/B sky130_fd_sc_hd__or2_2
XANTENNA__18749__S _18849_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20499__RESET_B repeater267/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13039_ _20670_/Q _13034_/X _12872_/X _13035_/X vssd1 vssd1 vccd1 vccd1 _20670_/D
+ sky130_fd_sc_hd__a22o_1
X_17916_ _18418_/X _17200_/X _18471_/X _17224_/X _17915_/X vssd1 vssd1 vccd1 vccd1
+ _17916_/X sky130_fd_sc_hd__o221a_1
XFILLER_239_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18896_ _18895_/X _13800_/Y _18896_/S vssd1 vssd1 vccd1 vccd1 _18896_/X sky130_fd_sc_hd__mux2_1
XFILLER_239_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17847_ _17833_/X _17852_/A _17838_/X _17843_/X _17846_/X vssd1 vssd1 vccd1 vccd1
+ _17847_/Y sky130_fd_sc_hd__o2111ai_4
XFILLER_208_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13482__A input48/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17778_ _20818_/Q vssd1 vssd1 vccd1 vccd1 _17778_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19256__S0 _21005_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_241_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19517_ _21462_/CLK _19517_/D vssd1 vssd1 vccd1 vccd1 _19517_/Q sky130_fd_sc_hd__dfxtp_1
X_16729_ _20991_/Q _11997_/B _11998_/B vssd1 vssd1 vccd1 vccd1 _16729_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__18484__S _18908_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_241_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20010__RESET_B repeater238/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_234_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19448_ _21234_/CLK _19448_/D vssd1 vssd1 vccd1 vccd1 _19448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16395__B1 _16231_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19379_ _19812_/CLK _19379_/D vssd1 vssd1 vccd1 vccd1 _19379_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__21287__RESET_B repeater207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21410_ _21417_/CLK _21410_/D repeater231/X vssd1 vssd1 vccd1 vccd1 _21410_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_194_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__21216__RESET_B repeater238/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21341_ _21341_/CLK _21341_/D repeater201/X vssd1 vssd1 vccd1 vccd1 _21341_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_163_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_131_HCLK_A clkbuf_4_4_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21272_ _21273_/CLK _21272_/D repeater245/X vssd1 vssd1 vccd1 vccd1 _21272_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_162_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20223_ _21484_/CLK _20223_/D repeater202/X vssd1 vssd1 vccd1 vccd1 _20223_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_144_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13657__A _13657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13381__B1 _13171_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20154_ _21242_/CLK _20154_/D repeater189/X vssd1 vssd1 vccd1 vccd1 _20154_/Q sky130_fd_sc_hd__dfrtp_1
X_09965_ _12725_/B vssd1 vssd1 vccd1 vccd1 _12605_/A sky130_fd_sc_hd__buf_2
XANTENNA__18659__S _18874_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20851__RESET_B repeater243/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20085_ _20496_/CLK _20085_/D repeater274/X vssd1 vssd1 vccd1 vccd1 _20085_/Q sky130_fd_sc_hd__dfrtp_1
X_09896_ _20010_/Q _09912_/A _09884_/A vssd1 vssd1 vccd1 vccd1 _17024_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__20169__RESET_B repeater190/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19247__S0 _20130_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20987_ _21319_/CLK _20987_/D repeater191/X vssd1 vssd1 vccd1 vccd1 _20987_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_25_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18394__S _18849_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10740_ _19928_/Q _16786_/A vssd1 vssd1 vccd1 vccd1 _16790_/A sky130_fd_sc_hd__or2_1
XFILLER_214_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10671_ _21338_/Q _10669_/X _10670_/X _10666_/A vssd1 vssd1 vccd1 vccd1 _21338_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_40_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12410_ _12410_/A vssd1 vssd1 vccd1 vccd1 _12462_/A sky130_fd_sc_hd__buf_1
XANTENNA__12947__B1 _12699_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_11_0_HCLK clkbuf_3_5_0_HCLK/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_11_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_13390_ _13410_/A vssd1 vssd1 vccd1 vccd1 _13390_/X sky130_fd_sc_hd__buf_1
XFILLER_223_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12341_ _12331_/A _12331_/B _12376_/A _12339_/Y vssd1 vssd1 vccd1 vccd1 _20978_/D
+ sky130_fd_sc_hd__a211oi_4
XFILLER_194_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15060_ _15060_/A _15214_/A vssd1 vssd1 vccd1 vccd1 _15061_/B sky130_fd_sc_hd__or2_2
XFILLER_4_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12272_ _12470_/A _20502_/Q _20944_/Q _12268_/Y _12271_/X vssd1 vssd1 vccd1 vccd1
+ _12278_/C sky130_fd_sc_hd__o221a_1
XFILLER_126_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14011_ _14011_/A _14028_/A vssd1 vssd1 vccd1 vccd1 _14026_/A sky130_fd_sc_hd__or2_2
XANTENNA__13567__A _13567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20939__RESET_B repeater278/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11223_ _21202_/Q _11219_/X _10889_/X _11220_/X vssd1 vssd1 vccd1 vccd1 _21202_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17039__A _21410_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_53_HCLK_A clkbuf_4_9_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11154_ _20891_/Q _17169_/B _16479_/A _17315_/A vssd1 vssd1 vccd1 vccd1 _16616_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_1_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17981__B _18001_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18569__S _18891_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13124__B1 _13001_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20592__RESET_B repeater259/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10105_ _10206_/A _20782_/Q _21385_/Q _10103_/Y _10104_/X vssd1 vssd1 vccd1 vccd1
+ _10112_/B sky130_fd_sc_hd__o221a_1
XFILLER_150_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18750_ _18749_/X _20263_/Q _18850_/S vssd1 vssd1 vccd1 vccd1 _18750_/X sky130_fd_sc_hd__mux2_2
X_11085_ _11085_/A vssd1 vssd1 vccd1 vccd1 _11086_/B sky130_fd_sc_hd__inv_2
X_15962_ _15962_/A vssd1 vssd1 vccd1 vccd1 _15962_/X sky130_fd_sc_hd__buf_1
XFILLER_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17701_ _19468_/Q vssd1 vssd1 vccd1 vccd1 _17701_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14913_ _14909_/Y _20078_/Q _14910_/Y _20103_/Q _14912_/X vssd1 vssd1 vccd1 vccd1
+ _14918_/C sky130_fd_sc_hd__o221a_1
X_10036_ _21380_/Q vssd1 vssd1 vccd1 vccd1 _10201_/A sky130_fd_sc_hd__inv_2
X_18681_ _18845_/A0 _17709_/Y _18879_/S vssd1 vssd1 vccd1 vccd1 _18681_/X sky130_fd_sc_hd__mux2_1
XANTENNA_output132_A _21248_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15893_ _16237_/A vssd1 vssd1 vccd1 vccd1 _15893_/X sky130_fd_sc_hd__clkbuf_2
X_17632_ _18736_/X _17703_/B vssd1 vssd1 vccd1 vccd1 _17632_/Y sky130_fd_sc_hd__nand2_1
X_14844_ _20090_/Q vssd1 vssd1 vccd1 vccd1 _14845_/A sky130_fd_sc_hd__inv_2
XFILLER_91_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19238__S0 _20130_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17563_ _21131_/Q vssd1 vssd1 vccd1 vccd1 _17563_/Y sky130_fd_sc_hd__inv_2
X_14775_ _14775_/A vssd1 vssd1 vccd1 vccd1 _14779_/A sky130_fd_sc_hd__buf_1
XFILLER_223_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11987_ _11983_/X _11985_/X _11883_/X _11986_/Y _19118_/X vssd1 vssd1 vccd1 vccd1
+ _11988_/A sky130_fd_sc_hd__o32a_1
XFILLER_216_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19302_ _20172_/CLK _19302_/D vssd1 vssd1 vccd1 vccd1 _19302_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16514_ _16688_/A _16510_/Y _16511_/Y _16494_/X _16513_/Y vssd1 vssd1 vccd1 vccd1
+ _20000_/D sky130_fd_sc_hd__o221ai_1
X_13726_ _20327_/Q vssd1 vssd1 vccd1 vccd1 _15769_/A sky130_fd_sc_hd__clkbuf_2
X_10938_ _21197_/Q _11864_/A _10933_/Y _10934_/X _10937_/X vssd1 vssd1 vccd1 vccd1
+ _10970_/B sky130_fd_sc_hd__o221a_1
X_17494_ _19506_/Q vssd1 vssd1 vccd1 vccd1 _17494_/Y sky130_fd_sc_hd__inv_2
X_19233_ _17488_/Y _17489_/Y _17490_/Y _17491_/Y _19275_/S0 _21004_/Q vssd1 vssd1
+ vccd1 vccd1 _19233_/X sky130_fd_sc_hd__mux4_2
XFILLER_231_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16445_ _19310_/Q _16441_/X _16340_/X _16442_/X vssd1 vssd1 vccd1 vccd1 _19310_/D
+ sky130_fd_sc_hd__a22o_1
X_10869_ _21265_/Q _10864_/X _09682_/X _10866_/X vssd1 vssd1 vccd1 vccd1 _21265_/D
+ sky130_fd_sc_hd__a22o_1
X_13657_ _13657_/A _13657_/B vssd1 vssd1 vccd1 vccd1 _13685_/A sky130_fd_sc_hd__or2_2
XANTENNA__09939__B _17231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12938__B1 _12849_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12608_ _20868_/Q _12574_/A _18220_/X _12575_/A vssd1 vssd1 vccd1 vccd1 _20868_/D
+ sky130_fd_sc_hd__a22o_1
X_19164_ _19726_/Q _19366_/Q _19782_/Q _19766_/Q _19280_/S0 _20122_/Q vssd1 vssd1
+ vccd1 vccd1 _19164_/X sky130_fd_sc_hd__mux4_2
XPHY_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16376_ _19349_/Q _16370_/X _16375_/X _16371_/X vssd1 vssd1 vccd1 vccd1 _19349_/D
+ sky130_fd_sc_hd__a22o_1
X_13588_ _13594_/A vssd1 vssd1 vccd1 vccd1 _13588_/X sky130_fd_sc_hd__buf_1
XFILLER_12_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18115_ _21486_/Q _15329_/X _13560_/X _15330_/X vssd1 vssd1 vccd1 vccd1 _21486_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_200_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15327_ _20029_/Q _15323_/X _13547_/X _15324_/X vssd1 vssd1 vccd1 vccd1 _20029_/D
+ sky130_fd_sc_hd__a22o_1
X_12539_ _11306_/B _12518_/A _11312_/A _12521_/A vssd1 vssd1 vccd1 vccd1 _20903_/D
+ sky130_fd_sc_hd__a22o_1
X_19095_ _16675_/X _21083_/Q _19870_/D vssd1 vssd1 vccd1 vccd1 _19095_/X sky130_fd_sc_hd__mux2_1
XFILLER_219_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18046_ _18331_/X _18021_/X _18314_/X _18045_/X vssd1 vssd1 vccd1 vccd1 _18046_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_145_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15258_ _20466_/Q _15060_/A _15257_/Y _15092_/X vssd1 vssd1 vccd1 vccd1 _15258_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_144_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13363__B1 _13146_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13477__A input51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14209_ _14209_/A vssd1 vssd1 vccd1 vccd1 _14209_/Y sky130_fd_sc_hd__inv_2
XFILLER_132_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15189_ _20061_/Q _15188_/Y _15076_/B _15177_/X vssd1 vssd1 vccd1 vccd1 _20061_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_98_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19997_ _21055_/CLK _19997_/D repeater220/X vssd1 vssd1 vccd1 vccd1 _19997_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_140_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18479__S _18903_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09750_ _21227_/Q vssd1 vssd1 vccd1 vccd1 _11052_/D sky130_fd_sc_hd__inv_2
X_18948_ _21051_/Q _21088_/Q _19843_/Q vssd1 vssd1 vccd1 vccd1 _18948_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20262__RESET_B repeater264/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09690__A _15329_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09681_ _15385_/A vssd1 vssd1 vccd1 vccd1 _12550_/A sky130_fd_sc_hd__clkbuf_4
X_18879_ _18878_/X _17188_/Y _18879_/S vssd1 vssd1 vccd1 vccd1 _18879_/X sky130_fd_sc_hd__mux2_1
X_20910_ _21196_/CLK _20910_/D repeater218/X vssd1 vssd1 vccd1 vccd1 _20910_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__17801__B1 _18673_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_215_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19229__S0 _20130_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_243_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20841_ _20841_/CLK _20841_/D repeater256/X vssd1 vssd1 vccd1 vccd1 _20841_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21468__RESET_B repeater204/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19103__S _19870_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20772_ _21406_/CLK _20772_/D repeater213/X vssd1 vssd1 vccd1 vccd1 _20772_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18942__S _18946_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12929__B1 _12928_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11601__B1 _21120_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21324_ _21341_/CLK _21324_/D repeater204/X vssd1 vssd1 vccd1 vccd1 _21324_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_191_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12157__A1 _12036_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13354__B1 _13219_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21255_ _21255_/CLK _21255_/D repeater240/X vssd1 vssd1 vccd1 vccd1 _21255_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_116_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20206_ _20623_/CLK _20206_/D repeater194/X vssd1 vssd1 vccd1 vccd1 _20206_/Q sky130_fd_sc_hd__dfrtp_1
X_21186_ _21193_/CLK _21186_/D repeater224/X vssd1 vssd1 vccd1 vccd1 _21186_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18389__S _18907_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20137_ _20137_/CLK _20137_/D repeater248/X vssd1 vssd1 vccd1 vccd1 _20137_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_132_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09948_ _10877_/A _17060_/A _12725_/B vssd1 vssd1 vccd1 vccd1 _13384_/C sky130_fd_sc_hd__or3_4
XFILLER_219_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20068_ _20070_/CLK _20068_/D repeater276/X vssd1 vssd1 vccd1 vccd1 _20068_/Q sky130_fd_sc_hd__dfrtp_1
X_09879_ _21440_/Q _21439_/Q _09870_/A vssd1 vssd1 vccd1 vccd1 _09879_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_38_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11910_ _11913_/A _11910_/B vssd1 vssd1 vccd1 vccd1 _11910_/X sky130_fd_sc_hd__or2_1
XFILLER_245_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12890_ input38/X vssd1 vssd1 vccd1 vccd1 _13600_/A sky130_fd_sc_hd__buf_2
XPHY_4411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11841_ _11841_/A vssd1 vssd1 vccd1 vccd1 _11842_/B sky130_fd_sc_hd__inv_2
XPHY_4444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19013__S _19019_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11772_ _19087_/X _11770_/X _21047_/Q _11771_/X vssd1 vssd1 vccd1 vccd1 _21047_/D
+ sky130_fd_sc_hd__a22o_1
X_14560_ _16077_/A vssd1 vssd1 vccd1 vccd1 _15816_/A sky130_fd_sc_hd__buf_1
XPHY_4488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10723_ _10723_/A _10723_/B _10723_/C vssd1 vssd1 vccd1 vccd1 _10726_/A sky130_fd_sc_hd__or3_4
X_13511_ _14264_/A vssd1 vssd1 vccd1 vccd1 _13511_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_213_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14491_ _20224_/Q _14490_/Y _14368_/B _14477_/X vssd1 vssd1 vccd1 vccd1 _20224_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__18852__S _18906_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16230_ _16240_/A vssd1 vssd1 vccd1 vccd1 _16230_/X sky130_fd_sc_hd__buf_1
X_10654_ _10654_/A _10693_/A vssd1 vssd1 vccd1 vccd1 _10655_/B sky130_fd_sc_hd__or2_2
X_13442_ _15421_/A vssd1 vssd1 vccd1 vccd1 _13442_/X sky130_fd_sc_hd__buf_2
XANTENNA__17976__B _17978_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_90_HCLK clkbuf_4_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20724_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__13593__B1 _13442_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16161_ _19456_/Q _16158_/X _16145_/X _16159_/X vssd1 vssd1 vccd1 vccd1 _19456_/D
+ sky130_fd_sc_hd__a22o_1
X_13373_ _20505_/Q _13371_/X _13240_/X _13372_/X vssd1 vssd1 vccd1 vccd1 _20505_/D
+ sky130_fd_sc_hd__a22o_1
X_10585_ _20743_/Q vssd1 vssd1 vccd1 vccd1 _10585_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15112_ _15112_/A vssd1 vssd1 vccd1 vccd1 _15112_/X sky130_fd_sc_hd__clkbuf_2
X_12324_ _12324_/A _12355_/A vssd1 vssd1 vccd1 vccd1 _12325_/B sky130_fd_sc_hd__or2_1
X_16092_ _19486_/Q _16087_/X _15916_/X _16088_/X vssd1 vssd1 vccd1 vccd1 _19486_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_181_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12148__B2 _20344_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19920_ _21379_/CLK _19920_/D repeater212/X vssd1 vssd1 vccd1 vccd1 _19920_/Q sky130_fd_sc_hd__dfrtp_1
X_15043_ _20059_/Q vssd1 vssd1 vccd1 vccd1 _15073_/A sky130_fd_sc_hd__inv_2
X_12255_ _12255_/A _12255_/B _12255_/C _12255_/D vssd1 vssd1 vccd1 vccd1 _12302_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_126_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11206_ _11225_/A vssd1 vssd1 vccd1 vccd1 _11206_/X sky130_fd_sc_hd__buf_1
XANTENNA__20702__RESET_B repeater190/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19851_ _20042_/CLK _19851_/D repeater219/X vssd1 vssd1 vccd1 vccd1 _19851_/Q sky130_fd_sc_hd__dfstp_1
X_12186_ _20341_/Q vssd1 vssd1 vccd1 vccd1 _12186_/Y sky130_fd_sc_hd__inv_2
XFILLER_134_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18299__S _18835_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18802_ _18801_/X _16891_/Y _18875_/S vssd1 vssd1 vccd1 vccd1 _18802_/X sky130_fd_sc_hd__mux2_2
X_11137_ _21219_/Q vssd1 vssd1 vccd1 vccd1 _15609_/B sky130_fd_sc_hd__buf_1
XFILLER_205_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19782_ _19828_/CLK _19782_/D vssd1 vssd1 vccd1 vccd1 _19782_/Q sky130_fd_sc_hd__dfxtp_1
X_16994_ _16994_/A _16994_/B vssd1 vssd1 vccd1 vccd1 _16994_/Y sky130_fd_sc_hd__nor2_1
XFILLER_237_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18733_ _17632_/Y _09734_/Y _18928_/S vssd1 vssd1 vccd1 vccd1 _18733_/X sky130_fd_sc_hd__mux2_1
X_15945_ _15945_/A vssd1 vssd1 vccd1 vccd1 _15945_/X sky130_fd_sc_hd__buf_1
X_11068_ _21239_/Q _11051_/X _11066_/A _09724_/Y _11067_/X vssd1 vssd1 vccd1 vccd1
+ _11069_/A sky130_fd_sc_hd__o32a_1
XFILLER_237_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10019_ _21106_/Q _21105_/Q _21107_/Q _21104_/Q _21108_/Q vssd1 vssd1 vccd1 vccd1
+ _11621_/A sky130_fd_sc_hd__a41o_1
XFILLER_92_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18664_ _18663_/X _20594_/Q _18907_/S vssd1 vssd1 vccd1 vccd1 _18664_/X sky130_fd_sc_hd__mux2_1
XFILLER_76_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21008__CLK _21009_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15876_ _15876_/A vssd1 vssd1 vccd1 vccd1 _15876_/X sky130_fd_sc_hd__buf_1
XFILLER_221_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17615_ _19627_/Q vssd1 vssd1 vccd1 vccd1 _17615_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14827_ _20105_/Q vssd1 vssd1 vccd1 vccd1 _14882_/A sky130_fd_sc_hd__inv_2
X_18595_ _18594_/X _17848_/Y _18874_/S vssd1 vssd1 vccd1 vccd1 _18595_/X sky130_fd_sc_hd__mux2_1
XFILLER_51_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17546_ _20815_/Q _18879_/S vssd1 vssd1 vccd1 vccd1 _17546_/Y sky130_fd_sc_hd__nand2_1
XFILLER_45_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14758_ _19123_/X _14758_/B vssd1 vssd1 vccd1 vccd1 _14758_/Y sky130_fd_sc_hd__nand2_1
XFILLER_44_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13709_ _20335_/Q _13706_/X _13707_/X _13708_/X vssd1 vssd1 vccd1 vccd1 _20335_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_20_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17477_ _18776_/X _17397_/X _18773_/X _17398_/X _17476_/X vssd1 vssd1 vccd1 vccd1
+ _17477_/X sky130_fd_sc_hd__o221a_1
XFILLER_149_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18762__S _18926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14689_ _14692_/A vssd1 vssd1 vccd1 vccd1 _14696_/A sky130_fd_sc_hd__inv_2
X_19216_ _19212_/X _19213_/X _19214_/X _19215_/X _21005_/Q _21006_/Q vssd1 vssd1 vccd1
+ vccd1 _19216_/X sky130_fd_sc_hd__mux4_2
X_16428_ _16428_/A vssd1 vssd1 vccd1 vccd1 _16428_/X sky130_fd_sc_hd__buf_1
XFILLER_177_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19147_ _19682_/Q _19810_/Q _19802_/Q _19794_/Q _19285_/S0 _21017_/Q vssd1 vssd1
+ vccd1 vccd1 _19147_/X sky130_fd_sc_hd__mux4_2
X_16359_ _17072_/B vssd1 vssd1 vccd1 vccd1 _17073_/B sky130_fd_sc_hd__inv_2
XFILLER_145_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09685__A _10892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15325__A1 _20031_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19078_ _16725_/X _20897_/Q _19908_/D vssd1 vssd1 vccd1 vccd1 _19078_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13336__B1 _13270_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18029_ _18029_/A _18032_/B vssd1 vssd1 vccd1 vccd1 _18029_/Y sky130_fd_sc_hd__nor2_1
XFILLER_133_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_246_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21040_ _21040_/CLK _21040_/D repeater247/X vssd1 vssd1 vccd1 vccd1 _21040_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_99_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09802_ _09802_/A vssd1 vssd1 vccd1 vccd1 _21457_/D sky130_fd_sc_hd__inv_2
XFILLER_114_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09733_ _21229_/Q vssd1 vssd1 vccd1 vccd1 _11054_/A sky130_fd_sc_hd__inv_2
XFILLER_86_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18937__S _18946_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11455__A _21043_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09664_ _21472_/Q _09657_/X _09663_/X _09660_/X vssd1 vssd1 vccd1 vccd1 _21472_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_54_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09595_ _13047_/A vssd1 vssd1 vccd1 vccd1 _12753_/A sky130_fd_sc_hd__buf_1
XPHY_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20824_ _21238_/CLK _20824_/D repeater251/X vssd1 vssd1 vccd1 vccd1 _20824_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21231__RESET_B repeater249/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20755_ _21481_/CLK _20755_/D repeater205/X vssd1 vssd1 vccd1 vccd1 _20755_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__10625__B2 _10619_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20686_ _21486_/CLK _20686_/D repeater199/X vssd1 vssd1 vccd1 vccd1 _20686_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_7_0_HCLK clkbuf_3_7_0_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_155_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15597__A _15603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10370_ _21373_/Q _10369_/Y _10364_/X _10289_/B vssd1 vssd1 vccd1 vccd1 _21373_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_164_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21307_ _21481_/CLK _21307_/D repeater206/X vssd1 vssd1 vccd1 vccd1 _21307_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_3_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12040_ _20977_/Q _12038_/Y _12304_/A _20364_/Q vssd1 vssd1 vccd1 vccd1 _12040_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_105_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21238_ _21238_/CLK _21238_/D repeater189/X vssd1 vssd1 vccd1 vccd1 _21238_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_120_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19008__S _19019_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21169_ _21184_/CLK _21169_/D repeater220/X vssd1 vssd1 vccd1 vccd1 _21169_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_172_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13991_ _14004_/A vssd1 vssd1 vccd1 vccd1 _13991_/X sky130_fd_sc_hd__buf_2
XANTENNA__18847__S _18898_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15730_ _16235_/A vssd1 vssd1 vccd1 vccd1 _15730_/X sky130_fd_sc_hd__buf_1
X_12942_ _12960_/A vssd1 vssd1 vccd1 vccd1 _12942_/X sky130_fd_sc_hd__buf_1
XFILLER_46_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19889__D _19889_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15661_ _15661_/A vssd1 vssd1 vccd1 vccd1 _15661_/X sky130_fd_sc_hd__buf_1
XPHY_4230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12873_ _20742_/Q _12867_/X _12872_/X _12868_/X vssd1 vssd1 vccd1 vccd1 _20742_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13580__A _13594_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17400_ _18810_/X _17397_/X _18807_/X _17398_/X _17399_/X vssd1 vssd1 vccd1 vccd1
+ _17400_/X sky130_fd_sc_hd__o221a_1
XPHY_4252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14612_ _14589_/A _14589_/B _14607_/X _14609_/Y vssd1 vssd1 vccd1 vccd1 _20200_/D
+ sky130_fd_sc_hd__a211oi_4
XFILLER_33_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18380_ _18379_/X _16914_/A _18680_/S vssd1 vssd1 vccd1 vccd1 _18380_/X sky130_fd_sc_hd__mux2_2
X_11824_ _11824_/A vssd1 vssd1 vccd1 vccd1 _11825_/B sky130_fd_sc_hd__inv_2
XPHY_4274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15592_ _15592_/A vssd1 vssd1 vccd1 vccd1 _15592_/X sky130_fd_sc_hd__clkbuf_2
XPHY_4285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17331_ _19640_/Q vssd1 vssd1 vccd1 vccd1 _17331_/Y sky130_fd_sc_hd__inv_2
XFILLER_187_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14543_ _14557_/A _15902_/B vssd1 vssd1 vccd1 vccd1 _14561_/A sky130_fd_sc_hd__or2_2
X_11755_ _11755_/A vssd1 vssd1 vccd1 vccd1 _11755_/Y sky130_fd_sc_hd__inv_2
XPHY_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18582__S _18884_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10706_ _10706_/A _10706_/B vssd1 vssd1 vccd1 vccd1 _10711_/A sky130_fd_sc_hd__or2_1
XPHY_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17262_ _19607_/Q vssd1 vssd1 vccd1 vccd1 _17262_/Y sky130_fd_sc_hd__inv_2
X_14474_ _14488_/A vssd1 vssd1 vccd1 vccd1 _14474_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__21450__CLK _21452_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11686_ _12550_/A vssd1 vssd1 vccd1 vccd1 _11686_/X sky130_fd_sc_hd__buf_1
XPHY_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19001_ _16995_/X _20422_/Q _19019_/S vssd1 vssd1 vccd1 vccd1 _19975_/D sky130_fd_sc_hd__mux2_1
X_16213_ _19431_/Q _16206_/X _16212_/X _16208_/X vssd1 vssd1 vccd1 vccd1 _19431_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__20954__RESET_B repeater186/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13425_ _20478_/Q _13417_/X _13424_/X _13420_/X vssd1 vssd1 vccd1 vccd1 _20478_/D
+ sky130_fd_sc_hd__a22o_1
X_10637_ _21337_/Q _10634_/Y _10708_/A _20748_/Q _10636_/X vssd1 vssd1 vccd1 vccd1
+ _10638_/D sky130_fd_sc_hd__o221a_1
X_17193_ _20810_/Q _17193_/B vssd1 vssd1 vccd1 vccd1 _17193_/Y sky130_fd_sc_hd__nor2_1
XFILLER_139_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16144_ _19465_/Q _16141_/X _16142_/X _16143_/X vssd1 vssd1 vccd1 vccd1 _19465_/D
+ sky130_fd_sc_hd__a22o_1
X_10568_ _21332_/Q vssd1 vssd1 vccd1 vccd1 _10569_/A sky130_fd_sc_hd__inv_2
XFILLER_143_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13356_ _20514_/Q _13351_/X _13223_/X _13352_/X vssd1 vssd1 vccd1 vccd1 _20514_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13318__B1 _13243_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12307_ _12307_/A _12386_/A vssd1 vssd1 vccd1 vccd1 _12308_/B sky130_fd_sc_hd__or2_2
X_16075_ _19495_/Q _16071_/X _15774_/X _16072_/X vssd1 vssd1 vccd1 vccd1 _19495_/D
+ sky130_fd_sc_hd__a22o_1
X_10499_ _20678_/Q vssd1 vssd1 vccd1 vccd1 _10499_/Y sky130_fd_sc_hd__inv_2
X_13287_ input53/X vssd1 vssd1 vccd1 vccd1 _13287_/X sky130_fd_sc_hd__buf_2
XFILLER_216_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19903_ _21185_/CLK _19903_/D repeater221/X vssd1 vssd1 vccd1 vccd1 _19903_/Q sky130_fd_sc_hd__dfrtp_1
X_15026_ _15019_/A _15019_/B _20076_/Q _14964_/X _14958_/X vssd1 vssd1 vccd1 vccd1
+ _20076_/D sky130_fd_sc_hd__o221a_1
X_12238_ _12420_/A _20511_/Q _20931_/Q _12234_/Y _12237_/X vssd1 vssd1 vccd1 vccd1
+ _12255_/A sky130_fd_sc_hd__o221a_1
XFILLER_96_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12169_ _20343_/Q vssd1 vssd1 vccd1 vccd1 _12169_/Y sky130_fd_sc_hd__inv_2
X_19834_ _19834_/CLK _19834_/D vssd1 vssd1 vccd1 vccd1 _19834_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16977_ _17013_/A _16977_/B vssd1 vssd1 vccd1 vccd1 _16977_/Y sky130_fd_sc_hd__nor2_1
X_19765_ _19765_/CLK _19765_/D vssd1 vssd1 vccd1 vccd1 _19765_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_209_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18757__S _18926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput5 HADDR[13] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_1
XFILLER_77_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18716_ _18845_/A0 _10441_/Y _18896_/S vssd1 vssd1 vccd1 vccd1 _18716_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15928_ _15928_/A vssd1 vssd1 vccd1 vccd1 _15928_/X sky130_fd_sc_hd__buf_1
XFILLER_237_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19696_ _19776_/CLK _19696_/D vssd1 vssd1 vccd1 vccd1 _19696_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18647_ _17079_/Y _15251_/Y _18908_/S vssd1 vssd1 vccd1 vccd1 _18647_/X sky130_fd_sc_hd__mux2_1
X_15859_ _19600_/Q _15856_/X _15791_/X _15857_/X vssd1 vssd1 vccd1 vccd1 _19600_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_64_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18578_ _18577_/X _16791_/A _18667_/S vssd1 vssd1 vccd1 vccd1 _18578_/X sky130_fd_sc_hd__mux2_1
XFILLER_240_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12818__B _17212_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17529_ _19340_/Q _19339_/Q _19338_/Q _19337_/Q vssd1 vssd1 vccd1 vccd1 _17529_/Y
+ sky130_fd_sc_hd__nor4_2
XANTENNA__10607__B2 _10606_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18492__S _18907_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20540_ _20592_/CLK _20540_/D repeater265/X vssd1 vssd1 vccd1 vccd1 _20540_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_20_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20471_ _20937_/CLK _20471_/D repeater279/X vssd1 vssd1 vccd1 vccd1 _20471_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_118_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20624__RESET_B repeater193/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18496__A0 _17079_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13309__B1 _13151_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18799__A1 _11123_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21023_ _21223_/CLK _21023_/D repeater241/X vssd1 vssd1 vccd1 vccd1 _21023_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17137__A _21056_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18667__S _18667_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21483__RESET_B repeater200/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09716_ _09792_/A _09803_/A _09793_/C _09716_/D vssd1 vssd1 vccd1 vccd1 _09787_/B
+ sky130_fd_sc_hd__or4_4
XANTENNA__19370__CLK _19706_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09647_ _21477_/Q _09643_/X _09645_/X _09646_/X vssd1 vssd1 vccd1 vccd1 _21477_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_71_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12728__B _13108_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20807_ _21011_/CLK _20807_/D repeater237/X vssd1 vssd1 vccd1 vccd1 _20807_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18723__A1 _13951_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11540_ _12502_/A _12502_/B _18969_/X vssd1 vssd1 vccd1 vccd1 _16568_/C sky130_fd_sc_hd__or3b_1
XPHY_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20738_ _21321_/CLK _20738_/D repeater205/X vssd1 vssd1 vccd1 vccd1 _20738_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17957__D _17957_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13548__B1 _13547_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11471_ _19096_/X _11468_/X _21162_/Q _11469_/X vssd1 vssd1 vccd1 vccd1 _21162_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_109_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20669_ _21306_/CLK _20669_/D repeater207/X vssd1 vssd1 vccd1 vccd1 _20669_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10422_ _21308_/Q vssd1 vssd1 vccd1 vccd1 _10422_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18487__A0 _17079_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13210_ _20587_/Q _13206_/X _13209_/X _13207_/X vssd1 vssd1 vccd1 vccd1 _20587_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_109_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14190_ _14190_/A vssd1 vssd1 vccd1 vccd1 _14190_/Y sky130_fd_sc_hd__inv_2
XFILLER_164_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13141_ _13141_/A vssd1 vssd1 vccd1 vccd1 _13167_/A sky130_fd_sc_hd__buf_1
X_10353_ _21352_/Q _17812_/A _21369_/Q _10352_/Y vssd1 vssd1 vccd1 vccd1 _10353_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_152_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13072_ _13072_/A vssd1 vssd1 vccd1 vccd1 _13072_/X sky130_fd_sc_hd__buf_1
Xclkbuf_leaf_120_HCLK clkbuf_opt_3_HCLK/A vssd1 vssd1 vccd1 vccd1 _20982_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_input56_A HWDATA[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10284_ _10284_/A _10377_/A vssd1 vssd1 vccd1 vccd1 _10285_/B sky130_fd_sc_hd__or2_1
X_12023_ _12029_/A vssd1 vssd1 vccd1 vccd1 _12023_/X sky130_fd_sc_hd__buf_1
X_16900_ _19954_/Q vssd1 vssd1 vccd1 vccd1 _16902_/A sky130_fd_sc_hd__inv_2
XANTENNA__13575__A _13595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17880_ _18439_/X _17856_/X _18428_/X _17569_/X _17879_/X vssd1 vssd1 vccd1 vccd1
+ _17880_/X sky130_fd_sc_hd__o221a_1
XFILLER_238_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16831_ _16848_/A vssd1 vssd1 vccd1 vccd1 _16831_/X sky130_fd_sc_hd__buf_1
XANTENNA__18577__S _18666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19550_ _19706_/CLK _19550_/D vssd1 vssd1 vccd1 vccd1 _19550_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_219_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16762_ _16779_/A vssd1 vssd1 vccd1 vccd1 _16762_/X sky130_fd_sc_hd__buf_1
XFILLER_46_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_108_HCLK_A clkbuf_4_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13974_ _13974_/A _13974_/B _13974_/C _13973_/X vssd1 vssd1 vccd1 vccd1 _13974_/X
+ sky130_fd_sc_hd__or4b_4
XFILLER_19_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18501_ _18500_/X _12222_/Y _18910_/S vssd1 vssd1 vccd1 vccd1 _18501_/X sky130_fd_sc_hd__mux2_1
XANTENNA__18411__A0 _18848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_219_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15713_ _19668_/Q _15709_/X _15661_/X _15711_/X vssd1 vssd1 vccd1 vccd1 _19668_/D
+ sky130_fd_sc_hd__a22o_1
X_19481_ _20890_/CLK _19481_/D vssd1 vssd1 vccd1 vccd1 _19481_/Q sky130_fd_sc_hd__dfxtp_1
X_12925_ input48/X vssd1 vssd1 vccd1 vccd1 _12925_/X sky130_fd_sc_hd__clkbuf_4
X_16693_ _16720_/A vssd1 vssd1 vccd1 vccd1 _16700_/A sky130_fd_sc_hd__buf_1
XFILLER_234_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18432_ _17896_/Y _20447_/Q _18906_/S vssd1 vssd1 vccd1 vccd1 _18432_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15644_ _19700_/Q _15640_/X _15473_/X _15642_/X vssd1 vssd1 vccd1 vccd1 _19700_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12856_ _20751_/Q _12848_/X _12855_/X _12851_/X vssd1 vssd1 vccd1 vccd1 _20751_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17281__D_N _17193_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18363_ _18362_/X _16994_/A _18680_/S vssd1 vssd1 vccd1 vccd1 _18363_/X sky130_fd_sc_hd__mux2_1
X_11807_ _11807_/A _11850_/A vssd1 vssd1 vccd1 vccd1 _11848_/B sky130_fd_sc_hd__nor2_1
X_15575_ _16325_/A _15624_/B _16451_/C vssd1 vssd1 vccd1 vccd1 _15584_/A sky130_fd_sc_hd__or3_4
XPHY_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12787_ _20788_/Q _12784_/X _09641_/X _12786_/X vssd1 vssd1 vccd1 vccd1 _20788_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17314_ _17575_/A vssd1 vssd1 vccd1 vccd1 _17862_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_202_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14526_ _20208_/Q vssd1 vssd1 vccd1 vccd1 _14526_/Y sky130_fd_sc_hd__inv_2
XFILLER_230_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11738_ _21059_/Q _11735_/X _11736_/X _11737_/X vssd1 vssd1 vccd1 vccd1 _21059_/D
+ sky130_fd_sc_hd__a22o_1
X_18294_ _18293_/X _20279_/Q _18904_/S vssd1 vssd1 vccd1 vccd1 _18294_/X sky130_fd_sc_hd__mux2_1
XFILLER_41_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17245_ _19383_/Q vssd1 vssd1 vccd1 vccd1 _17245_/Y sky130_fd_sc_hd__inv_2
X_14457_ _14382_/A _14382_/B _14383_/Y _14524_/C vssd1 vssd1 vccd1 vccd1 _20239_/D
+ sky130_fd_sc_hd__a211oi_2
X_11669_ _11669_/A vssd1 vssd1 vccd1 vccd1 _21091_/D sky130_fd_sc_hd__inv_2
XPHY_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18478__A0 _18848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13408_ _20486_/Q _13404_/X _13211_/X _13405_/X vssd1 vssd1 vccd1 vccd1 _20486_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_162_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17176_ _20108_/Q vssd1 vssd1 vccd1 vccd1 _17176_/Y sky130_fd_sc_hd__inv_2
X_14388_ _21483_/Q _14336_/A _20238_/Q _14387_/Y vssd1 vssd1 vccd1 vccd1 _14394_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_183_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16127_ _16127_/A vssd1 vssd1 vccd1 vccd1 _16127_/X sky130_fd_sc_hd__clkbuf_2
X_13339_ _13351_/A vssd1 vssd1 vccd1 vccd1 _13339_/X sky130_fd_sc_hd__buf_1
XFILLER_227_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15161__C1 _15160_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16058_ _19505_/Q _16056_/X _15769_/X _16057_/X vssd1 vssd1 vccd1 vccd1 _19505_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_170_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13485__A input47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13711__B1 _13710_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15009_ _15009_/A vssd1 vssd1 vccd1 vccd1 _15009_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18650__A0 _18848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19817_ _20172_/CLK _19817_/D vssd1 vssd1 vccd1 vccd1 _19817_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_229_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18487__S _18908_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19748_ _19811_/CLK _19748_/D vssd1 vssd1 vccd1 vccd1 _19748_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__19971__RESET_B repeater184/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19679_ _19820_/CLK _19679_/D vssd1 vssd1 vccd1 vccd1 _19679_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__18953__A1 _21083_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12829__A _12841_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11733__A _13163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_240_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20805__RESET_B repeater235/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12450__B1 _12445_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20523_ _20944_/CLK _20523_/D repeater277/X vssd1 vssd1 vccd1 vccd1 _20523_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18950__S _18962_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20454_ _20476_/CLK _20454_/D repeater279/X vssd1 vssd1 vccd1 vccd1 _20454_/Q sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_143_HCLK clkbuf_4_3_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _21218_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_21_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20385_ _20971_/CLK _20385_/D repeater280/X vssd1 vssd1 vccd1 vccd1 _20385_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_133_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19736__CLK _19765_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13702__B1 _13509_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21006_ _21009_/CLK _21006_/D repeater235/X vssd1 vssd1 vccd1 vccd1 _21006_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__18397__S _18879_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_248_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15455__B1 _15454_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10971_ _11800_/A vssd1 vssd1 vccd1 vccd1 _11964_/A sky130_fd_sc_hd__inv_2
XFILLER_16_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12710_ _20813_/Q _12707_/X _11739_/X _12708_/X vssd1 vssd1 vccd1 vccd1 _20813_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_71_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13690_ _20346_/Q _13686_/X _12853_/A _13688_/X vssd1 vssd1 vccd1 vccd1 _20346_/D
+ sky130_fd_sc_hd__a22o_1
X_12641_ input23/X _12637_/X _20845_/Q _12638_/X vssd1 vssd1 vccd1 vccd1 _20845_/D
+ sky130_fd_sc_hd__o22a_1
XPHY_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19021__S _19026_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_212_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15360_ _15366_/A vssd1 vssd1 vccd1 vccd1 _15367_/A sky130_fd_sc_hd__inv_2
XFILLER_12_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12572_ _13188_/A _12566_/X _18242_/X _18242_/S vssd1 vssd1 vccd1 vccd1 _20890_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12992__A1 _20695_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14311_ _14796_/A vssd1 vssd1 vccd1 vccd1 _14311_/X sky130_fd_sc_hd__clkbuf_2
XPHY_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11523_ _10894_/A _21144_/Q _11523_/S vssd1 vssd1 vccd1 vccd1 _21144_/D sky130_fd_sc_hd__mux2_1
XFILLER_8_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15291_ _19857_/Q _15291_/B vssd1 vssd1 vccd1 vccd1 _15292_/B sky130_fd_sc_hd__or2_1
XFILLER_178_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17030_ _21251_/Q _11017_/A _17029_/Y _21244_/Q _11584_/C vssd1 vssd1 vccd1 vccd1
+ _18993_/S sky130_fd_sc_hd__a221oi_2
X_14242_ _19902_/Q _14242_/B vssd1 vssd1 vccd1 vccd1 _14243_/B sky130_fd_sc_hd__or2_1
XPHY_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11454_ _21166_/Q _11454_/B vssd1 vssd1 vccd1 vccd1 _11454_/X sky130_fd_sc_hd__or2_2
XANTENNA__17984__B _18007_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12744__A1 _12968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10405_ _10405_/A _10405_/B _10405_/C vssd1 vssd1 vccd1 vccd1 _21354_/D sky130_fd_sc_hd__nor3_1
XANTENNA__13941__B1 _13939_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11385_ _11385_/A _21168_/Q _21184_/Q _11385_/D vssd1 vssd1 vccd1 vccd1 _11388_/B
+ sky130_fd_sc_hd__or4_4
X_14173_ _14205_/A vssd1 vssd1 vccd1 vccd1 _14191_/A sky130_fd_sc_hd__buf_1
XFILLER_180_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13124_ _20624_/Q _13120_/X _13001_/X _13121_/X vssd1 vssd1 vccd1 vccd1 _20624_/D
+ sky130_fd_sc_hd__a22o_1
X_10336_ _20713_/Q vssd1 vssd1 vccd1 vccd1 _10336_/Y sky130_fd_sc_hd__inv_2
X_18981_ _21425_/Q _21098_/Q _18983_/S vssd1 vssd1 vccd1 vccd1 _18981_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17932_ _17932_/A vssd1 vssd1 vccd1 vccd1 _17932_/X sky130_fd_sc_hd__clkbuf_2
X_13055_ _13073_/A vssd1 vssd1 vccd1 vccd1 _13055_/X sky130_fd_sc_hd__buf_1
X_10267_ _10267_/A _10409_/A vssd1 vssd1 vccd1 vccd1 _10268_/B sky130_fd_sc_hd__or2_2
XANTENNA__21334__RESET_B repeater203/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12006_ _12006_/A _19888_/D _12006_/C vssd1 vssd1 vccd1 vccd1 _12006_/X sky130_fd_sc_hd__or3_4
XFILLER_238_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17863_ _18576_/X _17839_/X _18562_/X _17840_/X vssd1 vssd1 vccd1 vccd1 _17863_/X
+ sky130_fd_sc_hd__o22a_1
X_10198_ _10149_/A _10149_/B _10196_/Y _10227_/C vssd1 vssd1 vccd1 vccd1 _21388_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_238_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19602_ _19821_/CLK _19602_/D vssd1 vssd1 vccd1 vccd1 _19602_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_213_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16814_ _16822_/C vssd1 vssd1 vccd1 vccd1 _16814_/Y sky130_fd_sc_hd__inv_2
X_17794_ _21193_/Q vssd1 vssd1 vccd1 vccd1 _17794_/Y sky130_fd_sc_hd__inv_2
X_19533_ _19784_/CLK _19533_/D vssd1 vssd1 vccd1 vccd1 _19533_/Q sky130_fd_sc_hd__dfxtp_1
X_16745_ _20771_/Q vssd1 vssd1 vccd1 vccd1 _16848_/A sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_24_HCLK clkbuf_4_9_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _21421_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_35_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13957_ _20647_/Q vssd1 vssd1 vccd1 vccd1 _13957_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18935__A1 _21141_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19283__S1 _21017_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19464_ _21234_/CLK _19464_/D vssd1 vssd1 vccd1 vccd1 _19464_/Q sky130_fd_sc_hd__dfxtp_1
X_12908_ _20731_/Q _12901_/X _12660_/X _12904_/X vssd1 vssd1 vccd1 vccd1 _20731_/D
+ sky130_fd_sc_hd__a22o_1
X_16676_ _21164_/Q _11452_/B _11453_/B vssd1 vssd1 vccd1 vccd1 _16676_/X sky130_fd_sc_hd__a21bo_1
X_13888_ _13971_/A _13993_/A vssd1 vssd1 vccd1 vccd1 _13889_/B sky130_fd_sc_hd__or2_2
X_18415_ _18414_/X _16936_/Y _18680_/S vssd1 vssd1 vccd1 vccd1 _18415_/X sky130_fd_sc_hd__mux2_2
X_15627_ _15633_/A vssd1 vssd1 vccd1 vccd1 _15627_/X sky130_fd_sc_hd__buf_1
X_12839_ _20759_/Q _12835_/X _09626_/X _12836_/X vssd1 vssd1 vccd1 vccd1 _20759_/D
+ sky130_fd_sc_hd__a22o_1
X_19395_ _21001_/CLK _19395_/D vssd1 vssd1 vccd1 vccd1 _19395_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18346_ _18345_/X _12153_/Y _18787_/S vssd1 vssd1 vccd1 vccd1 _18346_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15558_ _19742_/Q _15553_/X _15526_/X _15554_/X vssd1 vssd1 vccd1 vccd1 _19742_/D
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_166_HCLK clkbuf_opt_0_HCLK/A vssd1 vssd1 vccd1 vccd1 _21459_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__20216__RESET_B repeater202/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14509_ _14502_/A _14502_/B _14507_/Y _14469_/X vssd1 vssd1 vccd1 vccd1 _20217_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_174_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18277_ _19176_/X _21272_/Q _18281_/S vssd1 vssd1 vccd1 vccd1 _18277_/X sky130_fd_sc_hd__mux2_1
XFILLER_159_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18770__S _18880_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15489_ _16451_/A vssd1 vssd1 vccd1 vccd1 _16325_/A sky130_fd_sc_hd__buf_1
XFILLER_174_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17228_ _17228_/A vssd1 vssd1 vccd1 vccd1 _17732_/A sky130_fd_sc_hd__clkbuf_2
Xinput30 HADDR[7] vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__19759__CLK _19765_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput41 HWDATA[12] vssd1 vssd1 vccd1 vccd1 input41/X sky130_fd_sc_hd__buf_2
XANTENNA__19112__A1 _21071_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput52 HWDATA[22] vssd1 vssd1 vccd1 vccd1 input52/X sky130_fd_sc_hd__buf_2
Xinput63 HWDATA[3] vssd1 vssd1 vccd1 vccd1 input63/X sky130_fd_sc_hd__buf_6
XFILLER_116_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput74 RsRx_S1 vssd1 vssd1 vccd1 vccd1 input74/X sky130_fd_sc_hd__buf_6
XFILLER_7_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17159_ _17144_/X _17156_/X _17158_/X vssd1 vssd1 vccd1 vccd1 _17159_/Y sky130_fd_sc_hd__a21oi_1
X_20170_ _21120_/CLK _20170_/D repeater233/X vssd1 vssd1 vccd1 vccd1 _20170_/Q sky130_fd_sc_hd__dfrtp_1
X_09981_ _21413_/Q _09975_/A _09698_/X _09976_/A vssd1 vssd1 vccd1 vccd1 _21413_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_170_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15685__B1 _15590_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14104__A _20538_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18623__A0 _18848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21004__RESET_B repeater235/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19106__S _19870_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13943__A _20637_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_226_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09667__A1 _21471_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18945__S _18946_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19274__S1 _21004_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_154_HCLK_A clkbuf_opt_1_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12671__B1 _12670_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18680__S _18680_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20506_ _20947_/CLK _20506_/D repeater266/X vssd1 vssd1 vccd1 vccd1 _20506_/Q sky130_fd_sc_hd__dfrtp_4
X_21486_ _21486_/CLK _21486_/D repeater209/X vssd1 vssd1 vccd1 vccd1 _21486_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_147_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20437_ _20476_/CLK _20437_/D repeater279/X vssd1 vssd1 vccd1 vccd1 _20437_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_4_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11170_ _11170_/A vssd1 vssd1 vccd1 vccd1 _11170_/Y sky130_fd_sc_hd__inv_2
XFILLER_107_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20368_ _20422_/CLK _20368_/D repeater271/X vssd1 vssd1 vccd1 vccd1 _20368_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_106_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17665__B2 _17655_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10121_ _10041_/A _20776_/Q _10040_/A _20774_/Q _10120_/X vssd1 vssd1 vccd1 vccd1
+ _10122_/D sky130_fd_sc_hd__o221a_1
XFILLER_164_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20299_ _20693_/CLK _20299_/D repeater197/X vssd1 vssd1 vccd1 vccd1 _20299_/Q sky130_fd_sc_hd__dfrtp_1
X_10052_ _10206_/A _10205_/A _10052_/C _10207_/A vssd1 vssd1 vccd1 vccd1 _10053_/D
+ sky130_fd_sc_hd__or4_4
Xclkbuf_leaf_47_HCLK _20004_/CLK vssd1 vssd1 vccd1 vccd1 _21164_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_102_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_248_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19016__S _19019_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14860_ _20084_/Q vssd1 vssd1 vccd1 vccd1 _15004_/A sky130_fd_sc_hd__inv_2
XFILLER_235_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13811_ _13811_/A _13811_/B _13811_/C _13811_/D vssd1 vssd1 vccd1 vccd1 _13837_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_17_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14791_ _20119_/Q vssd1 vssd1 vccd1 vccd1 _14791_/Y sky130_fd_sc_hd__inv_2
XANTENNA_input19_A HADDR[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18855__S _18909_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19265__S1 _21004_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16530_ _16688_/B vssd1 vssd1 vccd1 vccd1 _16530_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20727__RESET_B repeater257/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13742_ _13736_/Y _20207_/Q _20608_/Q _13738_/X _13741_/X vssd1 vssd1 vccd1 vccd1
+ _13761_/A sky130_fd_sc_hd__o221a_1
X_10954_ _21204_/Q _11848_/A _21204_/Q _21031_/Q vssd1 vssd1 vccd1 vccd1 _10954_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_113_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16461_ _19303_/Q _16459_/X _16335_/X _16460_/X vssd1 vssd1 vccd1 vccd1 _19303_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_231_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13673_ _13679_/A vssd1 vssd1 vccd1 vccd1 _13673_/X sky130_fd_sc_hd__buf_1
XANTENNA_clkbuf_leaf_13_HCLK_A clkbuf_4_3_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10885_ _21257_/Q _10879_/X _10884_/X _10881_/X vssd1 vssd1 vccd1 vccd1 _21257_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_204_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18200_ _17281_/X _17959_/Y _18835_/S vssd1 vssd1 vccd1 vccd1 _18200_/X sky130_fd_sc_hd__mux2_1
XFILLER_231_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15412_ _15673_/A vssd1 vssd1 vccd1 vccd1 _15528_/A sky130_fd_sc_hd__buf_1
XPHY_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_76_HCLK_A clkbuf_4_13_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19180_ _19303_/Q _19825_/Q _19833_/Q _19417_/Q _19280_/S0 _20122_/Q vssd1 vssd1
+ vccd1 vccd1 _19180_/X sky130_fd_sc_hd__mux4_2
X_12624_ input5/X _12619_/X _20856_/Q _12620_/X vssd1 vssd1 vccd1 vccd1 _20856_/D
+ sky130_fd_sc_hd__o22a_1
XPHY_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16392_ _16399_/A vssd1 vssd1 vccd1 vccd1 _16392_/X sky130_fd_sc_hd__buf_1
XPHY_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_1_HCLK_A clkbuf_opt_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18131_ _18845_/A0 _13770_/Y _18896_/S vssd1 vssd1 vccd1 vccd1 _18131_/X sky130_fd_sc_hd__mux2_1
XPHY_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15343_ _15421_/A vssd1 vssd1 vccd1 vccd1 _15343_/X sky130_fd_sc_hd__buf_2
XANTENNA__17995__A _18064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12555_ _20896_/Q _12553_/X _11736_/X _12554_/X vssd1 vssd1 vccd1 vccd1 _20896_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_156_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18590__S _18907_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_repeater158_A _18850_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11506_ _10892_/A _11487_/X _11498_/A _11500_/Y _21148_/Q vssd1 vssd1 vccd1 vccd1
+ _21148_/D sky130_fd_sc_hd__a32o_1
X_18062_ _18258_/X _18021_/X _18255_/X _18045_/X vssd1 vssd1 vccd1 vccd1 _18062_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_156_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15274_ _20491_/Q _15084_/A _20470_/Q _15064_/A vssd1 vssd1 vccd1 vccd1 _15274_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_144_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12486_ _12486_/A vssd1 vssd1 vccd1 vccd1 _12486_/Y sky130_fd_sc_hd__inv_2
X_17013_ _17013_/A _17013_/B vssd1 vssd1 vccd1 vccd1 _17013_/Y sky130_fd_sc_hd__nor2_1
X_14225_ _14225_/A vssd1 vssd1 vccd1 vccd1 _14225_/Y sky130_fd_sc_hd__inv_2
X_11437_ _19917_/Q vssd1 vssd1 vccd1 vccd1 _11437_/Y sky130_fd_sc_hd__inv_2
XFILLER_208_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12932__A input45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18853__A0 _18852_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output87_A _17957_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14156_ _20533_/Q vssd1 vssd1 vccd1 vccd1 _14156_/Y sky130_fd_sc_hd__inv_2
X_11368_ _21174_/Q vssd1 vssd1 vccd1 vccd1 _11379_/B sky130_fd_sc_hd__buf_1
XFILLER_99_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13107_ _12978_/X _20632_/Q _13107_/S vssd1 vssd1 vccd1 vccd1 _20632_/D sky130_fd_sc_hd__mux2_1
X_10319_ _21344_/Q _10316_/Y _10278_/A _20722_/Q _10318_/X vssd1 vssd1 vccd1 vccd1
+ _10323_/C sky130_fd_sc_hd__o221a_1
X_18964_ _16618_/Y _14529_/B _18976_/S vssd1 vssd1 vccd1 vccd1 _18964_/X sky130_fd_sc_hd__mux2_1
X_14087_ _14087_/A _14087_/B vssd1 vssd1 vccd1 vccd1 _14198_/A sky130_fd_sc_hd__or2_1
X_11299_ _11299_/A _20905_/Q _11299_/C _11299_/D vssd1 vssd1 vccd1 vccd1 _11310_/D
+ sky130_fd_sc_hd__or4_4
XFILLER_224_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13038_ _20671_/Q _13034_/X _12957_/X _13035_/X vssd1 vssd1 vccd1 vccd1 _20671_/D
+ sky130_fd_sc_hd__a22o_1
X_17915_ _18495_/X _18024_/A _18486_/X _17869_/X vssd1 vssd1 vccd1 vccd1 _17915_/X
+ sky130_fd_sc_hd__o22a_1
X_18895_ _18894_/X _17181_/Y _18901_/S vssd1 vssd1 vccd1 vccd1 _18895_/X sky130_fd_sc_hd__mux2_1
XFILLER_239_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13763__A _20601_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17235__A _17235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17846_ _18593_/X _17214_/X _18599_/X _17203_/X _17845_/X vssd1 vssd1 vccd1 vccd1
+ _17846_/X sky130_fd_sc_hd__o221a_2
XANTENNA__16092__B1 _15916_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14989_ _14989_/A vssd1 vssd1 vccd1 vccd1 _14989_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__18765__S _18929_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17777_ _17777_/A _20116_/Q vssd1 vssd1 vccd1 vccd1 _17777_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__19256__S1 _21006_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19516_ _21445_/CLK _19516_/D vssd1 vssd1 vccd1 vccd1 _19516_/Q sky130_fd_sc_hd__dfxtp_1
X_16728_ _20990_/Q _11996_/B _11997_/B vssd1 vssd1 vccd1 vccd1 _16728_/X sky130_fd_sc_hd__a21bo_1
XFILLER_207_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20289__CLK _20592_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16659_ _16661_/A _18951_/X vssd1 vssd1 vccd1 vccd1 _19863_/D sky130_fd_sc_hd__and2_1
XFILLER_34_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19447_ _21234_/CLK _19447_/D vssd1 vssd1 vccd1 vccd1 _19447_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19378_ _19812_/CLK _19378_/D vssd1 vssd1 vccd1 vccd1 _19378_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20050__RESET_B repeater281/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18329_ _18845_/A0 _13801_/Y _18896_/S vssd1 vssd1 vccd1 vccd1 _18329_/X sky130_fd_sc_hd__mux2_1
X_21340_ _21341_/CLK _21340_/D repeater222/X vssd1 vssd1 vccd1 vccd1 _21340_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_175_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13003__A input54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21271_ _21444_/CLK _21271_/D repeater246/X vssd1 vssd1 vccd1 vccd1 _21271_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12842__A _12842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20222_ _21484_/CLK _20222_/D repeater202/X vssd1 vssd1 vccd1 vccd1 _20222_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__19192__S0 _19280_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13381__A1 _20499_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20153_ _21242_/CLK _20153_/D repeater189/X vssd1 vssd1 vccd1 vccd1 _20153_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_170_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09964_ _11199_/A vssd1 vssd1 vccd1 vccd1 _15312_/A sky130_fd_sc_hd__buf_1
XFILLER_134_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20084_ _20946_/CLK _20084_/D repeater274/X vssd1 vssd1 vccd1 vccd1 _20084_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_76_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09895_ _21257_/Q vssd1 vssd1 vccd1 vccd1 _09895_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17145__A _21080_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13673__A _13679_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21064__CLK _21134_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20891__RESET_B repeater248/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18675__S _18926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19247__S1 _20131_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20986_ _21141_/CLK _20986_/D repeater191/X vssd1 vssd1 vccd1 vccd1 _20986_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_3925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19924__CLK _21342_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20138__RESET_B repeater242/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09598__A _20887_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10670_ _10694_/A vssd1 vssd1 vccd1 vccd1 _10670_/X sky130_fd_sc_hd__buf_1
XFILLER_201_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12340_ _20979_/Q _12339_/Y _12206_/X _12333_/B vssd1 vssd1 vccd1 vccd1 _20979_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_216_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12271_ _12408_/A _12270_/Y _20948_/Q _20528_/Q vssd1 vssd1 vccd1 vccd1 _12271_/X
+ sky130_fd_sc_hd__a22o_1
X_21469_ _21477_/CLK _21469_/D repeater204/X vssd1 vssd1 vccd1 vccd1 _21469_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_107_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19183__S0 _19280_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14010_ _14030_/A _14031_/B _14010_/C vssd1 vssd1 vccd1 vccd1 _14028_/A sky130_fd_sc_hd__or3_1
XANTENNA__18835__A0 _17281_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11222_ _21203_/Q _11219_/X _10886_/X _11220_/X vssd1 vssd1 vccd1 vccd1 _21203_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_134_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11153_ _11153_/A vssd1 vssd1 vccd1 vccd1 _16479_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_1_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20979__RESET_B repeater187/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10104_ _21405_/Q _20802_/Q _21405_/Q _20802_/Q vssd1 vssd1 vccd1 vccd1 _10104_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_11084_ _11084_/A vssd1 vssd1 vccd1 vccd1 _21235_/D sky130_fd_sc_hd__inv_2
X_15961_ _15961_/A vssd1 vssd1 vccd1 vccd1 _15961_/X sky130_fd_sc_hd__buf_1
XFILLER_248_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20908__RESET_B repeater217/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17700_ _19460_/Q vssd1 vssd1 vccd1 vccd1 _17700_/Y sky130_fd_sc_hd__inv_2
X_14912_ _14895_/Y _20092_/Q _14911_/Y _20097_/Q vssd1 vssd1 vccd1 vccd1 _14912_/X
+ sky130_fd_sc_hd__o22a_1
X_10035_ _21405_/Q vssd1 vssd1 vccd1 vccd1 _10076_/C sky130_fd_sc_hd__inv_2
XFILLER_248_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18680_ _18679_/X _16910_/A _18680_/S vssd1 vssd1 vccd1 vccd1 _18680_/X sky130_fd_sc_hd__mux2_2
XFILLER_49_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15892_ _19588_/Q _15886_/X _15891_/X _15889_/X vssd1 vssd1 vccd1 vccd1 _19588_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_236_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14843_ _20091_/Q vssd1 vssd1 vccd1 vccd1 _14962_/A sky130_fd_sc_hd__inv_2
X_17631_ _19314_/Q _17631_/B vssd1 vssd1 vccd1 vccd1 _17631_/X sky130_fd_sc_hd__or2_1
XFILLER_64_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18585__S _18908_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19238__S1 _20131_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20431__CLK _21009_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output125_A _17088_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17562_ _20248_/Q vssd1 vssd1 vccd1 vccd1 _17562_/Y sky130_fd_sc_hd__inv_2
X_14774_ _15448_/A _14292_/X _19125_/X _14315_/Y _14773_/X vssd1 vssd1 vccd1 vccd1
+ _20128_/D sky130_fd_sc_hd__a41o_1
X_11986_ _20999_/Q vssd1 vssd1 vccd1 vccd1 _11986_/Y sky130_fd_sc_hd__inv_2
XFILLER_189_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16513_ _21092_/Q _16498_/Y _16512_/Y _11327_/X _16499_/X vssd1 vssd1 vccd1 vccd1
+ _16513_/Y sky130_fd_sc_hd__o2111ai_4
X_19301_ _19828_/CLK _19301_/D vssd1 vssd1 vccd1 vccd1 _19301_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_216_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13725_ _15764_/A _15766_/A _13725_/S vssd1 vssd1 vccd1 vccd1 _20328_/D sky130_fd_sc_hd__mux2_1
XFILLER_17_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10937_ _10935_/Y _21035_/Q _21208_/Q _11812_/A vssd1 vssd1 vccd1 vccd1 _10937_/X
+ sky130_fd_sc_hd__o22a_1
X_17493_ _19386_/Q vssd1 vssd1 vccd1 vccd1 _17493_/Y sky130_fd_sc_hd__inv_2
XFILLER_204_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16444_ _19311_/Q _16441_/X _16338_/X _16442_/X vssd1 vssd1 vccd1 vccd1 _19311_/D
+ sky130_fd_sc_hd__a22o_1
X_19232_ _17484_/Y _17485_/Y _17486_/Y _17487_/Y _19275_/S0 _21004_/Q vssd1 vssd1
+ vccd1 vccd1 _19232_/X sky130_fd_sc_hd__mux4_2
X_13656_ _20364_/Q _13651_/X _13454_/X _13652_/X vssd1 vssd1 vccd1 vccd1 _20364_/D
+ sky130_fd_sc_hd__a22o_1
X_10868_ _21266_/Q _10864_/X _09676_/X _10866_/X vssd1 vssd1 vccd1 vccd1 _21266_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_231_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19163_ _19542_/Q _19534_/Q _19526_/Q _19510_/Q _19280_/S0 _20122_/Q vssd1 vssd1
+ vccd1 vccd1 _19163_/X sky130_fd_sc_hd__mux4_1
X_12607_ _17060_/B _12600_/X _18221_/X _12601_/X vssd1 vssd1 vccd1 vccd1 _20869_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16375_ _21446_/Q vssd1 vssd1 vccd1 vccd1 _16375_/X sky130_fd_sc_hd__clkbuf_2
X_13587_ _20405_/Q _13580_/X _13586_/X _13581_/X vssd1 vssd1 vccd1 vccd1 _20405_/D
+ sky130_fd_sc_hd__a22o_1
X_10799_ _21302_/Q _10797_/Y _10798_/X _10779_/B vssd1 vssd1 vccd1 vccd1 _21302_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_219_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18114_ _21430_/Q _21112_/Q vssd1 vssd1 vccd1 vccd1 _18114_/X sky130_fd_sc_hd__and2_4
X_15326_ _20030_/Q _15323_/X _13545_/X _15324_/X vssd1 vssd1 vccd1 vccd1 _20030_/D
+ sky130_fd_sc_hd__a22o_1
X_12538_ _11311_/A _12521_/A _16568_/B _12518_/X vssd1 vssd1 vccd1 vccd1 _20904_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_200_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19094_ _16676_/X _21084_/Q _19870_/D vssd1 vssd1 vccd1 vccd1 _19094_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18045_ _18045_/A vssd1 vssd1 vccd1 vccd1 _18045_/X sky130_fd_sc_hd__buf_1
XFILLER_8_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15257_ _20474_/Q vssd1 vssd1 vccd1 vccd1 _15257_/Y sky130_fd_sc_hd__inv_2
X_12469_ _12490_/A _12469_/B _12469_/C vssd1 vssd1 vccd1 vccd1 _12488_/A sky130_fd_sc_hd__or3_1
XANTENNA__19174__S0 _19280_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14208_ _14083_/A _14083_/B _14204_/Y _14207_/X vssd1 vssd1 vccd1 vccd1 _20273_/D
+ sky130_fd_sc_hd__a211oi_2
X_15188_ _15188_/A vssd1 vssd1 vccd1 vccd1 _15188_/Y sky130_fd_sc_hd__inv_2
XFILLER_153_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15973__A _16235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14139_ _20545_/Q vssd1 vssd1 vccd1 vccd1 _14139_/Y sky130_fd_sc_hd__inv_2
XFILLER_235_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19996_ _21055_/CLK _19996_/D repeater220/X vssd1 vssd1 vccd1 vccd1 _19996_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_3_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18947_ _16682_/X _21051_/Q _18947_/S vssd1 vssd1 vccd1 vccd1 _18947_/X sky130_fd_sc_hd__mux2_1
XFILLER_101_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09680_ input65/X vssd1 vssd1 vccd1 vccd1 _15385_/A sky130_fd_sc_hd__buf_1
X_18878_ _18877_/X _17189_/Y _18901_/S vssd1 vssd1 vccd1 vccd1 _18878_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17829_ _18927_/S _17829_/B _18926_/S vssd1 vssd1 vccd1 vccd1 _17830_/A sky130_fd_sc_hd__or3_1
XANTENNA__19229__S1 _20131_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18495__S _18910_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20840_ _20841_/CLK _20840_/D repeater251/X vssd1 vssd1 vccd1 vccd1 _20840_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__20231__RESET_B repeater203/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20771_ _21374_/CLK _20771_/D repeater255/X vssd1 vssd1 vccd1 vccd1 _20771_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11741__A _13171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17317__B1 _18836_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21323_ _21341_/CLK _21323_/D repeater201/X vssd1 vssd1 vccd1 vccd1 _21323_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__13668__A _13680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19165__S0 _19280_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12157__A2 _20346_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18817__A0 _17079_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21254_ _21255_/CLK _21254_/D repeater240/X vssd1 vssd1 vccd1 vccd1 _21254_/Q sky130_fd_sc_hd__dfrtp_1
X_20205_ _20623_/CLK _20205_/D repeater194/X vssd1 vssd1 vccd1 vccd1 _20205_/Q sky130_fd_sc_hd__dfrtp_4
X_21185_ _21185_/CLK _21185_/D repeater221/X vssd1 vssd1 vccd1 vccd1 _21185_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_145_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20136_ _20136_/CLK _20136_/D repeater248/X vssd1 vssd1 vccd1 vccd1 _20136_/Q sky130_fd_sc_hd__dfrtp_4
X_09947_ _20869_/Q vssd1 vssd1 vccd1 vccd1 _12725_/B sky130_fd_sc_hd__buf_1
XFILLER_219_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11668__A1 _16654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20067_ _20070_/CLK _20067_/D repeater276/X vssd1 vssd1 vccd1 vccd1 _20067_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__12865__B1 _12697_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09878_ _09878_/A _09878_/B vssd1 vssd1 vccd1 vccd1 _09878_/Y sky130_fd_sc_hd__nor2_1
XFILLER_38_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20319__RESET_B repeater262/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_245_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater280 repeater281/X vssd1 vssd1 vccd1 vccd1 repeater280/X sky130_fd_sc_hd__buf_8
XPHY_4412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11840_ _11840_/A vssd1 vssd1 vccd1 vccd1 _21034_/D sky130_fd_sc_hd__inv_2
XPHY_4434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11771_ _11771_/A vssd1 vssd1 vccd1 vccd1 _11771_/X sky130_fd_sc_hd__buf_1
XFILLER_54_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20969_ _20971_/CLK _20969_/D repeater186/X vssd1 vssd1 vccd1 vccd1 _20969_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__13290__B1 _13209_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13510_ _20439_/Q _13505_/X _13509_/X _13507_/X vssd1 vssd1 vccd1 vccd1 _20439_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10722_ _10722_/A vssd1 vssd1 vccd1 vccd1 _10723_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_54_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14490_ _14490_/A vssd1 vssd1 vccd1 vccd1 _14490_/Y sky130_fd_sc_hd__inv_2
XPHY_3777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13441_ input64/X vssd1 vssd1 vccd1 vccd1 _15421_/A sky130_fd_sc_hd__clkbuf_2
X_10653_ _10653_/A _10653_/B vssd1 vssd1 vccd1 vccd1 _10693_/A sky130_fd_sc_hd__or2_1
XANTENNA__13042__B1 _12875_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__21178__RESET_B repeater216/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16160_ _19457_/Q _16158_/X _16142_/X _16159_/X vssd1 vssd1 vccd1 vccd1 _19457_/D
+ sky130_fd_sc_hd__a22o_1
X_13372_ _13378_/A vssd1 vssd1 vccd1 vccd1 _13372_/X sky130_fd_sc_hd__buf_1
X_10584_ _20750_/Q vssd1 vssd1 vccd1 vccd1 _10584_/Y sky130_fd_sc_hd__inv_2
XFILLER_70_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15111_ _20439_/Q vssd1 vssd1 vccd1 vccd1 _15111_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12323_ _12323_/A _12323_/B vssd1 vssd1 vccd1 vccd1 _12355_/A sky130_fd_sc_hd__or2_1
XFILLER_186_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16091_ _19487_/Q _16087_/X _15881_/X _16088_/X vssd1 vssd1 vccd1 vccd1 _19487_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_182_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18808__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15042_ _20060_/Q vssd1 vssd1 vccd1 vccd1 _15074_/A sky130_fd_sc_hd__inv_2
X_12254_ _12468_/A _20498_/Q _12422_/A _20513_/Q _12253_/X vssd1 vssd1 vccd1 vccd1
+ _12255_/D sky130_fd_sc_hd__o221a_1
XFILLER_141_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11205_ _11207_/A vssd1 vssd1 vccd1 vccd1 _11225_/A sky130_fd_sc_hd__clkbuf_2
X_19850_ _20042_/CLK _19850_/D repeater219/X vssd1 vssd1 vccd1 vccd1 _19850_/Q sky130_fd_sc_hd__dfstp_1
X_12185_ _12097_/X _20340_/Q _12119_/X _20356_/Q _12184_/X vssd1 vssd1 vccd1 vccd1
+ _12190_/C sky130_fd_sc_hd__o221a_1
X_18801_ _17281_/X _17374_/Y _18835_/S vssd1 vssd1 vccd1 vccd1 _18801_/X sky130_fd_sc_hd__mux2_1
X_11136_ _11136_/A vssd1 vssd1 vccd1 vccd1 _11136_/X sky130_fd_sc_hd__buf_1
XFILLER_95_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19781_ _20432_/CLK _19781_/D vssd1 vssd1 vccd1 vccd1 _19781_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_205_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16993_ _16997_/B vssd1 vssd1 vccd1 vccd1 _16999_/B sky130_fd_sc_hd__inv_2
XFILLER_95_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18732_ _17633_/Y _09907_/Y _20870_/Q vssd1 vssd1 vccd1 vccd1 _18732_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12856__B1 _12855_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15944_ _16335_/A vssd1 vssd1 vccd1 vccd1 _15944_/X sky130_fd_sc_hd__clkbuf_2
X_11067_ _11101_/A _11067_/B vssd1 vssd1 vccd1 vccd1 _11067_/X sky130_fd_sc_hd__and2_1
XFILLER_237_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16047__B1 _16016_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10018_ _11621_/B vssd1 vssd1 vccd1 vccd1 _14813_/D sky130_fd_sc_hd__buf_1
XFILLER_237_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15875_ _15875_/A vssd1 vssd1 vccd1 vccd1 _15875_/X sky130_fd_sc_hd__buf_1
X_18663_ _18078_/Y _20462_/Q _18906_/S vssd1 vssd1 vccd1 vccd1 _18663_/X sky130_fd_sc_hd__mux2_1
XFILLER_91_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17614_ _19346_/Q vssd1 vssd1 vccd1 vccd1 _17614_/Y sky130_fd_sc_hd__inv_2
X_14826_ _20106_/Q vssd1 vssd1 vccd1 vccd1 _14883_/A sky130_fd_sc_hd__inv_2
X_18594_ _17079_/Y _12083_/Y _18884_/S vssd1 vssd1 vccd1 vccd1 _18594_/X sky130_fd_sc_hd__mux2_1
XFILLER_240_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14757_ _14757_/A vssd1 vssd1 vccd1 vccd1 _14758_/B sky130_fd_sc_hd__buf_1
X_17545_ _17545_/A _17807_/B vssd1 vssd1 vccd1 vccd1 _17545_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__13281__B1 _13280_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11969_ _13179_/B vssd1 vssd1 vccd1 vccd1 _13717_/B sky130_fd_sc_hd__buf_1
XFILLER_220_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13708_ _13708_/A vssd1 vssd1 vccd1 vccd1 _13708_/X sky130_fd_sc_hd__buf_1
X_17476_ _18800_/X _17315_/X _18768_/X _17844_/A vssd1 vssd1 vccd1 vccd1 _17476_/X
+ sky130_fd_sc_hd__o22a_2
X_14688_ _14692_/A vssd1 vssd1 vccd1 vccd1 _14688_/X sky130_fd_sc_hd__buf_1
XFILLER_189_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19215_ _17678_/Y _17679_/Y _17680_/Y _17681_/Y _19275_/S0 _21004_/Q vssd1 vssd1
+ vccd1 vccd1 _19215_/X sky130_fd_sc_hd__mux4_1
XANTENNA__13033__B1 _13032_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16427_ _16427_/A vssd1 vssd1 vccd1 vccd1 _16427_/X sky130_fd_sc_hd__buf_1
X_13639_ _13651_/A vssd1 vssd1 vccd1 vccd1 _13639_/X sky130_fd_sc_hd__buf_1
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16358_ _19888_/D vssd1 vssd1 vccd1 vccd1 _17072_/B sky130_fd_sc_hd__buf_1
X_19146_ _19142_/X _19143_/X _19144_/X _19145_/X _21018_/Q _21019_/Q vssd1 vssd1 vccd1
+ vccd1 _19146_/X sky130_fd_sc_hd__mux4_2
XFILLER_173_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19996__RESET_B repeater220/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15309_ _20037_/Q _15302_/A _19867_/Q _15305_/X vssd1 vssd1 vccd1 vccd1 _20037_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_117_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16522__A1 _16495_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19077_ _16726_/X _20898_/Q _19908_/D vssd1 vssd1 vccd1 vccd1 _19077_/X sky130_fd_sc_hd__mux2_1
X_16289_ _16289_/A vssd1 vssd1 vccd1 vccd1 _16289_/X sky130_fd_sc_hd__buf_1
XANTENNA__19925__RESET_B repeater211/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19147__S0 _19285_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18028_ _18033_/A vssd1 vssd1 vccd1 vccd1 _18032_/B sky130_fd_sc_hd__buf_4
XFILLER_161_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09801_ _16620_/A _16620_/C _09806_/B _09716_/D _09800_/Y vssd1 vssd1 vccd1 vccd1
+ _09802_/A sky130_fd_sc_hd__o32a_1
XANTENNA__09960__B1 _09693_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19979_ _20809_/CLK _19979_/D repeater270/X vssd1 vssd1 vccd1 vccd1 _19979_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_115_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11736__A _13166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09732_ _21234_/Q _20154_/Q _11059_/A _09731_/Y vssd1 vssd1 vccd1 vccd1 _09732_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__20412__RESET_B repeater184/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09663_ _13311_/A vssd1 vssd1 vccd1 vccd1 _09663_/X sky130_fd_sc_hd__buf_6
XFILLER_227_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09594_ _20890_/Q vssd1 vssd1 vccd1 vccd1 _13047_/A sky130_fd_sc_hd__inv_2
XFILLER_227_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20823_ _20841_/CLK _20823_/D repeater251/X vssd1 vssd1 vccd1 vccd1 _20823_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18953__S _18962_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12567__A _20891_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_opt_4_HCLK_A clkbuf_opt_4_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20754_ _21477_/CLK _20754_/D repeater201/X vssd1 vssd1 vccd1 vccd1 _20754_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13024__B1 _12855_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20685_ _21302_/CLK _20685_/D repeater208/X vssd1 vssd1 vccd1 vccd1 _20685_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19138__S0 _19285_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21306_ _21306_/CLK _21306_/D repeater206/X vssd1 vssd1 vccd1 vccd1 _21306_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_108_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21237_ _21239_/CLK _21237_/D repeater249/X vssd1 vssd1 vccd1 vccd1 _21237_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_105_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21168_ _21184_/CLK _21168_/D repeater220/X vssd1 vssd1 vccd1 vccd1 _21168_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_131_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20119_ _21452_/CLK _20119_/D repeater247/X vssd1 vssd1 vccd1 vccd1 _20119_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_77_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12838__B1 _09621_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21099_ _21429_/CLK _21099_/D repeater231/X vssd1 vssd1 vccd1 vccd1 _21099_/Q sky130_fd_sc_hd__dfrtp_1
X_13990_ _13990_/A vssd1 vssd1 vccd1 vccd1 _14004_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_219_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09703__B1 _09702_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_219_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12941_ _20715_/Q _12935_/X _12857_/X _12937_/X vssd1 vssd1 vccd1 vccd1 _20715_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_234_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19024__S _19026_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15660_ _19693_/Q _15656_/X _15657_/X _15659_/X vssd1 vssd1 vccd1 vccd1 _19693_/D
+ sky130_fd_sc_hd__a22o_1
X_12872_ _13163_/A vssd1 vssd1 vccd1 vccd1 _12872_/X sky130_fd_sc_hd__buf_2
XPHY_4220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14611_ _20201_/Q _14609_/Y _14610_/X _14591_/B vssd1 vssd1 vccd1 vccd1 _20201_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_4253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11823_ _21038_/Q _11822_/Y _11818_/Y vssd1 vssd1 vccd1 vccd1 _21038_/D sky130_fd_sc_hd__o21ba_1
XPHY_4264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15591_ _19727_/Q _15584_/X _15590_/X _15586_/X vssd1 vssd1 vccd1 vccd1 _19727_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_199_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18863__S _18928_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21359__RESET_B repeater254/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17330_ _19496_/Q vssd1 vssd1 vccd1 vccd1 _17330_/Y sky130_fd_sc_hd__inv_2
XPHY_4297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14542_ _20136_/Q vssd1 vssd1 vccd1 vccd1 _14557_/A sky130_fd_sc_hd__inv_2
X_11754_ _21054_/Q vssd1 vssd1 vccd1 vccd1 _11754_/Y sky130_fd_sc_hd__inv_2
XPHY_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10705_ _10705_/A _10715_/A vssd1 vssd1 vccd1 vccd1 _10706_/B sky130_fd_sc_hd__or2_2
XFILLER_159_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17261_ _19623_/Q vssd1 vssd1 vccd1 vccd1 _17261_/Y sky130_fd_sc_hd__inv_2
X_14473_ _20234_/Q _14471_/Y _14472_/X _14378_/B vssd1 vssd1 vccd1 vccd1 _20234_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_187_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13015__B1 _12928_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11685_ _21086_/Q _11679_/X _11684_/X _11682_/X vssd1 vssd1 vccd1 vccd1 _21086_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19000_ _17000_/X _20423_/Q _19019_/S vssd1 vssd1 vccd1 vccd1 _19976_/D sky130_fd_sc_hd__mux2_1
X_16212_ _21447_/Q vssd1 vssd1 vccd1 vccd1 _16212_/X sky130_fd_sc_hd__buf_1
X_13424_ input42/X vssd1 vssd1 vccd1 vccd1 _13424_/X sky130_fd_sc_hd__clkbuf_2
X_10636_ _21325_/Q _10635_/Y _10577_/Y _20769_/Q vssd1 vssd1 vccd1 vccd1 _10636_/X
+ sky130_fd_sc_hd__o22a_1
X_17192_ _21242_/Q vssd1 vssd1 vccd1 vccd1 _17192_/Y sky130_fd_sc_hd__inv_2
X_16143_ _16143_/A vssd1 vssd1 vccd1 vccd1 _16143_/X sky130_fd_sc_hd__buf_1
XFILLER_10_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13355_ _20515_/Q _13351_/X _13221_/X _13352_/X vssd1 vssd1 vccd1 vccd1 _20515_/D
+ sky130_fd_sc_hd__a22o_1
X_10567_ _21333_/Q vssd1 vssd1 vccd1 vccd1 _10662_/A sky130_fd_sc_hd__inv_2
XANTENNA__19129__S0 _19285_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12306_ _12306_/A _12306_/B vssd1 vssd1 vccd1 vccd1 _12386_/A sky130_fd_sc_hd__or2_1
X_16074_ _19496_/Q _16071_/X _15772_/X _16072_/X vssd1 vssd1 vccd1 vccd1 _19496_/D
+ sky130_fd_sc_hd__a22o_1
X_13286_ _13293_/A vssd1 vssd1 vccd1 vccd1 _13286_/X sky130_fd_sc_hd__buf_1
X_10498_ _21280_/Q vssd1 vssd1 vccd1 vccd1 _10757_/A sky130_fd_sc_hd__inv_2
XFILLER_143_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19902_ _21185_/CLK _19902_/D repeater223/X vssd1 vssd1 vccd1 vccd1 _19902_/Q sky130_fd_sc_hd__dfrtp_1
X_15025_ _15025_/A _15025_/B _15025_/C vssd1 vssd1 vccd1 vccd1 _20077_/D sky130_fd_sc_hd__nor3_1
XFILLER_216_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12237_ _12475_/A _20507_/Q _20927_/Q _12236_/Y vssd1 vssd1 vccd1 vccd1 _12237_/X
+ sky130_fd_sc_hd__o22a_1
X_19833_ _19834_/CLK _19833_/D vssd1 vssd1 vccd1 vccd1 _19833_/Q sky130_fd_sc_hd__dfxtp_1
X_12168_ _20362_/Q vssd1 vssd1 vccd1 vccd1 _12168_/Y sky130_fd_sc_hd__inv_2
XFILLER_150_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11119_ _11076_/X _09739_/X _11100_/X _11118_/X vssd1 vssd1 vccd1 vccd1 _21226_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_84_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19764_ _19765_/CLK _19764_/D vssd1 vssd1 vccd1 vccd1 _19764_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16976_ _19971_/Q _16970_/A _16965_/A _16975_/Y _16972_/Y vssd1 vssd1 vccd1 vccd1
+ _16977_/B sky130_fd_sc_hd__o32a_1
X_12099_ _20958_/Q _20372_/Q _12097_/X _17806_/A vssd1 vssd1 vccd1 vccd1 _12103_/C
+ sky130_fd_sc_hd__o22a_1
XFILLER_232_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18715_ _18714_/X _10265_/A _18841_/S vssd1 vssd1 vccd1 vccd1 _18715_/X sky130_fd_sc_hd__mux2_1
Xinput6 HADDR[14] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_1
X_15927_ _15927_/A vssd1 vssd1 vccd1 vccd1 _15927_/X sky130_fd_sc_hd__buf_1
X_19695_ _19776_/CLK _19695_/D vssd1 vssd1 vccd1 vccd1 _19695_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_209_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18646_ _18085_/Y _17007_/Y _18875_/S vssd1 vssd1 vccd1 vccd1 _18646_/X sky130_fd_sc_hd__mux2_1
XFILLER_92_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15858_ _19601_/Q _15856_/X _15788_/X _15857_/X vssd1 vssd1 vccd1 vccd1 _19601_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_36_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16440__B1 _16332_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14809_ _20119_/Q _14311_/X _14794_/A _14808_/X vssd1 vssd1 vccd1 vccd1 _20119_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_17_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18577_ _18848_/A0 _17850_/Y _18666_/S vssd1 vssd1 vccd1 vccd1 _18577_/X sky130_fd_sc_hd__mux2_1
XANTENNA__18773__S _18841_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15789_ _15789_/A vssd1 vssd1 vccd1 vccd1 _15789_/X sky130_fd_sc_hd__buf_1
XFILLER_178_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17528_ _20120_/Q _17446_/A _17368_/X _17526_/Y vssd1 vssd1 vccd1 vccd1 _17528_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17897__B _17898_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21029__RESET_B repeater242/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17459_ _17457_/Y _17292_/A _17458_/Y _17381_/X vssd1 vssd1 vccd1 vccd1 _17459_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_20_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09696__A input49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20470_ _20470_/CLK _20470_/D repeater279/X vssd1 vssd1 vccd1 vccd1 _20470_/Q sky130_fd_sc_hd__dfrtp_1
X_19129_ _19686_/Q _19374_/Q _19670_/Q _19662_/Q _19285_/S0 _21017_/Q vssd1 vssd1
+ vccd1 vccd1 _19129_/X sky130_fd_sc_hd__mux4_1
XFILLER_145_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13309__A1 _20541_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21022_ _21223_/CLK _21022_/D repeater238/X vssd1 vssd1 vccd1 vccd1 _21022_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__14809__A1 _20119_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09715_ _21457_/Q vssd1 vssd1 vccd1 vccd1 _09716_/D sky130_fd_sc_hd__inv_2
XFILLER_19_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_80_HCLK clkbuf_opt_7_HCLK/A vssd1 vssd1 vccd1 vccd1 _21483_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_216_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17153__A _17153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09646_ _09660_/A vssd1 vssd1 vccd1 vccd1 _09646_/X sky130_fd_sc_hd__buf_1
XFILLER_71_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19665__CLK _19765_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18683__S _18884_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21452__RESET_B repeater247/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20806_ _21011_/CLK _20806_/D repeater235/X vssd1 vssd1 vccd1 vccd1 _20806_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20737_ _21342_/CLK _20737_/D repeater211/X vssd1 vssd1 vccd1 vccd1 _20737_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11470_ _19095_/X _11468_/X _21163_/Q _11469_/X vssd1 vssd1 vccd1 vccd1 _21163_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_183_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20668_ _21306_/CLK _20668_/D repeater207/X vssd1 vssd1 vccd1 vccd1 _20668_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10421_ _20698_/Q vssd1 vssd1 vccd1 vccd1 _10421_/Y sky130_fd_sc_hd__inv_2
X_20599_ _20693_/CLK _20599_/D repeater196/X vssd1 vssd1 vccd1 vccd1 _20599_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_136_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13140_ input44/X vssd1 vssd1 vccd1 vccd1 _13140_/X sky130_fd_sc_hd__clkbuf_4
X_10352_ _20728_/Q vssd1 vssd1 vccd1 vccd1 _10352_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19019__S _19019_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13071_ _20654_/Q _13066_/X _12922_/X _13067_/X vssd1 vssd1 vccd1 vccd1 _20654_/D
+ sky130_fd_sc_hd__a22o_1
X_10283_ _10283_/A _10283_/B vssd1 vssd1 vccd1 vccd1 _10377_/A sky130_fd_sc_hd__or2_1
X_12022_ _19074_/X _12017_/X _20991_/Q _12018_/X vssd1 vssd1 vccd1 vccd1 _20991_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_input49_A HWDATA[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16830_ _16830_/A _16830_/B vssd1 vssd1 vccd1 vccd1 _16830_/Y sky130_fd_sc_hd__nor2_1
X_16761_ _19920_/Q _16756_/A _19921_/Q vssd1 vssd1 vccd1 vccd1 _16761_/X sky130_fd_sc_hd__o21a_1
X_13973_ _13972_/X _20307_/Q _20306_/Q _20308_/Q vssd1 vssd1 vccd1 vccd1 _13973_/X
+ sky130_fd_sc_hd__and4b_1
XFILLER_234_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18500_ _18499_/X _17875_/Y _18666_/S vssd1 vssd1 vccd1 vccd1 _18500_/X sky130_fd_sc_hd__mux2_1
X_15712_ _19669_/Q _15709_/X _15657_/X _15711_/X vssd1 vssd1 vccd1 vccd1 _19669_/D
+ sky130_fd_sc_hd__a22o_1
X_12924_ _12924_/A vssd1 vssd1 vccd1 vccd1 _12924_/X sky130_fd_sc_hd__buf_1
XFILLER_206_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16692_ _19890_/Q _19891_/Q _14232_/B vssd1 vssd1 vccd1 vccd1 _16692_/X sky130_fd_sc_hd__a21bo_1
X_19480_ _19961_/CLK _19480_/D vssd1 vssd1 vccd1 vccd1 _19480_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_234_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18431_ _18430_/X _10274_/A _18841_/S vssd1 vssd1 vccd1 vccd1 _18431_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13236__B1 _13154_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15643_ _19701_/Q _15640_/X _15469_/X _15642_/X vssd1 vssd1 vccd1 vccd1 _19701_/D
+ sky130_fd_sc_hd__a22o_1
X_12855_ _12855_/A vssd1 vssd1 vccd1 vccd1 _12855_/X sky130_fd_sc_hd__clkbuf_2
XPHY_4050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18593__S _18880_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_repeater188_A repeater270/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11806_ _11806_/A _11855_/A vssd1 vssd1 vccd1 vccd1 _11850_/A sky130_fd_sc_hd__or2_1
X_18362_ _17281_/X _18044_/Y _18787_/S vssd1 vssd1 vccd1 vccd1 _18362_/X sky130_fd_sc_hd__mux2_1
X_15574_ _15574_/A _20125_/Q _15574_/C vssd1 vssd1 vccd1 vccd1 _16451_/C sky130_fd_sc_hd__or3_4
XFILLER_92_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12786_ _12804_/A vssd1 vssd1 vccd1 vccd1 _12786_/X sky130_fd_sc_hd__buf_1
XFILLER_187_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14525_ _14518_/A _14518_/B _20209_/Q _14464_/X _14458_/X vssd1 vssd1 vccd1 vccd1
+ _20209_/D sky130_fd_sc_hd__o221a_1
XPHY_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17313_ _17573_/A vssd1 vssd1 vccd1 vccd1 _17861_/A sky130_fd_sc_hd__clkbuf_2
XPHY_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11737_ _11737_/A vssd1 vssd1 vccd1 vccd1 _11737_/X sky130_fd_sc_hd__buf_1
XFILLER_14_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18293_ _17977_/Y _20654_/Q _18903_/S vssd1 vssd1 vccd1 vccd1 _18293_/X sky130_fd_sc_hd__mux2_1
XFILLER_230_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14456_ _14488_/A vssd1 vssd1 vccd1 vccd1 _14524_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA__14736__B1 _13710_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17244_ _19519_/Q vssd1 vssd1 vccd1 vccd1 _17244_/Y sky130_fd_sc_hd__inv_2
XPHY_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11668_ _16654_/A _11657_/A _11665_/Y _11509_/Y _11676_/S vssd1 vssd1 vccd1 vccd1
+ _11669_/A sky130_fd_sc_hd__o32a_1
XPHY_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13407_ _20487_/Q _13404_/X _13209_/X _13405_/X vssd1 vssd1 vccd1 vccd1 _20487_/D
+ sky130_fd_sc_hd__a22o_1
X_17175_ _17177_/A _17175_/B vssd1 vssd1 vccd1 vccd1 _18880_/S sky130_fd_sc_hd__nor2_8
X_10619_ _20752_/Q vssd1 vssd1 vccd1 vccd1 _10619_/Y sky130_fd_sc_hd__inv_2
XPHY_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14387_ _20030_/Q vssd1 vssd1 vccd1 vccd1 _14387_/Y sky130_fd_sc_hd__inv_2
XFILLER_155_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11599_ _11599_/A vssd1 vssd1 vccd1 vccd1 _11605_/A sky130_fd_sc_hd__inv_2
XFILLER_227_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16126_ _19471_/Q _16119_/X _16125_/X _16121_/X vssd1 vssd1 vccd1 vccd1 _19471_/D
+ sky130_fd_sc_hd__a22o_1
X_13338_ _20526_/Q _13331_/X _13274_/X _13334_/X vssd1 vssd1 vccd1 vccd1 _20526_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_182_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16057_ _16057_/A vssd1 vssd1 vccd1 vccd1 _16057_/X sky130_fd_sc_hd__buf_1
XANTENNA__12670__A input54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13269_ _20561_/Q _13264_/X _13265_/X _13268_/X vssd1 vssd1 vccd1 vccd1 _20561_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_142_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20075__RESET_B repeater276/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15008_ _15006_/A _15006_/B _15006_/Y _14989_/X vssd1 vssd1 vccd1 vccd1 _20086_/D
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__18768__S _18875_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19816_ _20172_/CLK _19816_/D vssd1 vssd1 vccd1 vccd1 _19816_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_243_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19747_ _19765_/CLK _19747_/D vssd1 vssd1 vccd1 vccd1 _19747_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16959_ _16963_/B vssd1 vssd1 vccd1 vccd1 _16966_/B sky130_fd_sc_hd__inv_2
XFILLER_37_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14672__C1 _11800_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_237_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19678_ _19811_/CLK _19678_/D vssd1 vssd1 vccd1 vccd1 _19678_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18629_ _18628_/X _12168_/Y _18909_/S vssd1 vssd1 vccd1 vccd1 _18629_/X sky130_fd_sc_hd__mux2_1
XFILLER_213_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13006__A input53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_240_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18166__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_212_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20522_ _20944_/CLK _20522_/D repeater277/X vssd1 vssd1 vccd1 vccd1 _20522_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__14727__B1 _13712_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20845__RESET_B repeater243/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20453_ _20476_/CLK _20453_/D repeater280/X vssd1 vssd1 vccd1 vccd1 _20453_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_192_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20384_ _20972_/CLK _20384_/D repeater280/X vssd1 vssd1 vccd1 vccd1 _20384_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_107_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_114_HCLK_A clkbuf_opt_3_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput140 _21043_/Q vssd1 vssd1 vccd1 vccd1 scl_oen_o_S4 sky130_fd_sc_hd__clkbuf_2
XANTENNA__12580__A _12580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_217_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18678__S _18926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15891__A _16235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21005_ _21009_/CLK _21005_/D repeater235/X vssd1 vssd1 vccd1 vccd1 _21005_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_87_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10970_ _10931_/X _10970_/B _10970_/C _10970_/D vssd1 vssd1 vccd1 vccd1 _11800_/A
+ sky130_fd_sc_hd__and4b_4
XFILLER_55_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09629_ _21483_/Q _09620_/X _09628_/X _09624_/X vssd1 vssd1 vccd1 vccd1 _21483_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_55_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13218__B1 _13216_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12640_ input26/X _12637_/X _20846_/Q _12638_/X vssd1 vssd1 vccd1 vccd1 _20846_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_43_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12571_ _17169_/A _12566_/X _18217_/X _18242_/S vssd1 vssd1 vccd1 vccd1 _20891_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_23_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12755__A _17083_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_212_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14310_ _14792_/A _16481_/B vssd1 vssd1 vccd1 vccd1 _14796_/A sky130_fd_sc_hd__nand2_2
XFILLER_12_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11522_ _11522_/A vssd1 vssd1 vccd1 vccd1 _21145_/D sky130_fd_sc_hd__inv_2
XPHY_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_opt_5_HCLK clkbuf_opt_7_HCLK/A vssd1 vssd1 vccd1 vccd1 _19904_/CLK sky130_fd_sc_hd__clkbuf_16
X_15290_ _19856_/Q _15290_/B vssd1 vssd1 vccd1 vccd1 _15291_/B sky130_fd_sc_hd__or2_1
XPHY_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14241_ _19901_/Q _14241_/B vssd1 vssd1 vccd1 vccd1 _14242_/B sky130_fd_sc_hd__or2_1
XFILLER_7_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11453_ _21165_/Q _11453_/B vssd1 vssd1 vccd1 vccd1 _11454_/B sky130_fd_sc_hd__or2_1
XFILLER_11_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15391__B1 _15346_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10404_ _10346_/X _10406_/A _10269_/A vssd1 vssd1 vccd1 vccd1 _10405_/C sky130_fd_sc_hd__o21a_1
XANTENNA__13941__A1 _20637_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14172_ _14176_/A vssd1 vssd1 vccd1 vccd1 _14205_/A sky130_fd_sc_hd__inv_2
X_11384_ _11385_/A _11384_/B _11384_/C vssd1 vssd1 vccd1 vccd1 _11786_/A sky130_fd_sc_hd__nor3_4
XFILLER_194_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13123_ _20625_/Q _13120_/X _12999_/X _13121_/X vssd1 vssd1 vccd1 vccd1 _20625_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13586__A input68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17058__A _21042_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10335_ _21370_/Q _10333_/Y _10260_/A _20703_/Q _10334_/X vssd1 vssd1 vccd1 vccd1
+ _10340_/C sky130_fd_sc_hd__o221a_1
X_18980_ _21426_/Q _21099_/Q _18983_/S vssd1 vssd1 vccd1 vccd1 _18980_/X sky130_fd_sc_hd__mux2_1
XFILLER_180_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20538__CLK _20592_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17931_ _18024_/A vssd1 vssd1 vccd1 vccd1 _17931_/X sky130_fd_sc_hd__buf_1
XFILLER_112_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13054_ _13080_/A vssd1 vssd1 vccd1 vccd1 _13073_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_78_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10266_ _10266_/A _10266_/B vssd1 vssd1 vccd1 vccd1 _10409_/A sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_36_HCLK_A _20004_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18588__S _18908_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12005_ _19888_/Q vssd1 vssd1 vccd1 vccd1 _12006_/C sky130_fd_sc_hd__inv_2
XFILLER_79_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_99_HCLK_A clkbuf_4_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17862_ _17862_/A vssd1 vssd1 vccd1 vccd1 _17862_/X sky130_fd_sc_hd__buf_1
XFILLER_39_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10197_ _21389_/Q _10196_/Y _10166_/A _10151_/B vssd1 vssd1 vccd1 vccd1 _21389_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_120_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19601_ _21021_/CLK _19601_/D vssd1 vssd1 vccd1 vccd1 _19601_/Q sky130_fd_sc_hd__dfxtp_1
X_16813_ _19934_/Q _16813_/B vssd1 vssd1 vccd1 vccd1 _16822_/C sky130_fd_sc_hd__or2_2
XFILLER_238_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17793_ _19878_/Q vssd1 vssd1 vccd1 vccd1 _17793_/Y sky130_fd_sc_hd__inv_2
XFILLER_213_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21374__RESET_B repeater257/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19532_ _21462_/CLK _19532_/D vssd1 vssd1 vccd1 vccd1 _19532_/Q sky130_fd_sc_hd__dfxtp_1
X_16744_ _16744_/A _16744_/B vssd1 vssd1 vccd1 vccd1 _19913_/D sky130_fd_sc_hd__nor2_1
XANTENNA__18396__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13956_ _20649_/Q _13882_/A _13954_/Y _20306_/Q _13955_/Y vssd1 vssd1 vccd1 vccd1
+ _13961_/C sky130_fd_sc_hd__o221a_1
XANTENNA__21303__RESET_B repeater207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19463_ _21234_/CLK _19463_/D vssd1 vssd1 vccd1 vccd1 _19463_/Q sky130_fd_sc_hd__dfxtp_1
X_12907_ _20732_/Q _12901_/X _12658_/X _12904_/X vssd1 vssd1 vccd1 vccd1 _20732_/D
+ sky130_fd_sc_hd__a22o_1
X_16675_ _21163_/Q _11451_/B _11452_/B vssd1 vssd1 vccd1 vccd1 _16675_/X sky130_fd_sc_hd__a21bo_1
X_13887_ _13971_/B _13887_/B vssd1 vssd1 vccd1 vccd1 _13993_/A sky130_fd_sc_hd__or2_1
X_18414_ _17281_/X _17885_/Y _18835_/S vssd1 vssd1 vccd1 vccd1 _18414_/X sky130_fd_sc_hd__mux2_1
X_12838_ _20760_/Q _12835_/X _09621_/X _12836_/X vssd1 vssd1 vccd1 vccd1 _20760_/D
+ sky130_fd_sc_hd__a22o_1
X_15626_ _15632_/A vssd1 vssd1 vccd1 vccd1 _15633_/A sky130_fd_sc_hd__inv_2
XFILLER_22_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19394_ _21001_/CLK _19394_/D vssd1 vssd1 vccd1 vccd1 _19394_/Q sky130_fd_sc_hd__dfxtp_1
X_18345_ _17079_/Y _12054_/Y _18908_/S vssd1 vssd1 vccd1 vccd1 _18345_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15557_ _19743_/Q _15553_/X _15524_/X _15554_/X vssd1 vssd1 vccd1 vccd1 _19743_/D
+ sky130_fd_sc_hd__a22o_1
X_12769_ _20798_/Q _12765_/X _12668_/X _12766_/X vssd1 vssd1 vccd1 vccd1 _20798_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_230_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14508_ _20218_/Q _14507_/Y _14504_/B _14477_/X vssd1 vssd1 vccd1 vccd1 _20218_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_202_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14709__B1 _12855_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_1_0_HCLK_A clkbuf_2_1_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18276_ _19171_/X _21271_/Q _18281_/S vssd1 vssd1 vccd1 vccd1 _18276_/X sky130_fd_sc_hd__mux2_1
X_15488_ _19774_/Q _15479_/X _15487_/X _15481_/X vssd1 vssd1 vccd1 vccd1 _19774_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_174_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput20 HADDR[27] vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__buf_1
X_17227_ _17853_/A vssd1 vssd1 vccd1 vccd1 _17227_/X sky130_fd_sc_hd__buf_1
X_14439_ _21481_/Q vssd1 vssd1 vccd1 vccd1 _14439_/Y sky130_fd_sc_hd__inv_2
Xinput31 HADDR[8] vssd1 vssd1 vccd1 vccd1 input31/X sky130_fd_sc_hd__clkbuf_1
XFILLER_175_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput42 HWDATA[13] vssd1 vssd1 vccd1 vccd1 input42/X sky130_fd_sc_hd__buf_2
Xinput53 HWDATA[23] vssd1 vssd1 vccd1 vccd1 input53/X sky130_fd_sc_hd__clkbuf_4
Xinput64 HWDATA[4] vssd1 vssd1 vccd1 vccd1 input64/X sky130_fd_sc_hd__buf_6
Xinput75 scl_i_S4 vssd1 vssd1 vccd1 vccd1 input75/X sky130_fd_sc_hd__clkbuf_1
X_17158_ _17548_/A vssd1 vssd1 vccd1 vccd1 _17158_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_7_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16109_ _20331_/Q vssd1 vssd1 vccd1 vccd1 _16109_/X sky130_fd_sc_hd__clkbuf_2
X_17089_ _21343_/Q _20700_/Q vssd1 vssd1 vccd1 vccd1 _17089_/X sky130_fd_sc_hd__and2_2
X_09980_ _21414_/Q _09975_/X _09693_/X _09976_/X vssd1 vssd1 vccd1 vccd1 _21414_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_131_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13696__B1 _12863_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18498__S _18910_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13448__B1 _13446_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18387__A0 _17079_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_1_HCLK clkbuf_1_0_1_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_226_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10682__B1 _10677_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_241_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18139__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_110_HCLK clkbuf_opt_3_HCLK/A vssd1 vssd1 vccd1 vccd1 _20070_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_80_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18961__S _18962_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20505_ _20930_/CLK _20505_/D repeater268/X vssd1 vssd1 vccd1 vccd1 _20505_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12725__D _13383_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21485_ _21485_/CLK _21485_/D repeater200/X vssd1 vssd1 vccd1 vccd1 _21485_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_146_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20436_ _20937_/CLK _20436_/D repeater278/X vssd1 vssd1 vccd1 vccd1 _20436_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_106_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17665__A2 _17646_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20367_ _20951_/CLK _20367_/D repeater271/X vssd1 vssd1 vccd1 vccd1 _20367_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_122_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10120_ _10077_/A _10119_/Y _21406_/Q _20803_/Q vssd1 vssd1 vccd1 vccd1 _10120_/X
+ sky130_fd_sc_hd__a22o_1
X_20298_ _20316_/CLK _20298_/D repeater197/X vssd1 vssd1 vccd1 vccd1 _20298_/Q sky130_fd_sc_hd__dfrtp_1
X_10051_ _21386_/Q vssd1 vssd1 vccd1 vccd1 _10207_/A sky130_fd_sc_hd__inv_2
XANTENNA__18201__S _18680_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13439__B1 _13243_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13810_ _20609_/Q _14575_/A _17542_/A _20180_/Q _13809_/X vssd1 vssd1 vccd1 vccd1
+ _13811_/D sky130_fd_sc_hd__o221a_1
XFILLER_180_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14790_ _14783_/A _14288_/X _19126_/X _20121_/Q vssd1 vssd1 vccd1 vccd1 _20121_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_63_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13741_ _17810_/A _20184_/Q _17941_/A _20193_/Q vssd1 vssd1 vccd1 vccd1 _13741_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_44_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10953_ _21031_/Q vssd1 vssd1 vccd1 vccd1 _11848_/A sky130_fd_sc_hd__buf_1
XANTENNA__19862__RESET_B repeater226/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_216_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19032__S _19046_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13672_ _20356_/Q _13667_/X _13557_/X _13668_/X vssd1 vssd1 vccd1 vccd1 _20356_/D
+ sky130_fd_sc_hd__a22o_1
X_16460_ _16460_/A vssd1 vssd1 vccd1 vccd1 _16460_/X sky130_fd_sc_hd__buf_1
X_10884_ _12544_/A vssd1 vssd1 vccd1 vccd1 _10884_/X sky130_fd_sc_hd__buf_2
XFILLER_188_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12623_ input6/X _12619_/X _20857_/Q _12620_/X vssd1 vssd1 vccd1 vccd1 _20857_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_71_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15411_ _21015_/Q vssd1 vssd1 vccd1 vccd1 _15673_/A sky130_fd_sc_hd__buf_1
X_16391_ _16433_/A _16485_/A vssd1 vssd1 vccd1 vccd1 _16399_/A sky130_fd_sc_hd__or2_2
XANTENNA__17060__B _17060_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10589__A2_N _20760_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13611__B1 _13545_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18871__S _18899_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15342_ _19835_/Q _15337_/X _14264_/X _15339_/X vssd1 vssd1 vccd1 vccd1 _19835_/D
+ sky130_fd_sc_hd__a22o_1
X_18130_ _18129_/X _12291_/Y _18910_/S vssd1 vssd1 vccd1 vccd1 _18130_/X sky130_fd_sc_hd__mux2_1
XPHY_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12554_ _12554_/A vssd1 vssd1 vccd1 vccd1 _12554_/X sky130_fd_sc_hd__buf_1
XFILLER_196_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18550__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11505_ _11504_/X _11487_/X _19111_/S _11500_/Y _21149_/Q vssd1 vssd1 vccd1 vccd1
+ _21149_/D sky130_fd_sc_hd__a32o_1
XPHY_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15273_ _15269_/Y _20059_/Q _15270_/Y _20049_/Q _15272_/X vssd1 vssd1 vccd1 vccd1
+ _15284_/A sky130_fd_sc_hd__o221a_1
X_18061_ _20424_/Q vssd1 vssd1 vccd1 vccd1 _18061_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15364__B1 _14264_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12485_ _12472_/A _12472_/B _12483_/Y _12445_/X vssd1 vssd1 vccd1 vccd1 _20924_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_156_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17012_ _19980_/Q _17008_/A _17011_/Y _17008_/Y vssd1 vssd1 vccd1 vccd1 _17013_/B
+ sky130_fd_sc_hd__o22a_1
X_14224_ _14074_/A _14074_/B _14222_/Y _14185_/X vssd1 vssd1 vccd1 vccd1 _20263_/D
+ sky130_fd_sc_hd__a211oi_4
X_11436_ _11385_/A _11420_/A _11786_/A _11421_/X vssd1 vssd1 vccd1 vccd1 _21169_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_171_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11925__B1 _21006_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14155_ _14155_/A _14155_/B _14155_/C _14155_/D vssd1 vssd1 vccd1 vccd1 _14171_/C
+ sky130_fd_sc_hd__and4_1
X_11367_ _21184_/Q _11367_/B _11379_/C vssd1 vssd1 vccd1 vccd1 _11387_/B sky130_fd_sc_hd__or3_4
XFILLER_113_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13106_ _13108_/A _13106_/B vssd1 vssd1 vccd1 vccd1 _13107_/S sky130_fd_sc_hd__or2_1
X_10318_ _21372_/Q _10317_/Y _10287_/A _20731_/Q vssd1 vssd1 vccd1 vccd1 _10318_/X
+ sky130_fd_sc_hd__o22a_1
X_18963_ _16620_/X _16619_/Y _18976_/S vssd1 vssd1 vccd1 vccd1 _18963_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14086_ _14086_/A _14201_/A vssd1 vssd1 vccd1 vccd1 _14087_/B sky130_fd_sc_hd__or2_1
XFILLER_113_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11298_ _11311_/B _11306_/B _11311_/A vssd1 vssd1 vccd1 vccd1 _11301_/A sky130_fd_sc_hd__or3b_1
XFILLER_239_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_160_HCLK_A clkbuf_opt_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_224_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18605__A1 _14403_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13037_ _20672_/Q _13034_/X _12954_/X _13035_/X vssd1 vssd1 vccd1 vccd1 _20672_/D
+ sky130_fd_sc_hd__a22o_1
X_17914_ _18416_/X _17227_/X _18426_/X _17817_/X vssd1 vssd1 vccd1 vccd1 _17914_/X
+ sky130_fd_sc_hd__o22a_1
X_10249_ _21354_/Q vssd1 vssd1 vccd1 vccd1 _10269_/A sky130_fd_sc_hd__inv_2
X_18894_ _18893_/X _13735_/Y _18910_/S vssd1 vssd1 vccd1 vccd1 _18894_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17845_ _18614_/X _17324_/X _18612_/X _18064_/A vssd1 vssd1 vccd1 vccd1 _17845_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_121_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17776_ _21438_/Q _17776_/B vssd1 vssd1 vccd1 vccd1 _17776_/Y sky130_fd_sc_hd__nand2_1
XFILLER_240_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14988_ _20093_/Q _14987_/Y _14872_/B _14978_/X vssd1 vssd1 vccd1 vccd1 _20093_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_208_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19515_ _21462_/CLK _19515_/D vssd1 vssd1 vccd1 vccd1 _19515_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_133_HCLK clkbuf_4_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20930_/CLK sky130_fd_sc_hd__clkbuf_16
X_16727_ _20989_/Q _11995_/B _11996_/B vssd1 vssd1 vccd1 vccd1 _16727_/X sky130_fd_sc_hd__a21bo_1
X_13939_ _20640_/Q vssd1 vssd1 vccd1 vccd1 _13939_/Y sky130_fd_sc_hd__inv_2
XFILLER_223_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19446_ _20137_/CLK _19446_/D vssd1 vssd1 vccd1 vccd1 _19446_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16658_ _19863_/Q _15297_/B _15298_/B vssd1 vssd1 vccd1 vccd1 _16658_/X sky130_fd_sc_hd__a21bo_1
XFILLER_34_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13602__A0 _13600_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15609_ _15609_/A _15609_/B _16616_/B vssd1 vssd1 vccd1 vccd1 _16344_/C sky130_fd_sc_hd__or3_4
X_19377_ _19706_/CLK _19377_/D vssd1 vssd1 vccd1 vccd1 _19377_/Q sky130_fd_sc_hd__dfxtp_1
X_16589_ _16740_/A _16535_/X _19992_/Q _16588_/Y vssd1 vssd1 vccd1 vccd1 _19992_/D
+ sky130_fd_sc_hd__a31o_1
XANTENNA__18781__S _18849_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18328_ _18327_/X _21352_/Q _18841_/S vssd1 vssd1 vccd1 vccd1 _18328_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18259_ _17079_/Y _12048_/Y _18908_/S vssd1 vssd1 vccd1 vccd1 _18259_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19097__A1 _21081_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21270_ _21444_/CLK _21270_/D repeater246/X vssd1 vssd1 vccd1 vccd1 _21270_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__14323__A1_N _20124_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20221_ _21484_/CLK _20221_/D repeater202/X vssd1 vssd1 vccd1 vccd1 _20221_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__19192__S1 _20122_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20152_ _21242_/CLK _20152_/D repeater189/X vssd1 vssd1 vccd1 vccd1 _20152_/Q sky130_fd_sc_hd__dfrtp_1
X_09963_ _20870_/Q vssd1 vssd1 vccd1 vccd1 _11199_/A sky130_fd_sc_hd__inv_2
XANTENNA__13669__B1 _13550_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__21296__RESET_B repeater208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20083_ _20590_/CLK _20083_/D repeater260/X vssd1 vssd1 vccd1 vccd1 _20083_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_112_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09894_ _20012_/Q _09887_/B _09893_/Y _20013_/Q _09887_/Y vssd1 vssd1 vccd1 vccd1
+ _20013_/D sky130_fd_sc_hd__a32o_1
XFILLER_85_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21225__RESET_B repeater249/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17804__C1 _17802_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18072__A2 _17205_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_82_HCLK_A clkbuf_4_13_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18956__S _18962_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20985_ _21141_/CLK _20985_/D repeater191/X vssd1 vssd1 vccd1 vccd1 _20985_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_3915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17161__A _21127_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18780__A0 _18848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20860__RESET_B repeater243/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_213_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18691__S _18898_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_241_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20178__RESET_B repeater200/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20107__RESET_B repeater259/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12270_ _20528_/Q vssd1 vssd1 vccd1 vccd1 _12270_/Y sky130_fd_sc_hd__inv_2
X_21468_ _21477_/CLK _21468_/D repeater204/X vssd1 vssd1 vccd1 vccd1 _21468_/Q sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_14_HCLK clkbuf_opt_2_HCLK/A vssd1 vssd1 vccd1 vccd1 _19765_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_209_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11221_ _21204_/Q _11219_/X _10884_/X _11220_/X vssd1 vssd1 vccd1 vccd1 _21204_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_135_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20419_ _20957_/CLK _20419_/D repeater187/X vssd1 vssd1 vccd1 vccd1 _20419_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__19183__S1 _20122_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21399_ _21405_/CLK _21399_/D repeater252/X vssd1 vssd1 vccd1 vccd1 _21399_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_134_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11152_ _19986_/Q vssd1 vssd1 vccd1 vccd1 _17169_/B sky130_fd_sc_hd__inv_2
XFILLER_96_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10103_ _20782_/Q vssd1 vssd1 vccd1 vccd1 _10103_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19027__S _19058_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15960_ _19554_/Q _15954_/X _15941_/X _15956_/X vssd1 vssd1 vccd1 vccd1 _19554_/D
+ sky130_fd_sc_hd__a22o_1
X_11083_ _11075_/B _11079_/X _11081_/Y _11082_/X _11060_/A vssd1 vssd1 vccd1 vccd1
+ _11084_/A sky130_fd_sc_hd__o32a_1
XFILLER_68_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input31_A HADDR[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_156_HCLK clkbuf_opt_1_HCLK/A vssd1 vssd1 vccd1 vccd1 _21452_/CLK sky130_fd_sc_hd__clkbuf_16
X_14911_ _20586_/Q vssd1 vssd1 vccd1 vccd1 _14911_/Y sky130_fd_sc_hd__inv_2
X_10034_ _10034_/A _10034_/B vssd1 vssd1 vccd1 vccd1 _10163_/A sky130_fd_sc_hd__or2_1
XFILLER_237_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15891_ _16235_/A vssd1 vssd1 vccd1 vccd1 _15891_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__18866__S _18926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17630_ _20175_/Q _17446_/X _17628_/X _17629_/X _17529_/Y vssd1 vssd1 vccd1 vccd1
+ _17630_/Y sky130_fd_sc_hd__o221ai_4
X_14842_ _20092_/Q vssd1 vssd1 vccd1 vccd1 _14961_/D sky130_fd_sc_hd__inv_2
XFILLER_84_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17561_ _21140_/Q vssd1 vssd1 vccd1 vccd1 _17561_/Y sky130_fd_sc_hd__inv_2
X_14773_ _14775_/A _14318_/X _15919_/A vssd1 vssd1 vccd1 vccd1 _14773_/X sky130_fd_sc_hd__o21a_1
XFILLER_90_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11985_ _15397_/A _11984_/X _15397_/A _11984_/X vssd1 vssd1 vccd1 vccd1 _11985_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_205_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19300_ _19828_/CLK _19300_/D vssd1 vssd1 vccd1 vccd1 _19300_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_244_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17071__A _19889_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16512_ _21093_/Q vssd1 vssd1 vccd1 vccd1 _16512_/Y sky130_fd_sc_hd__inv_2
XFILLER_205_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10936_ _21035_/Q vssd1 vssd1 vccd1 vccd1 _11812_/A sky130_fd_sc_hd__inv_2
X_13724_ _20328_/Q vssd1 vssd1 vccd1 vccd1 _15766_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_32_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17492_ _19522_/Q vssd1 vssd1 vccd1 vccd1 _17492_/Y sky130_fd_sc_hd__inv_2
XFILLER_189_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18771__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19231_ _19227_/X _19228_/X _19229_/X _19230_/X _20132_/Q _20133_/Q vssd1 vssd1 vccd1
+ vccd1 _19231_/X sky130_fd_sc_hd__mux4_2
XFILLER_16_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16443_ _19312_/Q _16441_/X _16335_/X _16442_/X vssd1 vssd1 vccd1 vccd1 _19312_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_231_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_repeater170_A _18897_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10867_ _21267_/Q _10864_/X _09670_/X _10866_/X vssd1 vssd1 vccd1 vccd1 _21267_/D
+ sky130_fd_sc_hd__a22o_1
X_13655_ _20365_/Q _13651_/X _13452_/X _13652_/X vssd1 vssd1 vccd1 vccd1 _20365_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_20_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19162_ _19702_/Q _19566_/Q _19558_/Q _19550_/Q _19280_/S0 _20122_/Q vssd1 vssd1
+ vccd1 vccd1 _19162_/X sky130_fd_sc_hd__mux4_2
X_12606_ _12606_/A vssd1 vssd1 vccd1 vccd1 _17060_/B sky130_fd_sc_hd__clkbuf_2
X_16374_ _19350_/Q _16370_/X _16212_/X _16371_/X vssd1 vssd1 vccd1 vccd1 _19350_/D
+ sky130_fd_sc_hd__a22o_1
X_13586_ input68/X vssd1 vssd1 vccd1 vccd1 _13586_/X sky130_fd_sc_hd__clkbuf_4
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10798_ _10812_/A vssd1 vssd1 vccd1 vccd1 _10798_/X sky130_fd_sc_hd__clkbuf_2
XPHY_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18113_ _21268_/Q _21240_/Q vssd1 vssd1 vccd1 vccd1 _18113_/X sky130_fd_sc_hd__and2_4
X_12537_ _11290_/A _12524_/X _11301_/A _12528_/X vssd1 vssd1 vccd1 vccd1 _20905_/D
+ sky130_fd_sc_hd__o22ai_1
X_15325_ _20031_/Q _15323_/X _13543_/X _15324_/X vssd1 vssd1 vccd1 vccd1 _20031_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_219_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19093_ _16677_/X _21085_/Q _19870_/D vssd1 vssd1 vccd1 vccd1 _19093_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12943__A _12961_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18044_ _20422_/Q vssd1 vssd1 vccd1 vccd1 _18044_/Y sky130_fd_sc_hd__inv_2
X_15256_ _20488_/Q _20067_/Q _15255_/Y _15081_/A vssd1 vssd1 vccd1 vccd1 _15259_/C
+ sky130_fd_sc_hd__o22a_1
X_12468_ _12468_/A vssd1 vssd1 vccd1 vccd1 _12490_/A sky130_fd_sc_hd__buf_1
XFILLER_126_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11419_ _11783_/B _11418_/X _11364_/X _11403_/A vssd1 vssd1 vccd1 vccd1 _21180_/D
+ sky130_fd_sc_hd__o22ai_1
XANTENNA__19174__S1 _20122_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11559__A _16332_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14207_ _14207_/A vssd1 vssd1 vccd1 vccd1 _14207_/X sky130_fd_sc_hd__buf_2
X_15187_ _15076_/A _15076_/B _15184_/Y _15179_/X vssd1 vssd1 vccd1 vccd1 _20062_/D
+ sky130_fd_sc_hd__a211oi_2
X_12399_ _12470_/A _12469_/C _12399_/C _12399_/D vssd1 vssd1 vccd1 vccd1 _12418_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_235_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14138_ _14124_/X _14138_/B _14138_/C _14138_/D vssd1 vssd1 vccd1 vccd1 _14171_/B
+ sky130_fd_sc_hd__and4b_1
X_19995_ _21196_/CLK _19995_/D repeater218/X vssd1 vssd1 vccd1 vccd1 _19995_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_180_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18946_ _19890_/Q _16690_/Y _18946_/S vssd1 vssd1 vccd1 vccd1 _18946_/X sky130_fd_sc_hd__mux2_1
X_14069_ _20259_/Q vssd1 vssd1 vccd1 vccd1 _14070_/A sky130_fd_sc_hd__inv_2
XFILLER_239_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18877_ _18876_/X _10731_/Y _18910_/S vssd1 vssd1 vccd1 vccd1 _18877_/X sky130_fd_sc_hd__mux2_1
XANTENNA__18776__S _18880_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17828_ _14702_/A _17818_/X _17838_/A _17819_/X _17827_/X vssd1 vssd1 vccd1 vccd1
+ _17828_/Y sky130_fd_sc_hd__o221ai_4
XANTENNA__10885__B1 _10884_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17759_ _19324_/Q vssd1 vssd1 vccd1 vccd1 _17759_/Y sky130_fd_sc_hd__inv_2
X_20770_ _21406_/CLK _20770_/D repeater213/X vssd1 vssd1 vccd1 vccd1 _20770_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_63_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_223_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19429_ _20331_/CLK _19429_/D vssd1 vssd1 vccd1 vccd1 _19429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_195_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20271__RESET_B repeater263/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_37_HCLK _20004_/CLK vssd1 vssd1 vccd1 vccd1 _20042_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__15328__B1 _13550_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12853__A _12853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21322_ _21341_/CLK _21322_/D repeater222/X vssd1 vssd1 vccd1 vccd1 _21322_/Q sky130_fd_sc_hd__dfrtp_1
Xclkbuf_2_0_0_HCLK clkbuf_2_1_0_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_1_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_135_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19165__S1 _20122_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21253_ _21255_/CLK _21253_/D repeater240/X vssd1 vssd1 vccd1 vccd1 _21253_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_209_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20204_ _20623_/CLK _20204_/D repeater194/X vssd1 vssd1 vccd1 vccd1 _20204_/Q sky130_fd_sc_hd__dfrtp_1
X_21184_ _21184_/CLK _21184_/D repeater220/X vssd1 vssd1 vccd1 vccd1 _21184_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_78_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20135_ _20136_/CLK _20135_/D repeater248/X vssd1 vssd1 vccd1 vccd1 _20135_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_89_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09946_ _20870_/Q vssd1 vssd1 vccd1 vccd1 _17060_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_225_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11668__A2 _11657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20066_ _20066_/CLK _20066_/D hold8/X vssd1 vssd1 vccd1 vccd1 _20066_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_219_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18686__S _18896_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09877_ _09846_/C _09876_/X _09873_/X vssd1 vssd1 vccd1 vccd1 _21441_/D sky130_fd_sc_hd__a21oi_1
XFILLER_58_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10876__B1 _09702_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_3_4_0_HCLK_A clkbuf_3_5_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater270 repeater272/X vssd1 vssd1 vccd1 vccd1 repeater270/X sky130_fd_sc_hd__buf_8
XPHY_4402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater281 hold8/X vssd1 vssd1 vccd1 vccd1 repeater281/X sky130_fd_sc_hd__buf_8
XFILLER_245_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11770_ _11770_/A vssd1 vssd1 vccd1 vccd1 _11770_/X sky130_fd_sc_hd__buf_1
XPHY_4468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20968_ _20971_/CLK _20968_/D repeater186/X vssd1 vssd1 vccd1 vccd1 _20968_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__13290__A1 _20552_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10721_ _21314_/Q _10725_/A _10718_/A _10712_/X vssd1 vssd1 vccd1 vccd1 _21314_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_3767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20899_ _21141_/CLK _20899_/D repeater212/X vssd1 vssd1 vccd1 vccd1 _20899_/Q sky130_fd_sc_hd__dfstp_1
XPHY_3789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13440_ _20470_/Q _13436_/X _13245_/X _13437_/X vssd1 vssd1 vccd1 vccd1 _20470_/D
+ sky130_fd_sc_hd__a22o_1
X_10652_ _10652_/A _10697_/A vssd1 vssd1 vccd1 vccd1 _10653_/B sky130_fd_sc_hd__or2_1
XANTENNA__18505__A0 _18848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13371_ _13377_/A vssd1 vssd1 vccd1 vccd1 _13371_/X sky130_fd_sc_hd__buf_1
X_10583_ _20745_/Q vssd1 vssd1 vccd1 vccd1 _10583_/Y sky130_fd_sc_hd__inv_2
XFILLER_166_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16235__A _16235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15110_ _15110_/A _15110_/B _15106_/X _15109_/X vssd1 vssd1 vccd1 vccd1 _15158_/A
+ sky130_fd_sc_hd__or4bb_4
X_12322_ _12322_/A _12358_/A vssd1 vssd1 vccd1 vccd1 _12323_/B sky130_fd_sc_hd__or2_2
XFILLER_154_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16090_ _19488_/Q _16087_/X _15879_/X _16088_/X vssd1 vssd1 vccd1 vccd1 _19488_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_182_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15041_ _20061_/Q vssd1 vssd1 vccd1 vccd1 _15075_/A sky130_fd_sc_hd__inv_2
X_12253_ _20949_/Q _12251_/Y _20941_/Q _12252_/Y vssd1 vssd1 vccd1 vccd1 _12253_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_181_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21147__RESET_B repeater212/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11204_ _15885_/A _14702_/A vssd1 vssd1 vccd1 vccd1 _11207_/A sky130_fd_sc_hd__or2_1
X_12184_ _12311_/A _20339_/Q _20957_/Q _12183_/Y vssd1 vssd1 vccd1 vccd1 _12184_/X
+ sky130_fd_sc_hd__o22a_1
X_18800_ _18799_/X _19246_/X _18930_/S vssd1 vssd1 vccd1 vccd1 _18800_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13594__A _13594_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11135_ _15466_/B vssd1 vssd1 vccd1 vccd1 _11176_/B sky130_fd_sc_hd__buf_1
X_19780_ _20432_/CLK _19780_/D vssd1 vssd1 vccd1 vccd1 _19780_/Q sky130_fd_sc_hd__dfxtp_1
X_16992_ _19975_/Q _16992_/B vssd1 vssd1 vccd1 vccd1 _16997_/B sky130_fd_sc_hd__or2_1
XFILLER_150_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18731_ _17634_/Y _10008_/Y _20870_/Q vssd1 vssd1 vccd1 vccd1 _18731_/X sky130_fd_sc_hd__mux2_1
X_15943_ _15943_/A vssd1 vssd1 vccd1 vccd1 _15943_/X sky130_fd_sc_hd__buf_1
X_11066_ _11066_/A _11066_/B vssd1 vssd1 vccd1 vccd1 _11067_/B sky130_fd_sc_hd__nand2_1
XANTENNA__18596__S _18910_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10017_ _10017_/A _10017_/B _20023_/D _10016_/X vssd1 vssd1 vccd1 vccd1 _11621_/B
+ sky130_fd_sc_hd__or4b_4
XANTENNA__10867__B1 _09670_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18662_ _18661_/X _20527_/Q _18910_/S vssd1 vssd1 vccd1 vccd1 _18662_/X sky130_fd_sc_hd__mux2_1
X_15874_ _19594_/Q _15864_/X _15873_/X _15867_/X vssd1 vssd1 vccd1 vccd1 _19594_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_36_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17613_ _19322_/Q vssd1 vssd1 vccd1 vccd1 _17613_/Y sky130_fd_sc_hd__inv_2
XFILLER_91_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14825_ _20108_/Q _14185_/X _14824_/Y vssd1 vssd1 vccd1 vccd1 _20108_/D sky130_fd_sc_hd__o21a_1
X_18593_ _18592_/X _10505_/X _18880_/S vssd1 vssd1 vccd1 vccd1 _18593_/X sky130_fd_sc_hd__mux2_2
XFILLER_221_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17544_ _17544_/A _17807_/B vssd1 vssd1 vccd1 vccd1 _17544_/Y sky130_fd_sc_hd__nor2_1
XFILLER_63_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20711__RESET_B repeater254/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14756_ _20133_/Q _14754_/Y _14755_/Y _14754_/A vssd1 vssd1 vccd1 vccd1 _20133_/D
+ sky130_fd_sc_hd__o22a_1
X_11968_ _13182_/B vssd1 vssd1 vccd1 vccd1 _13179_/B sky130_fd_sc_hd__inv_2
XFILLER_205_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13707_ _15424_/A vssd1 vssd1 vccd1 vccd1 _13707_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_220_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10919_ _21033_/Q vssd1 vssd1 vccd1 vccd1 _11810_/A sky130_fd_sc_hd__inv_2
X_17475_ _17471_/Y _17472_/X _17473_/Y _17474_/X vssd1 vssd1 vccd1 vccd1 _17475_/X
+ sky130_fd_sc_hd__o22a_1
X_11899_ _19114_/X _10992_/X _10988_/X vssd1 vssd1 vccd1 vccd1 _11900_/B sky130_fd_sc_hd__a21oi_1
X_14687_ _10985_/Y _14674_/X _18975_/X _12742_/A _16526_/B vssd1 vssd1 vccd1 vccd1
+ _14692_/A sky130_fd_sc_hd__o2111a_1
XFILLER_177_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19214_ _17674_/Y _17675_/Y _17676_/Y _17677_/Y _19275_/S0 _21004_/Q vssd1 vssd1
+ vccd1 vccd1 _19214_/X sky130_fd_sc_hd__mux4_2
X_16426_ _19321_/Q _16420_/X _15873_/A _16422_/X vssd1 vssd1 vccd1 vccd1 _19321_/D
+ sky130_fd_sc_hd__a22o_1
X_13638_ _20376_/Q _13632_/X _13426_/X _13634_/X vssd1 vssd1 vccd1 vccd1 _20376_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_60_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19145_ _19657_/Q _19649_/Q _19633_/Q _19817_/Q _19285_/S0 _21017_/Q vssd1 vssd1
+ vccd1 vccd1 _19145_/X sky130_fd_sc_hd__mux4_2
X_16357_ _19358_/Q _16352_/X _16295_/X _16353_/X vssd1 vssd1 vccd1 vccd1 _19358_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_201_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13569_ _20415_/Q _13566_/X _13485_/X _13567_/X vssd1 vssd1 vccd1 vccd1 _20415_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12673__A input53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15308_ _20038_/Q _15302_/A _20037_/Q _15305_/X vssd1 vssd1 vccd1 vccd1 _20038_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_200_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19076_ _16727_/X _20899_/Q _19908_/D vssd1 vssd1 vccd1 vccd1 _19076_/X sky130_fd_sc_hd__mux2_1
X_16288_ _20327_/Q vssd1 vssd1 vccd1 vccd1 _16288_/X sky130_fd_sc_hd__clkbuf_2
X_18027_ _18018_/X _18027_/B _18027_/C vssd1 vssd1 vccd1 vccd1 _18027_/Y sky130_fd_sc_hd__nand3b_4
XANTENNA__19147__S1 _21017_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15239_ _20483_/Q vssd1 vssd1 vccd1 vccd1 _15239_/Y sky130_fd_sc_hd__inv_2
XFILLER_173_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19965__RESET_B repeater184/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09800_ _09804_/C _09800_/B vssd1 vssd1 vccd1 vccd1 _09800_/Y sky130_fd_sc_hd__nor2_1
XFILLER_99_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19978_ _20809_/CLK _19978_/D repeater270/X vssd1 vssd1 vccd1 vccd1 _19978_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_113_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09731_ _20154_/Q vssd1 vssd1 vccd1 vccd1 _09731_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18929_ _18928_/X _11986_/Y _18929_/S vssd1 vssd1 vccd1 vccd1 _18929_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_0_HCLK HCLK vssd1 vssd1 vccd1 vccd1 clkbuf_0_HCLK/X sky130_fd_sc_hd__clkbuf_16
X_09662_ input69/X vssd1 vssd1 vccd1 vccd1 _13311_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_28_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_242_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20822_ _21374_/CLK _20822_/D repeater256/X vssd1 vssd1 vccd1 vccd1 _20822_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20753_ _21342_/CLK _20753_/D repeater210/X vssd1 vssd1 vccd1 vccd1 _20753_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__15549__B1 _15548_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20684_ _21480_/CLK _20684_/D repeater208/X vssd1 vssd1 vccd1 vccd1 _20684_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_210_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13679__A _13679_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21305_ _21480_/CLK _21305_/D repeater206/X vssd1 vssd1 vccd1 vccd1 _21305_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__19138__S1 _21017_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21236_ _21239_/CLK _21236_/D repeater189/X vssd1 vssd1 vccd1 vccd1 _21236_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_104_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21167_ _21167_/CLK _21167_/D repeater225/X vssd1 vssd1 vccd1 vccd1 _21167_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_131_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14303__A _20890_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20118_ _21452_/CLK _20118_/D repeater247/X vssd1 vssd1 vccd1 vccd1 _20118_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_131_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12838__A1 _20760_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09929_ _20014_/Q _21431_/Q _09929_/S vssd1 vssd1 vccd1 vccd1 _21431_/D sky130_fd_sc_hd__mux2_1
X_21098_ _21429_/CLK _21098_/D repeater231/X vssd1 vssd1 vccd1 vccd1 _21098_/Q sky130_fd_sc_hd__dfrtp_1
X_20049_ _20480_/CLK _20049_/D repeater281/X vssd1 vssd1 vccd1 vccd1 _20049_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_92_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12940_ _20716_/Q _12935_/X _12855_/X _12937_/X vssd1 vssd1 vccd1 vccd1 _20716_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_219_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12871_ _20743_/Q _12867_/X _12550_/X _12868_/X vssd1 vssd1 vccd1 vccd1 _20743_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16985__C1 _16984_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20193__RESET_B repeater200/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14610_ _14624_/A vssd1 vssd1 vccd1 vccd1 _14610_/X sky130_fd_sc_hd__buf_1
XPHY_4243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11822_ _11822_/A _11822_/B vssd1 vssd1 vccd1 vccd1 _11822_/Y sky130_fd_sc_hd__nor2_1
XPHY_4254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15590_ _15793_/A vssd1 vssd1 vccd1 vccd1 _15590_/X sky130_fd_sc_hd__clkbuf_2
XPHY_4265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20122__RESET_B repeater247/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_230_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11753_ _21053_/Q _11761_/A _11753_/C vssd1 vssd1 vccd1 vccd1 _11755_/A sky130_fd_sc_hd__or3_1
XFILLER_26_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14541_ _14541_/A vssd1 vssd1 vccd1 vccd1 _14541_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10704_ _10704_/A _10704_/B vssd1 vssd1 vccd1 vccd1 _10715_/A sky130_fd_sc_hd__or2_1
XPHY_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19040__S _19046_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17260_ _19342_/Q vssd1 vssd1 vccd1 vccd1 _17260_/Y sky130_fd_sc_hd__inv_2
X_14472_ _14566_/B vssd1 vssd1 vccd1 vccd1 _14472_/X sky130_fd_sc_hd__buf_1
X_11684_ _12548_/A vssd1 vssd1 vccd1 vccd1 _11684_/X sky130_fd_sc_hd__clkbuf_2
XPHY_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16211_ _19432_/Q _16206_/X _16210_/X _16208_/X vssd1 vssd1 vccd1 vccd1 _19432_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__21399__RESET_B repeater252/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10635_ _20753_/Q vssd1 vssd1 vccd1 vccd1 _10635_/Y sky130_fd_sc_hd__inv_2
XPHY_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13589__A _13595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13423_ _20479_/Q _13417_/X _13422_/X _13420_/X vssd1 vssd1 vccd1 vccd1 _20479_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_174_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17191_ _20397_/Q vssd1 vssd1 vccd1 vccd1 _17191_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12774__B1 _09621_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16142_ _21449_/Q vssd1 vssd1 vccd1 vccd1 _16142_/X sky130_fd_sc_hd__buf_1
X_13354_ _20516_/Q _13351_/X _13219_/X _13352_/X vssd1 vssd1 vccd1 vccd1 _20516_/D
+ sky130_fd_sc_hd__a22o_1
X_10566_ _10654_/A _10653_/A _10566_/C _10566_/D vssd1 vssd1 vccd1 vccd1 _10573_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_155_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12305_ _12305_/A _12389_/A vssd1 vssd1 vccd1 vccd1 _12306_/B sky130_fd_sc_hd__or2_2
XFILLER_154_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19129__S1 _21017_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16073_ _19497_/Q _16071_/X _15769_/X _16072_/X vssd1 vssd1 vccd1 vccd1 _19497_/D
+ sky130_fd_sc_hd__a22o_1
X_13285_ _20554_/Q _13276_/X _13284_/X _13278_/X vssd1 vssd1 vccd1 vccd1 _20554_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_115_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10497_ _20670_/Q vssd1 vssd1 vccd1 vccd1 _17544_/A sky130_fd_sc_hd__inv_2
XFILLER_182_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19901_ _21185_/CLK _19901_/D repeater224/X vssd1 vssd1 vccd1 vccd1 _19901_/Q sky130_fd_sc_hd__dfrtp_1
Xclkbuf_4_9_0_HCLK clkbuf_4_9_0_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_9_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_5_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12236_ _20507_/Q vssd1 vssd1 vccd1 vccd1 _12236_/Y sky130_fd_sc_hd__inv_2
X_15024_ _15019_/A _15019_/B _15019_/C vssd1 vssd1 vccd1 vccd1 _15025_/B sky130_fd_sc_hd__o21a_1
X_19832_ _19834_/CLK _19832_/D vssd1 vssd1 vccd1 vccd1 _19832_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12167_ _20965_/Q _12164_/Y _12318_/A _20347_/Q _12166_/X vssd1 vssd1 vccd1 vccd1
+ _12175_/B sky130_fd_sc_hd__a221o_1
XFILLER_123_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11118_ _21225_/Q _09744_/X _21226_/Q _11117_/X vssd1 vssd1 vccd1 vccd1 _11118_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__20963__RESET_B repeater185/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19763_ _19765_/CLK _19763_/D vssd1 vssd1 vccd1 vccd1 _19763_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16975_ _19971_/Q vssd1 vssd1 vccd1 vccd1 _16975_/Y sky130_fd_sc_hd__inv_2
X_12098_ _20372_/Q vssd1 vssd1 vccd1 vccd1 _17806_/A sky130_fd_sc_hd__inv_2
XFILLER_96_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18714_ _18713_/X _10123_/Y _18879_/S vssd1 vssd1 vccd1 vccd1 _18714_/X sky130_fd_sc_hd__mux2_1
XFILLER_232_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11049_ _20138_/Q vssd1 vssd1 vccd1 vccd1 _11050_/A sky130_fd_sc_hd__inv_2
X_15926_ _19570_/Q _15920_/X _15785_/X _15922_/X vssd1 vssd1 vccd1 vccd1 _19570_/D
+ sky130_fd_sc_hd__a22o_1
X_19694_ _19776_/CLK _19694_/D vssd1 vssd1 vccd1 vccd1 _19694_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11501__A1 _11486_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput7 HADDR[15] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_1
XFILLER_209_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18645_ _18644_/X _10289_/A _18886_/S vssd1 vssd1 vccd1 vccd1 _18645_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15857_ _15857_/A vssd1 vssd1 vccd1 vccd1 _15857_/X sky130_fd_sc_hd__buf_1
XANTENNA__12668__A input55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_224_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14808_ _14803_/A _14803_/B _14804_/A _14807_/X vssd1 vssd1 vccd1 vccd1 _14808_/X
+ sky130_fd_sc_hd__o211a_1
X_18576_ _18575_/X _14079_/A _18904_/S vssd1 vssd1 vccd1 vccd1 _18576_/X sky130_fd_sc_hd__mux2_1
XFILLER_224_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15788_ _15788_/A vssd1 vssd1 vccd1 vccd1 _15788_/X sky130_fd_sc_hd__buf_2
X_17527_ _17368_/X _17526_/Y _20119_/Q vssd1 vssd1 vccd1 vccd1 _17527_/X sky130_fd_sc_hd__o21a_1
X_14739_ _17684_/A _16433_/A vssd1 vssd1 vccd1 vccd1 _14740_/S sky130_fd_sc_hd__or2_1
XFILLER_189_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17458_ _21047_/Q vssd1 vssd1 vccd1 vccd1 _17458_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16409_ _19332_/Q _16406_/X _16196_/X _16408_/X vssd1 vssd1 vccd1 vccd1 _19332_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_192_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17389_ _21188_/Q vssd1 vssd1 vccd1 vccd1 _17389_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19128_ _19758_/Q _19750_/Q _19742_/Q _19734_/Q _19285_/S0 _21017_/Q vssd1 vssd1
+ vccd1 vccd1 _19128_/X sky130_fd_sc_hd__mux4_2
XFILLER_173_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19059_ _21192_/Q _21134_/Q _19910_/Q vssd1 vssd1 vccd1 vccd1 _19059_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21021_ _21021_/CLK _21021_/D repeater238/X vssd1 vssd1 vccd1 vccd1 _21021_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_99_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09714_ _21456_/Q vssd1 vssd1 vccd1 vccd1 _09793_/C sky130_fd_sc_hd__inv_2
XFILLER_56_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09645_ _12853_/A vssd1 vssd1 vccd1 vccd1 _09645_/X sky130_fd_sc_hd__buf_4
XFILLER_82_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_137_HCLK_A clkbuf_4_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20805_ _21011_/CLK _20805_/D repeater235/X vssd1 vssd1 vccd1 vccd1 _20805_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_212_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20736_ _21349_/CLK _20736_/D repeater210/X vssd1 vssd1 vccd1 vccd1 _20736_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_196_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20667_ _21306_/CLK _20667_/D repeater207/X vssd1 vssd1 vccd1 vccd1 _20667_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_177_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10420_ _21344_/Q _10177_/A _10418_/A _10364_/X vssd1 vssd1 vccd1 vccd1 _21344_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_164_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20598_ _21011_/CLK _20598_/D repeater235/X vssd1 vssd1 vccd1 vccd1 _20598_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_164_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10351_ _20711_/Q vssd1 vssd1 vccd1 vccd1 _17812_/A sky130_fd_sc_hd__inv_2
XFILLER_136_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18204__S _18886_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13070_ _20655_/Q _13066_/X _12920_/X _13067_/X vssd1 vssd1 vccd1 vccd1 _20655_/D
+ sky130_fd_sc_hd__a22o_1
X_10282_ _10282_/A _10380_/A vssd1 vssd1 vccd1 vccd1 _10283_/B sky130_fd_sc_hd__or2_2
XFILLER_140_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12021_ _19073_/X _12017_/X _20992_/Q _12018_/X vssd1 vssd1 vccd1 vccd1 _20992_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11657__A _11657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21219_ _21222_/CLK _21219_/D repeater235/X vssd1 vssd1 vccd1 vccd1 _21219_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_104_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11166__A1_N _11123_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20374__RESET_B repeater186/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19035__S _19046_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16760_ _16760_/A vssd1 vssd1 vccd1 vccd1 _16766_/B sky130_fd_sc_hd__inv_2
XANTENNA__12287__A2 _20501_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13972_ _13972_/A _13972_/B _13972_/C _13972_/D vssd1 vssd1 vccd1 vccd1 _13972_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_86_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15711_ _15717_/A vssd1 vssd1 vccd1 vccd1 _15711_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_246_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12923_ _20723_/Q _12915_/X _12922_/X _12916_/X vssd1 vssd1 vccd1 vccd1 _20723_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_207_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16691_ _16691_/A _18946_/X vssd1 vssd1 vccd1 vccd1 _19890_/D sky130_fd_sc_hd__nor2_1
XANTENNA__18874__S _18874_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18430_ _18429_/X _10129_/Y _18885_/S vssd1 vssd1 vccd1 vccd1 _18430_/X sky130_fd_sc_hd__mux2_1
X_15642_ _15648_/A vssd1 vssd1 vccd1 vccd1 _15642_/X sky130_fd_sc_hd__buf_1
XFILLER_234_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12854_ _20752_/Q _12848_/X _12853_/X _12851_/X vssd1 vssd1 vccd1 vccd1 _20752_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18361_ _18360_/X _16863_/A _18667_/S vssd1 vssd1 vccd1 vccd1 _18361_/X sky130_fd_sc_hd__mux2_1
X_11805_ _11805_/A _11859_/A vssd1 vssd1 vccd1 vccd1 _11855_/A sky130_fd_sc_hd__or2_1
XPHY_4084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output100_A _18090_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15573_ _19734_/Q _15568_/X _15526_/X _15569_/X vssd1 vssd1 vccd1 vccd1 _19734_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12785_ _12785_/A vssd1 vssd1 vccd1 vccd1 _12804_/A sky130_fd_sc_hd__clkbuf_2
XPHY_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11798__A1 input70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17312_ _17310_/Y _17196_/X _17311_/Y _17232_/X vssd1 vssd1 vccd1 vccd1 _17312_/X
+ sky130_fd_sc_hd__o22a_1
X_14524_ _14524_/A _14524_/B _14524_/C vssd1 vssd1 vccd1 vccd1 _20210_/D sky130_fd_sc_hd__nor3_1
XPHY_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11736_ _13166_/A vssd1 vssd1 vccd1 vccd1 _11736_/X sky130_fd_sc_hd__clkbuf_2
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18292_ _18291_/X _20518_/Q _18910_/S vssd1 vssd1 vccd1 vccd1 _18292_/X sky130_fd_sc_hd__mux2_1
XFILLER_230_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_59_HCLK_A clkbuf_4_14_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17243_ _19407_/Q vssd1 vssd1 vccd1 vccd1 _17243_/Y sky130_fd_sc_hd__inv_2
XPHY_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14455_ _14464_/B vssd1 vssd1 vccd1 vccd1 _14488_/A sky130_fd_sc_hd__buf_1
XANTENNA_repeater250_A repeater251/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11667_ _16634_/A _11667_/B vssd1 vssd1 vccd1 vccd1 _11676_/S sky130_fd_sc_hd__or2_2
XFILLER_128_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21162__RESET_B repeater226/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13406_ _20488_/Q _13404_/X _13287_/X _13405_/X vssd1 vssd1 vccd1 vccd1 _20488_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10618_ _20763_/Q vssd1 vssd1 vccd1 vccd1 _10618_/Y sky130_fd_sc_hd__inv_2
X_17174_ _20497_/Q _17174_/B vssd1 vssd1 vccd1 vccd1 _17174_/Y sky130_fd_sc_hd__nor2_1
XPHY_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14386_ _21482_/Q _20228_/Q _14385_/Y _14461_/C vssd1 vssd1 vccd1 vccd1 _14401_/A
+ sky130_fd_sc_hd__o22a_1
X_11598_ _11598_/A vssd1 vssd1 vccd1 vccd1 _11598_/X sky130_fd_sc_hd__buf_1
XFILLER_6_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16125_ _20325_/Q vssd1 vssd1 vccd1 vccd1 _16125_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_227_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10549_ _21321_/Q vssd1 vssd1 vccd1 vccd1 _10551_/C sky130_fd_sc_hd__inv_2
X_13337_ _20527_/Q _13331_/X _13272_/X _13334_/X vssd1 vssd1 vccd1 vccd1 _20527_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_4_7_0_HCLK_A clkbuf_4_7_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12951__A _12961_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16056_ _16056_/A vssd1 vssd1 vccd1 vccd1 _16056_/X sky130_fd_sc_hd__buf_1
XFILLER_142_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13268_ _13294_/A vssd1 vssd1 vccd1 vccd1 _13268_/X sky130_fd_sc_hd__buf_1
XFILLER_131_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13172__B1 _13171_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15007_ _20087_/Q _15006_/Y _14978_/A _14866_/B vssd1 vssd1 vccd1 vccd1 _20087_/D
+ sky130_fd_sc_hd__o211a_1
X_12219_ _12432_/C _20524_/Q _12256_/A _20504_/Q _12218_/X vssd1 vssd1 vccd1 vccd1
+ _12232_/B sky130_fd_sc_hd__o221a_1
X_13199_ _20593_/Q _13192_/X _12993_/X _13195_/X vssd1 vssd1 vccd1 vccd1 _20593_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_243_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19815_ _20172_/CLK _19815_/D vssd1 vssd1 vccd1 vccd1 _19815_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13782__A _20609_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16958_ _16958_/A _19968_/Q _16958_/C vssd1 vssd1 vccd1 vccd1 _16963_/B sky130_fd_sc_hd__or3_1
X_19746_ _19765_/CLK _19746_/D vssd1 vssd1 vccd1 vccd1 _19746_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09679__B1 _09676_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20044__RESET_B repeater276/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15909_ _19579_/Q _15904_/X _15871_/X _15906_/X vssd1 vssd1 vccd1 vccd1 _19579_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_225_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19677_ _19813_/CLK _19677_/D vssd1 vssd1 vccd1 vccd1 _19677_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__18784__S _18784_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16889_ _16889_/A _16889_/B vssd1 vssd1 vccd1 vccd1 _16889_/X sky130_fd_sc_hd__or2_1
XANTENNA__15216__A2 _14970_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18628_ _17079_/Y _12042_/Y _18908_/S vssd1 vssd1 vccd1 vccd1 _18628_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18559_ _18558_/X _16931_/A _18680_/S vssd1 vssd1 vccd1 vccd1 _18559_/X sky130_fd_sc_hd__mux2_2
XFILLER_178_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20521_ _20943_/CLK _20521_/D repeater275/X vssd1 vssd1 vccd1 vccd1 _20521_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_166_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10646__A _20699_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15924__B1 _15891_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20452_ _20480_/CLK _20452_/D repeater183/X vssd1 vssd1 vccd1 vccd1 _20452_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_21_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19210__S0 _20130_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19980__RESET_B repeater270/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20383_ _20971_/CLK _20383_/D repeater183/X vssd1 vssd1 vccd1 vccd1 _20383_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_119_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15152__A1 _20441_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput130 _20003_/Q vssd1 vssd1 vccd1 vccd1 RsTx_S0 sky130_fd_sc_hd__clkbuf_2
Xoutput141 _21185_/Q vssd1 vssd1 vccd1 vccd1 scl_oen_o_S5 sky130_fd_sc_hd__clkbuf_2
XANTENNA__18959__S _18962_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20814__RESET_B repeater212/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_217_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21004_ _21009_/CLK _21004_/D repeater235/X vssd1 vssd1 vccd1 vccd1 _21004_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_130_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17164__A _21136_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19277__S0 _19280_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18694__S _18850_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09628_ input50/X vssd1 vssd1 vccd1 vccd1 _09628_/X sky130_fd_sc_hd__buf_4
XFILLER_244_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11229__B1 _10898_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_231_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18157__A1 _20760_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11940__A _11940_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12570_ _12575_/A vssd1 vssd1 vccd1 vccd1 _18242_/S sky130_fd_sc_hd__buf_6
XFILLER_212_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_239_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11521_ _16711_/A _11497_/A _17064_/A _11520_/Y _11523_/S vssd1 vssd1 vccd1 vccd1
+ _11522_/A sky130_fd_sc_hd__o32a_1
XFILLER_12_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20719_ _20724_/CLK _20719_/D repeater264/X vssd1 vssd1 vccd1 vccd1 _20719_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12729__A0 _11179_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14240_ _19900_/Q _14240_/B vssd1 vssd1 vccd1 vccd1 _14241_/B sky130_fd_sc_hd__or2_1
X_11452_ _21164_/Q _11452_/B vssd1 vssd1 vccd1 vccd1 _11453_/B sky130_fd_sc_hd__or2_1
XFILLER_149_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19201__S0 _20132_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10403_ _21355_/Q _10405_/A _10395_/X _10271_/B vssd1 vssd1 vccd1 vccd1 _21355_/D
+ sky130_fd_sc_hd__o211a_1
X_14171_ _14171_/A _14171_/B _14171_/C _14171_/D vssd1 vssd1 vccd1 vccd1 _14176_/A
+ sky130_fd_sc_hd__and4_1
X_11383_ _11384_/C _11384_/B _11385_/A vssd1 vssd1 vccd1 vccd1 _11410_/B sky130_fd_sc_hd__and3b_1
XFILLER_180_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13122_ _20626_/Q _13120_/X _12996_/X _13121_/X vssd1 vssd1 vccd1 vccd1 _20626_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_input61_A HWDATA[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10334_ _10284_/A _20728_/Q _10270_/A _20714_/Q vssd1 vssd1 vccd1 vccd1 _10334_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_180_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18869__S _18929_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17930_ _18425_/X _17926_/X _18413_/X _17927_/X _17929_/X vssd1 vssd1 vccd1 vccd1
+ _17936_/B sky130_fd_sc_hd__o221a_2
XFILLER_97_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13053_ _13078_/A vssd1 vssd1 vccd1 vccd1 _13080_/A sky130_fd_sc_hd__inv_2
XFILLER_180_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10265_ _10265_/A _10412_/A vssd1 vssd1 vccd1 vccd1 _10266_/B sky130_fd_sc_hd__or2_2
XFILLER_133_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12004_ _21185_/Q vssd1 vssd1 vccd1 vccd1 _12006_/A sky130_fd_sc_hd__inv_2
XFILLER_133_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17861_ _17861_/A vssd1 vssd1 vccd1 vccd1 _17861_/X sky130_fd_sc_hd__buf_1
X_10196_ _10196_/A vssd1 vssd1 vccd1 vccd1 _10196_/Y sky130_fd_sc_hd__inv_2
X_16812_ _19934_/Q vssd1 vssd1 vccd1 vccd1 _16815_/A sky130_fd_sc_hd__inv_2
X_19600_ _21021_/CLK _19600_/D vssd1 vssd1 vccd1 vccd1 _19600_/Q sky130_fd_sc_hd__dfxtp_1
X_17792_ _21143_/Q vssd1 vssd1 vccd1 vccd1 _17792_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19268__S0 _20130_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19531_ _21462_/CLK _19531_/D vssd1 vssd1 vccd1 vccd1 _19531_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_207_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16743_ _16556_/Y _16554_/Y _16585_/A vssd1 vssd1 vccd1 vccd1 _19910_/D sky130_fd_sc_hd__o21a_1
XFILLER_47_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13955_ _20655_/Q _13971_/A _20651_/Q _13884_/A vssd1 vssd1 vccd1 vccd1 _13955_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_246_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19462_ _21234_/CLK _19462_/D vssd1 vssd1 vccd1 vccd1 _19462_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12906_ _20733_/Q _12901_/X _12656_/X _12904_/X vssd1 vssd1 vccd1 vccd1 _20733_/D
+ sky130_fd_sc_hd__a22o_1
X_16674_ _21162_/Q _11450_/B _11451_/B vssd1 vssd1 vccd1 vccd1 _16674_/X sky130_fd_sc_hd__a21bo_1
XFILLER_47_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13886_ _13972_/A _13996_/A vssd1 vssd1 vccd1 vccd1 _13887_/B sky130_fd_sc_hd__or2_2
XFILLER_34_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18413_ _18412_/X _14085_/A _18850_/S vssd1 vssd1 vccd1 vccd1 _18413_/X sky130_fd_sc_hd__mux2_1
X_15625_ _15632_/A vssd1 vssd1 vccd1 vccd1 _15625_/X sky130_fd_sc_hd__buf_1
X_12837_ _20761_/Q _12835_/X _12673_/X _12836_/X vssd1 vssd1 vccd1 vccd1 _20761_/D
+ sky130_fd_sc_hd__a22o_1
X_19393_ _21222_/CLK _19393_/D vssd1 vssd1 vccd1 vccd1 _19393_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__21343__RESET_B repeater205/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10127__A2_N _20787_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_120_HCLK_A clkbuf_opt_3_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18344_ _18343_/X _14911_/Y _18907_/S vssd1 vssd1 vccd1 vccd1 _18344_/X sky130_fd_sc_hd__mux2_2
XFILLER_15_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15556_ _19744_/Q _15553_/X _15521_/X _15554_/X vssd1 vssd1 vccd1 vccd1 _19744_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12768_ _20799_/Q _12765_/X _12666_/X _12766_/X vssd1 vssd1 vccd1 vccd1 _20799_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14507_ _14507_/A vssd1 vssd1 vccd1 vccd1 _14507_/Y sky130_fd_sc_hd__inv_2
X_11719_ _21068_/Q _11713_/X _11560_/X _11715_/X vssd1 vssd1 vccd1 vccd1 _21068_/D
+ sky130_fd_sc_hd__a22o_1
X_18275_ _19166_/X _21270_/Q _18281_/S vssd1 vssd1 vccd1 vccd1 _18275_/X sky130_fd_sc_hd__mux2_1
X_15487_ _16127_/A vssd1 vssd1 vccd1 vccd1 _15487_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_202_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12699_ _13313_/A vssd1 vssd1 vccd1 vccd1 _12699_/X sky130_fd_sc_hd__clkbuf_4
XPHY_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17226_ _17226_/A vssd1 vssd1 vccd1 vccd1 _17853_/A sky130_fd_sc_hd__buf_1
X_14438_ _21466_/Q vssd1 vssd1 vccd1 vccd1 _14438_/Y sky130_fd_sc_hd__inv_2
XFILLER_174_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput10 HADDR[18] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__clkbuf_1
Xinput21 HADDR[28] vssd1 vssd1 vccd1 vccd1 input21/X sky130_fd_sc_hd__buf_1
Xclkbuf_leaf_70_HCLK clkbuf_opt_7_HCLK/A vssd1 vssd1 vccd1 vccd1 _21484_/CLK sky130_fd_sc_hd__clkbuf_16
Xinput32 HADDR[9] vssd1 vssd1 vccd1 vccd1 input32/X sky130_fd_sc_hd__clkbuf_1
Xinput43 HWDATA[14] vssd1 vssd1 vccd1 vccd1 input43/X sky130_fd_sc_hd__clkbuf_2
XFILLER_190_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput54 HWDATA[24] vssd1 vssd1 vccd1 vccd1 input54/X sky130_fd_sc_hd__clkbuf_4
XFILLER_156_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17157_ _17169_/A _17169_/B _17169_/C _17157_/D vssd1 vssd1 vccd1 vccd1 _17548_/A
+ sky130_fd_sc_hd__or4_4
X_14369_ _14461_/B _14486_/A vssd1 vssd1 vccd1 vccd1 _14370_/B sky130_fd_sc_hd__or2_2
Xinput65 HWDATA[5] vssd1 vssd1 vccd1 vccd1 input65/X sky130_fd_sc_hd__clkbuf_4
Xinput76 scl_i_S5 vssd1 vssd1 vccd1 vccd1 input76/X sky130_fd_sc_hd__clkbuf_1
XFILLER_171_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16108_ _16119_/A vssd1 vssd1 vccd1 vccd1 _16108_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__15134__A1 _20456_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17088_ _20633_/Q _20323_/Q vssd1 vssd1 vccd1 vccd1 _17088_/X sky130_fd_sc_hd__and2_2
XFILLER_143_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16331__B1 _16237_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18779__S _18898_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13145__B1 _13144_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16039_ _19516_/Q _16035_/X _15973_/X _16037_/X vssd1 vssd1 vccd1 vccd1 _19516_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__20296__RESET_B repeater262/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20225__RESET_B repeater202/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19259__S0 _20130_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19729_ _19784_/CLK _19729_/D vssd1 vssd1 vccd1 vccd1 _19729_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16398__B1 _16332_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_225_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12959__B1 _12872_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20900__SET_B repeater212/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21013__RESET_B repeater238/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_42_HCLK_A clkbuf_4_11_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20504_ _20930_/CLK _20504_/D repeater267/X vssd1 vssd1 vccd1 vccd1 _20504_/Q sky130_fd_sc_hd__dfrtp_2
X_21484_ _21484_/CLK _21484_/D repeater200/X vssd1 vssd1 vccd1 vccd1 _21484_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_166_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20435_ _20937_/CLK _20435_/D repeater278/X vssd1 vssd1 vccd1 vccd1 _20435_/Q sky130_fd_sc_hd__dfrtp_1
X_20366_ _20951_/CLK _20366_/D repeater271/X vssd1 vssd1 vccd1 vccd1 _20366_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__16322__B1 _16012_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18689__S _18896_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13136__B1 _12930_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20297_ _20661_/CLK _20297_/D repeater262/X vssd1 vssd1 vccd1 vccd1 _20297_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_88_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10050_ _21387_/Q vssd1 vssd1 vccd1 vccd1 _10052_/C sky130_fd_sc_hd__inv_2
XFILLER_248_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11654__B _17157_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13740_ _20616_/Q vssd1 vssd1 vccd1 vccd1 _17941_/A sky130_fd_sc_hd__inv_2
XFILLER_17_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10952_ _21030_/Q vssd1 vssd1 vccd1 vccd1 _11807_/A sky130_fd_sc_hd__inv_2
XFILLER_244_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13671_ _20357_/Q _13667_/X _13555_/X _13668_/X vssd1 vssd1 vccd1 vccd1 _20357_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_73_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10883_ _21258_/Q _10879_/X _09666_/X _10881_/X vssd1 vssd1 vccd1 vccd1 _21258_/D
+ sky130_fd_sc_hd__a22o_1
X_15410_ _19806_/Q _15405_/X _15355_/X _15406_/X vssd1 vssd1 vccd1 vccd1 _19806_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12622_ input7/X _12619_/X _20858_/Q _12620_/X vssd1 vssd1 vccd1 vccd1 _20858_/D
+ sky130_fd_sc_hd__o22a_1
XPHY_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16390_ _19341_/Q _16385_/X _16375_/X _16386_/X vssd1 vssd1 vccd1 vccd1 _19341_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13611__A1 _20393_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_93_HCLK clkbuf_4_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20929_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15341_ _19836_/Q _15337_/X _14262_/X _15339_/X vssd1 vssd1 vccd1 vccd1 _19836_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12553_ _12553_/A vssd1 vssd1 vccd1 vccd1 _12553_/X sky130_fd_sc_hd__buf_1
XPHY_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20505__CLK _20930_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11504_ _15385_/A vssd1 vssd1 vccd1 vccd1 _11504_/X sky130_fd_sc_hd__buf_4
X_18060_ _20838_/Q vssd1 vssd1 vccd1 vccd1 _18060_/Y sky130_fd_sc_hd__inv_2
XFILLER_156_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15272_ _20480_/Q _15073_/A _17938_/A _20061_/Q vssd1 vssd1 vccd1 vccd1 _15272_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12484_ _20925_/Q _12483_/Y _12474_/B _12480_/X vssd1 vssd1 vccd1 vccd1 _20925_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12178__B2 _20341_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17011_ _19980_/Q vssd1 vssd1 vccd1 vccd1 _17011_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13375__B1 _13245_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14223_ _20264_/Q _14222_/Y _14076_/B _14191_/X vssd1 vssd1 vccd1 vccd1 _20264_/D
+ sky130_fd_sc_hd__o211a_1
X_11435_ _11386_/B _11421_/A _11410_/B _11420_/X vssd1 vssd1 vccd1 vccd1 _21170_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__20736__RESET_B repeater210/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11366_ _21173_/Q _11390_/C _11366_/C vssd1 vssd1 vccd1 vccd1 _11379_/C sky130_fd_sc_hd__or3_1
X_14154_ _20540_/Q _14079_/A _17541_/A _20263_/Q _14153_/X vssd1 vssd1 vccd1 vccd1
+ _14155_/D sky130_fd_sc_hd__o221a_1
XFILLER_152_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18599__S _18886_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13105_ _12978_/X _20633_/Q _13105_/S vssd1 vssd1 vccd1 vccd1 _20633_/D sky130_fd_sc_hd__mux2_1
X_10317_ _20731_/Q vssd1 vssd1 vccd1 vccd1 _10317_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11297_ _20904_/Q vssd1 vssd1 vccd1 vccd1 _11311_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_18962_ _19852_/Q _16633_/Y _18962_/S vssd1 vssd1 vccd1 vccd1 _18962_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14085_ _14085_/A _14085_/B vssd1 vssd1 vccd1 vccd1 _14201_/A sky130_fd_sc_hd__or2_1
X_13036_ _20673_/Q _13034_/X _12950_/X _13035_/X vssd1 vssd1 vccd1 vccd1 _20673_/D
+ sky130_fd_sc_hd__a22o_1
X_17913_ _20412_/Q vssd1 vssd1 vccd1 vccd1 _17913_/Y sky130_fd_sc_hd__inv_2
X_10248_ _21355_/Q vssd1 vssd1 vccd1 vccd1 _10270_/A sky130_fd_sc_hd__inv_2
X_18893_ _17182_/Y _14518_/A _18899_/S vssd1 vssd1 vccd1 vccd1 _18893_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17844_ _17844_/A vssd1 vssd1 vccd1 vccd1 _18064_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_227_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10179_ _10179_/A vssd1 vssd1 vccd1 vccd1 _10179_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17775_ _18674_/X _17775_/B vssd1 vssd1 vccd1 vccd1 _17775_/Y sky130_fd_sc_hd__nand2_1
XFILLER_82_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14987_ _14987_/A vssd1 vssd1 vccd1 vccd1 _14987_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_235_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16726_ _20988_/Q _11994_/B _11995_/B vssd1 vssd1 vccd1 vccd1 _16726_/X sky130_fd_sc_hd__a21bo_1
X_19514_ _19789_/CLK _19514_/D vssd1 vssd1 vccd1 vccd1 _19514_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_208_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13938_ _13935_/Y _20319_/Q _13936_/Y _20295_/Q _13937_/Y vssd1 vssd1 vccd1 vccd1
+ _13947_/B sky130_fd_sc_hd__o221a_1
XFILLER_223_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19445_ _19834_/CLK _19445_/D vssd1 vssd1 vccd1 vccd1 _19445_/Q sky130_fd_sc_hd__dfxtp_1
X_16657_ _16661_/A _18952_/X vssd1 vssd1 vccd1 vccd1 _19862_/D sky130_fd_sc_hd__and2_1
XFILLER_90_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13869_ _20291_/Q vssd1 vssd1 vccd1 vccd1 _14009_/A sky130_fd_sc_hd__inv_2
XFILLER_223_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15608_ _19718_/Q _15603_/X _15487_/X _15604_/X vssd1 vssd1 vccd1 vccd1 _19718_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_222_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19376_ _19706_/CLK _19376_/D vssd1 vssd1 vccd1 vccd1 _19376_/Q sky130_fd_sc_hd__dfxtp_1
X_16588_ _16588_/A vssd1 vssd1 vccd1 vccd1 _16588_/Y sky130_fd_sc_hd__inv_2
XFILLER_148_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18327_ _17812_/Y _20781_/Q _18885_/S vssd1 vssd1 vccd1 vccd1 _18327_/X sky130_fd_sc_hd__mux2_1
XFILLER_188_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15539_ _19752_/Q _15536_/X _15521_/X _15537_/X vssd1 vssd1 vccd1 vccd1 _19752_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_203_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18258_ _18257_/X _14592_/A _18748_/S vssd1 vssd1 vccd1 vccd1 _18258_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18082__B _18083_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17209_ _17209_/A vssd1 vssd1 vccd1 vccd1 _17889_/A sky130_fd_sc_hd__buf_1
XFILLER_191_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18189_ _18845_/A0 _13775_/Y _18896_/S vssd1 vssd1 vccd1 vccd1 _18189_/X sky130_fd_sc_hd__mux2_1
XFILLER_116_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20220_ _20220_/CLK _20220_/D repeater203/X vssd1 vssd1 vccd1 vccd1 _20220_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__20406__RESET_B repeater184/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13118__B1 _12991_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20151_ _21218_/CLK _20151_/D repeater250/X vssd1 vssd1 vccd1 vccd1 _20151_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_131_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09962_ _21422_/Q _09957_/X _09702_/X _09958_/X vssd1 vssd1 vccd1 vccd1 _21422_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17707__A _20504_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18302__S _18667_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20082_ _20590_/CLK _20082_/D repeater260/X vssd1 vssd1 vccd1 vccd1 _20082_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_131_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09893_ _20013_/Q vssd1 vssd1 vccd1 vccd1 _09893_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20984_ _21141_/CLK _20984_/D repeater191/X vssd1 vssd1 vccd1 vccd1 _20984_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_3905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11490__A _15847_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_241_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21467_ _21481_/CLK _21467_/D repeater205/X vssd1 vssd1 vccd1 vccd1 _21467_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_153_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14306__A _15574_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18296__A0 _18848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11220_ _11226_/A vssd1 vssd1 vccd1 vccd1 _11220_/X sky130_fd_sc_hd__buf_1
X_20418_ _20957_/CLK _20418_/D repeater187/X vssd1 vssd1 vccd1 vccd1 _20418_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__20147__RESET_B repeater242/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21398_ _21405_/CLK _21398_/D repeater253/X vssd1 vssd1 vccd1 vccd1 _21398_/Q sky130_fd_sc_hd__dfrtp_1
X_11151_ _11151_/A _11151_/B _11151_/C _11926_/A vssd1 vssd1 vccd1 vccd1 _11151_/X
+ sky130_fd_sc_hd__or4b_1
X_20349_ _20476_/CLK _20349_/D repeater280/X vssd1 vssd1 vccd1 vccd1 _20349_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__18212__S _18669_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10102_ _10155_/A _20791_/Q _21394_/Q _10099_/Y _10101_/X vssd1 vssd1 vccd1 vccd1
+ _10102_/X sky130_fd_sc_hd__a221o_1
X_11082_ _11101_/A vssd1 vssd1 vccd1 vccd1 _11082_/X sky130_fd_sc_hd__buf_1
XFILLER_0_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14910_ _20592_/Q vssd1 vssd1 vccd1 vccd1 _14910_/Y sky130_fd_sc_hd__inv_2
X_10033_ _21403_/Q vssd1 vssd1 vccd1 vccd1 _10034_/B sky130_fd_sc_hd__inv_2
XFILLER_209_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15890_ _19589_/Q _15886_/X _15887_/X _15889_/X vssd1 vssd1 vccd1 vccd1 _19589_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_103_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_248_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input24_A HADDR[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14841_ _20093_/Q vssd1 vssd1 vccd1 vccd1 _14961_/B sky130_fd_sc_hd__inv_2
XFILLER_217_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19043__S _19046_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17560_ _17560_/A vssd1 vssd1 vccd1 vccd1 _17560_/X sky130_fd_sc_hd__clkbuf_4
X_14772_ _19125_/X vssd1 vssd1 vccd1 vccd1 _14775_/A sky130_fd_sc_hd__inv_2
XFILLER_29_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11984_ _10994_/X _11910_/B _10994_/X _11910_/B vssd1 vssd1 vccd1 vccd1 _11984_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_84_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16511_ _20000_/Q vssd1 vssd1 vccd1 vccd1 _16511_/Y sky130_fd_sc_hd__inv_2
XFILLER_205_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13723_ _15762_/A _15764_/A _13725_/S vssd1 vssd1 vccd1 vccd1 _20329_/D sky130_fd_sc_hd__mux2_1
XFILLER_17_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10935_ _21208_/Q vssd1 vssd1 vccd1 vccd1 _10935_/Y sky130_fd_sc_hd__inv_2
X_17491_ _19410_/Q vssd1 vssd1 vccd1 vccd1 _17491_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18882__S _18910_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19230_ _17521_/Y _17522_/Y _17523_/Y _17524_/Y _20130_/Q _20131_/Q vssd1 vssd1 vccd1
+ vccd1 _19230_/X sky130_fd_sc_hd__mux4_2
XFILLER_32_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16442_ _16442_/A vssd1 vssd1 vccd1 vccd1 _16442_/X sky130_fd_sc_hd__buf_1
XFILLER_189_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13654_ _20366_/Q _13651_/X _13449_/X _13652_/X vssd1 vssd1 vccd1 vccd1 _20366_/D
+ sky130_fd_sc_hd__a22o_1
X_10866_ _10872_/A vssd1 vssd1 vccd1 vccd1 _10866_/X sky130_fd_sc_hd__buf_1
XFILLER_31_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13596__B1 _13446_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19161_ _19157_/X _19158_/X _19159_/X _19160_/X _21018_/Q _21019_/Q vssd1 vssd1 vccd1
+ vccd1 _19161_/X sky130_fd_sc_hd__mux4_2
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12605_ _12605_/A vssd1 vssd1 vccd1 vccd1 _12606_/A sky130_fd_sc_hd__buf_1
XANTENNA__20917__RESET_B repeater218/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13104__B _13104_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16373_ _19351_/Q _16370_/X _16210_/X _16371_/X vssd1 vssd1 vccd1 vccd1 _19351_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13585_ _20406_/Q _13580_/X _13584_/X _13581_/X vssd1 vssd1 vccd1 vccd1 _20406_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_repeater163_A _18910_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10797_ _10797_/A vssd1 vssd1 vccd1 vccd1 _10797_/Y sky130_fd_sc_hd__inv_2
XFILLER_200_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18112_ _18112_/A _18112_/B vssd1 vssd1 vccd1 vccd1 _18112_/Y sky130_fd_sc_hd__nor2_8
XFILLER_200_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15324_ _15330_/A vssd1 vssd1 vccd1 vccd1 _15324_/X sky130_fd_sc_hd__buf_1
X_12536_ _12527_/A _12525_/Y _19989_/Q _11299_/A _12520_/X vssd1 vssd1 vccd1 vccd1
+ _20906_/D sky130_fd_sc_hd__a32o_1
X_19092_ _16678_/X _21086_/Q _19870_/D vssd1 vssd1 vccd1 vccd1 _19092_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17731__C1 _17730_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13348__B1 _13209_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18043_ _20836_/Q vssd1 vssd1 vccd1 vccd1 _18043_/Y sky130_fd_sc_hd__inv_2
XFILLER_184_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15255_ _20488_/Q vssd1 vssd1 vccd1 vccd1 _15255_/Y sky130_fd_sc_hd__inv_2
X_12467_ _12419_/A _12419_/B _12465_/Y _12496_/C vssd1 vssd1 vccd1 vccd1 _20930_/D
+ sky130_fd_sc_hd__a211oi_4
XANTENNA_output92_A _17999_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14206_ _20274_/Q _14204_/Y _14205_/X _14085_/B vssd1 vssd1 vccd1 vccd1 _20274_/D
+ sky130_fd_sc_hd__o211a_1
X_11418_ _11418_/A vssd1 vssd1 vccd1 vccd1 _11418_/X sky130_fd_sc_hd__buf_1
X_15186_ _15098_/X _15184_/Y _15185_/X _15078_/B vssd1 vssd1 vccd1 vccd1 _20063_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_99_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12398_ _12475_/A _12474_/A _12398_/C _12476_/A vssd1 vssd1 vccd1 vccd1 _12399_/D
+ sky130_fd_sc_hd__or4_4
XANTENNA__12571__A1 _17169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12571__B2 _18242_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14137_ _14133_/Y _20277_/Q _20536_/Q _14076_/A _14136_/X vssd1 vssd1 vccd1 vccd1
+ _14138_/D sky130_fd_sc_hd__o221a_1
XFILLER_126_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11349_ _21179_/Q _21178_/Q _11362_/B vssd1 vssd1 vccd1 vccd1 _11366_/C sky130_fd_sc_hd__or3_1
X_19994_ _21055_/CLK _19994_/D repeater220/X vssd1 vssd1 vccd1 vccd1 _19994_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_141_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18945_ _16692_/X _20896_/Q _18946_/S vssd1 vssd1 vccd1 vccd1 _18945_/X sky130_fd_sc_hd__mux2_1
X_14068_ _20260_/Q vssd1 vssd1 vccd1 vccd1 _14071_/A sky130_fd_sc_hd__inv_2
XFILLER_113_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_100_HCLK clkbuf_4_13_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20322_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_239_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13019_ _13040_/A vssd1 vssd1 vccd1 vccd1 _13019_/X sky130_fd_sc_hd__buf_1
XFILLER_239_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18876_ _17190_/Y _16758_/A _18899_/S vssd1 vssd1 vccd1 vccd1 _18876_/X sky130_fd_sc_hd__mux2_1
XFILLER_227_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17827_ _17827_/A _17827_/B _17827_/C vssd1 vssd1 vccd1 vccd1 _17827_/X sky130_fd_sc_hd__and3_2
X_17758_ _19453_/Q vssd1 vssd1 vccd1 vccd1 _17758_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18211__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18077__B _18078_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16709_ _16709_/A _18938_/X vssd1 vssd1 vccd1 vccd1 _19898_/D sky130_fd_sc_hd__and2_1
X_17689_ _19347_/Q vssd1 vssd1 vccd1 vccd1 _17689_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18792__S _18927_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19428_ _20331_/CLK _19428_/D vssd1 vssd1 vccd1 vccd1 _19428_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17970__C1 _17969_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13587__B1 _13586_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19359_ _19521_/CLK _19359_/D vssd1 vssd1 vccd1 vccd1 _19359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15328__A1 _20028_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21321_ _21321_/CLK _21321_/D repeater205/X vssd1 vssd1 vccd1 vccd1 _21321_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_148_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21252_ _21438_/CLK _21252_/D repeater239/X vssd1 vssd1 vccd1 vccd1 _21252_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_116_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20203_ _20626_/CLK _20203_/D repeater193/X vssd1 vssd1 vccd1 vccd1 _20203_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_145_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21183_ _21183_/CLK _21183_/D repeater216/X vssd1 vssd1 vccd1 vccd1 _21183_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20134_ _20241_/CLK _20134_/D repeater248/X vssd1 vssd1 vccd1 vccd1 _20134_/Q sky130_fd_sc_hd__dfrtp_1
X_09945_ _20871_/Q vssd1 vssd1 vccd1 vccd1 _10877_/A sky130_fd_sc_hd__buf_1
XFILLER_131_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__21446__RESET_B repeater248/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20065_ _20070_/CLK _20065_/D hold8/X vssd1 vssd1 vccd1 vccd1 _20065_/Q sky130_fd_sc_hd__dfrtp_2
X_09876_ _09876_/A _09878_/A _09878_/B vssd1 vssd1 vccd1 vccd1 _09876_/X sky130_fd_sc_hd__or3_2
XFILLER_161_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrepeater260 repeater267/X vssd1 vssd1 vccd1 vccd1 repeater260/X sky130_fd_sc_hd__buf_8
Xrepeater271 repeater272/X vssd1 vssd1 vccd1 vccd1 repeater271/X sky130_fd_sc_hd__clkbuf_8
XFILLER_100_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18202__A0 _18848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10628__B2 _10626_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20967_ _20971_/CLK _20967_/D repeater186/X vssd1 vssd1 vccd1 vccd1 _20967_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_3735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10720_ _10720_/A vssd1 vssd1 vccd1 vccd1 _10725_/A sky130_fd_sc_hd__inv_2
XFILLER_198_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20898_ _21141_/CLK _20898_/D repeater212/X vssd1 vssd1 vccd1 vccd1 _20898_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__13578__B1 _13424_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10651_ _10651_/A _10651_/B vssd1 vssd1 vccd1 vccd1 _10697_/A sky130_fd_sc_hd__or2_1
XFILLER_13_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20399__RESET_B repeater270/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18207__S _18907_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20328__RESET_B repeater190/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10582_ _10543_/A _20744_/Q _10664_/C _20764_/Q _10581_/X vssd1 vssd1 vccd1 vccd1
+ _10591_/B sky130_fd_sc_hd__o221a_1
XFILLER_155_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13370_ _20506_/Q _13365_/X _13313_/X _13366_/X vssd1 vssd1 vccd1 vccd1 _20506_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_221_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12321_ _12321_/A _12321_/B vssd1 vssd1 vccd1 vccd1 _12358_/A sky130_fd_sc_hd__or2_1
XFILLER_127_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15040_ _20062_/Q vssd1 vssd1 vccd1 vccd1 _15076_/A sky130_fd_sc_hd__inv_2
X_12252_ _20521_/Q vssd1 vssd1 vccd1 vccd1 _12252_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_123_HCLK clkbuf_4_4_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20981_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_107_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19038__S _19046_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11203_ _16488_/A vssd1 vssd1 vccd1 vccd1 _14702_/A sky130_fd_sc_hd__buf_2
XFILLER_108_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12183_ _20339_/Q vssd1 vssd1 vccd1 vccd1 _12183_/Y sky130_fd_sc_hd__inv_2
X_11134_ _21219_/Q vssd1 vssd1 vccd1 vccd1 _15466_/B sky130_fd_sc_hd__inv_2
XFILLER_122_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16991_ _19975_/Q vssd1 vssd1 vccd1 vccd1 _16994_/A sky130_fd_sc_hd__inv_2
XANTENNA__18877__S _18910_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13502__B1 _13432_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15942_ _19562_/Q _15935_/X _15941_/X _15937_/X vssd1 vssd1 vccd1 vccd1 _19562_/D
+ sky130_fd_sc_hd__a22o_1
X_11065_ _11100_/A vssd1 vssd1 vccd1 vccd1 _11066_/B sky130_fd_sc_hd__inv_2
X_18730_ _18729_/X _12223_/Y _18910_/S vssd1 vssd1 vccd1 vccd1 _18730_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10016_ _09996_/Y _09998_/Y _21419_/Q _17036_/A _10015_/X vssd1 vssd1 vccd1 vccd1
+ _10016_/X sky130_fd_sc_hd__o221a_1
XANTENNA__21116__RESET_B repeater233/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18661_ _18077_/Y _20361_/Q _18909_/S vssd1 vssd1 vccd1 vccd1 _18661_/X sky130_fd_sc_hd__mux2_1
XANTENNA_output130_A _20003_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15873_ _15873_/A vssd1 vssd1 vccd1 vccd1 _15873_/X sky130_fd_sc_hd__buf_1
XFILLER_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17795__A2 _17141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17612_ _19451_/Q vssd1 vssd1 vccd1 vccd1 _17612_/Y sky130_fd_sc_hd__inv_2
X_14824_ _20562_/Q vssd1 vssd1 vccd1 vccd1 _14824_/Y sky130_fd_sc_hd__inv_2
X_18592_ _18591_/X _10593_/Y _18879_/S vssd1 vssd1 vccd1 vccd1 _18592_/X sky130_fd_sc_hd__mux2_1
XFILLER_224_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17543_ _17808_/A vssd1 vssd1 vccd1 vccd1 _17807_/B sky130_fd_sc_hd__buf_4
X_14755_ _20133_/Q vssd1 vssd1 vccd1 vccd1 _14755_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_repeater280_A repeater281/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11967_ _20597_/Q vssd1 vssd1 vccd1 vccd1 _13182_/B sky130_fd_sc_hd__buf_1
XFILLER_91_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13706_ _13706_/A vssd1 vssd1 vccd1 vccd1 _13706_/X sky130_fd_sc_hd__buf_1
X_17474_ _17474_/A vssd1 vssd1 vccd1 vccd1 _17474_/X sky130_fd_sc_hd__buf_1
X_10918_ _10918_/A _10918_/B vssd1 vssd1 vccd1 vccd1 _12735_/A sky130_fd_sc_hd__or2_2
X_14686_ _14686_/A _14686_/B vssd1 vssd1 vccd1 vccd1 _16526_/B sky130_fd_sc_hd__or2_2
XFILLER_60_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11898_ _10994_/X _11897_/A _10993_/Y _11900_/A vssd1 vssd1 vccd1 vccd1 _21019_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_232_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16425_ _19322_/Q _16420_/X _15871_/A _16422_/X vssd1 vssd1 vccd1 vccd1 _19322_/D
+ sky130_fd_sc_hd__a22o_1
X_19213_ _17670_/Y _17671_/Y _17672_/Y _17673_/Y _19275_/S0 _21004_/Q vssd1 vssd1
+ vccd1 vccd1 _19213_/X sky130_fd_sc_hd__mux4_2
XANTENNA__20751__RESET_B repeater210/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13637_ _20377_/Q _13632_/X _13424_/X _13634_/X vssd1 vssd1 vccd1 vccd1 _20377_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_220_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10849_ _10849_/A vssd1 vssd1 vccd1 vccd1 _10849_/X sky130_fd_sc_hd__buf_1
XANTENNA__12954__A _14262_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15330__A _15330_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19144_ _19689_/Q _19377_/Q _19673_/Q _19665_/Q _19285_/S0 _21017_/Q vssd1 vssd1
+ vccd1 vccd1 _19144_/X sky130_fd_sc_hd__mux4_1
XANTENNA__20069__RESET_B repeater276/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16356_ _19359_/Q _16352_/X _16293_/X _16353_/X vssd1 vssd1 vccd1 vccd1 _19359_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_185_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13568_ _20416_/Q _13566_/X _13482_/X _13567_/X vssd1 vssd1 vccd1 vccd1 _20416_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09966__C _12605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15307_ _20039_/Q _15302_/X _20038_/Q _15305_/X vssd1 vssd1 vccd1 vccd1 _20039_/D
+ sky130_fd_sc_hd__a22o_1
X_12519_ _20916_/Q _12521_/A _12502_/B _12518_/X vssd1 vssd1 vccd1 vccd1 _20916_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_185_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19075_ _16728_/X _20900_/Q _19908_/D vssd1 vssd1 vccd1 vccd1 _19075_/X sky130_fd_sc_hd__mux2_1
XFILLER_157_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16287_ _16287_/A vssd1 vssd1 vccd1 vccd1 _16287_/X sky130_fd_sc_hd__buf_1
X_13499_ _13514_/A vssd1 vssd1 vccd1 vccd1 _13499_/X sky130_fd_sc_hd__buf_1
XFILLER_246_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18026_ _18261_/X _18024_/X _18323_/X _17995_/X _18025_/X vssd1 vssd1 vccd1 vccd1
+ _18027_/C sky130_fd_sc_hd__o221a_1
X_15238_ _20493_/Q vssd1 vssd1 vccd1 vccd1 _15238_/Y sky130_fd_sc_hd__inv_2
XFILLER_173_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15169_ _15169_/A vssd1 vssd1 vccd1 vccd1 _15169_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19977_ _20809_/CLK _19977_/D repeater188/X vssd1 vssd1 vccd1 vccd1 _19977_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18787__S _18787_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09730_ _21234_/Q vssd1 vssd1 vccd1 vccd1 _11059_/A sky130_fd_sc_hd__inv_2
XFILLER_113_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18928_ _18927_/X _10933_/Y _18928_/S vssd1 vssd1 vccd1 vccd1 _18928_/X sky130_fd_sc_hd__mux2_1
X_09661_ _21473_/Q _09657_/X _09659_/X _09660_/X vssd1 vssd1 vccd1 vccd1 _21473_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_83_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18859_ _17279_/X _21251_/Q _20870_/Q vssd1 vssd1 vccd1 vccd1 _18859_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19934__RESET_B repeater251/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17786__A2 _17141_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20821_ _21401_/CLK _20821_/D repeater256/X vssd1 vssd1 vccd1 vccd1 _20821_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_208_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18735__A1 _19221_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20752_ _21294_/CLK _20752_/D repeater209/X vssd1 vssd1 vccd1 vccd1 _20752_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_35_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20683_ _21302_/CLK _20683_/D repeater208/X vssd1 vssd1 vccd1 vccd1 _20683_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18499__A0 _17079_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_146_HCLK clkbuf_opt_1_HCLK/A vssd1 vssd1 vccd1 vccd1 _20241_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_40_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14509__C1 _14469_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21304_ _21306_/CLK _21304_/D repeater206/X vssd1 vssd1 vccd1 vccd1 _21304_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__19739__CLK _19765_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21235_ _21235_/CLK _21235_/D repeater189/X vssd1 vssd1 vccd1 vccd1 _21235_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_105_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21166_ _21167_/CLK _21166_/D repeater225/X vssd1 vssd1 vccd1 vccd1 _21166_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_78_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18697__S _18907_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14303__B _20889_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__21280__RESET_B repeater207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20117_ _21453_/CLK _20117_/D repeater247/X vssd1 vssd1 vccd1 vccd1 _20117_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_104_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09928_ _21431_/Q _21432_/Q _09929_/S vssd1 vssd1 vccd1 vccd1 _21432_/D sky130_fd_sc_hd__mux2_1
X_21097_ _21423_/CLK _21097_/D repeater231/X vssd1 vssd1 vccd1 vccd1 _21097_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_246_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18423__A0 _17079_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20048_ _20470_/CLK _20048_/D repeater280/X vssd1 vssd1 vccd1 vccd1 _20048_/Q sky130_fd_sc_hd__dfrtp_1
X_09859_ _09859_/A _09859_/B vssd1 vssd1 vccd1 vccd1 _09859_/Y sky130_fd_sc_hd__nor2_1
XFILLER_92_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12870_ _20744_/Q _12867_/X _12548_/X _12868_/X vssd1 vssd1 vccd1 vccd1 _20744_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_65_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11821_ _11827_/A vssd1 vssd1 vccd1 vccd1 _11822_/B sky130_fd_sc_hd__clkbuf_2
XPHY_4244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14540_ _15902_/B vssd1 vssd1 vccd1 vccd1 _14541_/A sky130_fd_sc_hd__buf_1
XFILLER_242_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11752_ _19873_/Q vssd1 vssd1 vccd1 vccd1 _11753_/C sky130_fd_sc_hd__inv_2
XPHY_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10703_ _10703_/A _10718_/A vssd1 vssd1 vccd1 vccd1 _10704_/B sky130_fd_sc_hd__or2_1
XFILLER_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14471_ _14471_/A vssd1 vssd1 vccd1 vccd1 _14471_/Y sky130_fd_sc_hd__inv_2
XPHY_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11683_ _21087_/Q _11679_/X _11680_/X _11682_/X vssd1 vssd1 vccd1 vccd1 _21087_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16210_ _21448_/Q vssd1 vssd1 vccd1 vccd1 _16210_/X sky130_fd_sc_hd__buf_1
XPHY_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13422_ input43/X vssd1 vssd1 vccd1 vccd1 _13422_/X sky130_fd_sc_hd__clkbuf_2
X_10634_ _20765_/Q vssd1 vssd1 vccd1 vccd1 _10634_/Y sky130_fd_sc_hd__inv_2
X_17190_ _20772_/Q _17193_/B vssd1 vssd1 vccd1 vccd1 _17190_/Y sky130_fd_sc_hd__nor2_1
XPHY_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12774__A1 _20795_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16141_ _16141_/A vssd1 vssd1 vccd1 vccd1 _16141_/X sky130_fd_sc_hd__buf_1
XFILLER_6_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13353_ _20517_/Q _13351_/X _13216_/X _13352_/X vssd1 vssd1 vccd1 vccd1 _20517_/D
+ sky130_fd_sc_hd__a22o_1
X_10565_ _10657_/A _10656_/A _10658_/A _10655_/A vssd1 vssd1 vccd1 vccd1 _10566_/D
+ sky130_fd_sc_hd__or4_4
XFILLER_10_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12304_ _12304_/A _12410_/A vssd1 vssd1 vccd1 vccd1 _12389_/A sky130_fd_sc_hd__or2_2
XFILLER_5_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16072_ _16072_/A vssd1 vssd1 vccd1 vccd1 _16072_/X sky130_fd_sc_hd__clkbuf_2
X_13284_ input54/X vssd1 vssd1 vccd1 vccd1 _13284_/X sky130_fd_sc_hd__clkbuf_2
X_10496_ _10496_/A _10496_/B _10496_/C _10496_/D vssd1 vssd1 vccd1 vccd1 _10523_/C
+ sky130_fd_sc_hd__and4_1
X_19900_ _21193_/CLK _19900_/D repeater224/X vssd1 vssd1 vccd1 vccd1 _19900_/Q sky130_fd_sc_hd__dfrtp_1
X_15023_ _14853_/B _15022_/A _20078_/Q _15025_/A _14958_/X vssd1 vssd1 vccd1 vccd1
+ _20078_/D sky130_fd_sc_hd__o221a_1
XANTENNA__21368__RESET_B repeater257/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12235_ _20927_/Q vssd1 vssd1 vccd1 vccd1 _12475_/A sky130_fd_sc_hd__inv_2
XANTENNA__20396__CLK _20930_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19831_ _19834_/CLK _19831_/D vssd1 vssd1 vccd1 vccd1 _19831_/Q sky130_fd_sc_hd__dfxtp_1
X_12166_ _20968_/Q _20350_/Q _12321_/A _12165_/Y vssd1 vssd1 vccd1 vccd1 _12166_/X
+ sky130_fd_sc_hd__o22a_1
X_11117_ _11112_/X _11113_/X _09739_/X vssd1 vssd1 vccd1 vccd1 _11117_/X sky130_fd_sc_hd__o21a_1
X_19762_ _21009_/CLK _19762_/D vssd1 vssd1 vccd1 vccd1 _19762_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_19_HCLK_A clkbuf_4_3_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16974_ _17013_/A _16974_/B vssd1 vssd1 vccd1 vccd1 _16974_/Y sky130_fd_sc_hd__nor2_1
X_12097_ _12312_/A vssd1 vssd1 vccd1 vccd1 _12097_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__18400__S _18879_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_237_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18414__A0 _17281_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_27_HCLK clkbuf_opt_4_HCLK/A vssd1 vssd1 vccd1 vccd1 _21417_/CLK sky130_fd_sc_hd__clkbuf_16
X_18713_ _18845_/A0 _10303_/Y _18884_/S vssd1 vssd1 vccd1 vccd1 _18713_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15925_ _19571_/Q _15920_/X _15893_/X _15922_/X vssd1 vssd1 vccd1 vccd1 _19571_/D
+ sky130_fd_sc_hd__a22o_1
X_11048_ _17027_/A _21240_/Q _21241_/Q vssd1 vssd1 vccd1 vccd1 _21240_/D sky130_fd_sc_hd__a21o_1
X_19693_ _19813_/CLK _19693_/D vssd1 vssd1 vccd1 vccd1 _19693_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_7_HCLK_A clkbuf_opt_2_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15228__B1 _17896_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput8 HADDR[16] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__clkbuf_1
XFILLER_76_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15856_ _15856_/A vssd1 vssd1 vccd1 vccd1 _15856_/X sky130_fd_sc_hd__buf_1
X_18644_ _18643_/X _10119_/Y _18644_/S vssd1 vssd1 vccd1 vccd1 _18644_/X sky130_fd_sc_hd__mux2_1
XFILLER_80_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14807_ _19125_/S _14807_/B vssd1 vssd1 vccd1 vccd1 _14807_/X sky130_fd_sc_hd__or2_2
XFILLER_224_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15787_ _15787_/A vssd1 vssd1 vccd1 vccd1 _15787_/X sky130_fd_sc_hd__buf_1
X_18575_ _18574_/X _17849_/Y _18903_/S vssd1 vssd1 vccd1 vccd1 _18575_/X sky130_fd_sc_hd__mux2_1
XFILLER_51_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12999_ input56/X vssd1 vssd1 vccd1 vccd1 _12999_/X sky130_fd_sc_hd__buf_2
X_17526_ _14795_/Y _19334_/Q _17525_/X vssd1 vssd1 vccd1 vccd1 _17526_/Y sky130_fd_sc_hd__o21ai_1
X_14738_ _20139_/Q _14732_/A _13714_/X _14733_/A vssd1 vssd1 vccd1 vccd1 _20139_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_33_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_169_HCLK clkbuf_opt_0_HCLK/A vssd1 vssd1 vccd1 vccd1 _21461_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_44_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17457_ _21067_/Q vssd1 vssd1 vccd1 vccd1 _17457_/Y sky130_fd_sc_hd__inv_2
X_14669_ _14659_/A _14659_/B _14660_/A _14663_/Y vssd1 vssd1 vccd1 vccd1 _14669_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_189_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16408_ _16414_/A vssd1 vssd1 vccd1 vccd1 _16408_/X sky130_fd_sc_hd__buf_1
X_17388_ _20246_/Q vssd1 vssd1 vccd1 vccd1 _17388_/Y sky130_fd_sc_hd__inv_2
XFILLER_118_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16339_ _19368_/Q _16334_/X _16338_/X _16336_/X vssd1 vssd1 vccd1 vccd1 _19368_/D
+ sky130_fd_sc_hd__a22o_1
X_19127_ _19678_/Q _19806_/Q _19798_/Q _19790_/Q _19285_/S0 _21017_/Q vssd1 vssd1
+ vccd1 vccd1 _19127_/X sky130_fd_sc_hd__mux4_2
XFILLER_118_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19058_ _16748_/Y _20811_/Q _19058_/S vssd1 vssd1 vccd1 vccd1 _19918_/D sky130_fd_sc_hd__mux2_1
XANTENNA__15164__C1 _15201_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18090__B _18090_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18009_ _20419_/Q _18084_/B vssd1 vssd1 vccd1 vccd1 _18009_/Y sky130_fd_sc_hd__nand2_1
XFILLER_160_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18102__C1 _18101_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21038__RESET_B repeater242/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21020_ _21021_/CLK _21020_/D repeater238/X vssd1 vssd1 vccd1 vccd1 _21020_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_114_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17715__A _21086_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18310__S _18897_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09713_ _21454_/Q vssd1 vssd1 vccd1 vccd1 _09803_/A sky130_fd_sc_hd__inv_2
XANTENNA__17208__B2 _17203_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18956__A1 _21080_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20119__CLK _21452_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09644_ input43/X vssd1 vssd1 vccd1 vccd1 _12853_/A sky130_fd_sc_hd__buf_4
XFILLER_216_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20804_ _21407_/CLK _20804_/D repeater252/X vssd1 vssd1 vccd1 vccd1 _20804_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_224_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16719__B1 _18946_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20735_ _21294_/CLK _20735_/D repeater210/X vssd1 vssd1 vccd1 vccd1 _20735_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20666_ _21306_/CLK _20666_/D repeater207/X vssd1 vssd1 vccd1 vccd1 _20666_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13953__B1 _13951_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20597_ _21011_/CLK _20597_/D repeater235/X vssd1 vssd1 vccd1 vccd1 _20597_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_192_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10350_ _10280_/A _20724_/Q _10346_/X _20712_/Q _10349_/X vssd1 vssd1 vccd1 vccd1
+ _10360_/B sky130_fd_sc_hd__o221a_1
XFILLER_109_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21461__RESET_B repeater245/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13705__B1 _13704_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10281_ _10281_/A _10281_/B vssd1 vssd1 vccd1 vccd1 _10380_/A sky130_fd_sc_hd__or2_1
XFILLER_105_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12020_ _19072_/X _12017_/X _20993_/Q _12018_/X vssd1 vssd1 vccd1 vccd1 _20993_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_3_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21218_ _21218_/CLK _21218_/D repeater242/X vssd1 vssd1 vccd1 vccd1 _21218_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__15458__B1 _15421_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21149_ _21151_/CLK _21149_/D repeater223/X vssd1 vssd1 vccd1 vccd1 _21149_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18220__S _18236_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13971_ _13971_/A _13971_/B _13971_/C _13971_/D vssd1 vssd1 vccd1 vccd1 _13972_/D
+ sky130_fd_sc_hd__or4_1
XFILLER_93_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15710_ _15716_/A vssd1 vssd1 vccd1 vccd1 _15717_/A sky130_fd_sc_hd__inv_2
XFILLER_246_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12922_ input50/X vssd1 vssd1 vccd1 vccd1 _12922_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_86_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16690_ _20895_/Q vssd1 vssd1 vccd1 vccd1 _16690_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12692__B1 _09652_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15641_ _15647_/A vssd1 vssd1 vccd1 vccd1 _15648_/A sky130_fd_sc_hd__inv_2
X_12853_ _12853_/A vssd1 vssd1 vccd1 vccd1 _12853_/X sky130_fd_sc_hd__clkbuf_2
XPHY_4030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19051__S _19058_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15630__B1 _15550_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18360_ _18848_/A0 _18053_/Y _18666_/S vssd1 vssd1 vccd1 vccd1 _18360_/X sky130_fd_sc_hd__mux2_1
X_11804_ _11863_/A _11864_/A _11804_/C _11804_/D vssd1 vssd1 vccd1 vccd1 _11859_/A
+ sky130_fd_sc_hd__or4_4
XPHY_4074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15572_ _19735_/Q _15568_/X _15524_/X _15569_/X vssd1 vssd1 vccd1 vccd1 _19735_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12784_ _12803_/A vssd1 vssd1 vccd1 vccd1 _12784_/X sky130_fd_sc_hd__buf_1
XFILLER_221_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19904__CLK _19904_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17311_ _18858_/X vssd1 vssd1 vccd1 vccd1 _17311_/Y sky130_fd_sc_hd__inv_2
X_14523_ _14518_/A _14518_/B _14518_/C vssd1 vssd1 vccd1 vccd1 _14524_/B sky130_fd_sc_hd__o21a_1
XPHY_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11735_ _11735_/A vssd1 vssd1 vccd1 vccd1 _11735_/X sky130_fd_sc_hd__buf_1
X_18291_ _17975_/Y _20352_/Q _18787_/S vssd1 vssd1 vccd1 vccd1 _18291_/X sky130_fd_sc_hd__mux2_1
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_202_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18890__S _18896_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17242_ _19391_/Q vssd1 vssd1 vccd1 vccd1 _17242_/Y sky130_fd_sc_hd__inv_2
XPHY_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14454_ _20240_/Q _14383_/Y _14384_/Y _14383_/A _14453_/X vssd1 vssd1 vccd1 vccd1
+ _20240_/D sky130_fd_sc_hd__o221a_1
XFILLER_159_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11666_ _21071_/Q vssd1 vssd1 vccd1 vccd1 _16634_/A sky130_fd_sc_hd__inv_2
XPHY_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13405_ _13411_/A vssd1 vssd1 vccd1 vccd1 _13405_/X sky130_fd_sc_hd__buf_1
XPHY_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10617_ _21336_/Q _10614_/Y _10702_/A _20742_/Q _10616_/X vssd1 vssd1 vccd1 vccd1
+ _10622_/C sky130_fd_sc_hd__o221a_1
X_17173_ _20396_/Q _17174_/B vssd1 vssd1 vccd1 vccd1 _17173_/Y sky130_fd_sc_hd__nor2_1
X_14385_ _21482_/Q vssd1 vssd1 vccd1 vccd1 _14385_/Y sky130_fd_sc_hd__inv_2
XPHY_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11597_ _11599_/A vssd1 vssd1 vccd1 vccd1 _11598_/A sky130_fd_sc_hd__buf_1
X_16124_ _19472_/Q _16119_/X _16123_/X _16121_/X vssd1 vssd1 vccd1 vccd1 _19472_/D
+ sky130_fd_sc_hd__a22o_1
X_13336_ _20528_/Q _13331_/X _13270_/X _13334_/X vssd1 vssd1 vccd1 vccd1 _20528_/D
+ sky130_fd_sc_hd__a22o_1
X_10548_ _21318_/Q vssd1 vssd1 vccd1 vccd1 _10706_/A sky130_fd_sc_hd__inv_2
XFILLER_6_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16055_ _19506_/Q _16049_/X _15766_/X _16051_/X vssd1 vssd1 vccd1 vccd1 _19506_/D
+ sky130_fd_sc_hd__a22o_1
X_13267_ _13301_/A vssd1 vssd1 vccd1 vccd1 _13294_/A sky130_fd_sc_hd__buf_1
X_10479_ _20669_/Q vssd1 vssd1 vccd1 vccd1 _10479_/Y sky130_fd_sc_hd__inv_2
XFILLER_142_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15006_ _15006_/A _15006_/B vssd1 vssd1 vccd1 vccd1 _15006_/Y sky130_fd_sc_hd__nor2_1
X_12218_ _12490_/C _20499_/Q _12430_/A _20521_/Q vssd1 vssd1 vccd1 vccd1 _12218_/X
+ sky130_fd_sc_hd__o22a_1
X_13198_ _20594_/Q _13192_/X _12991_/X _13195_/X vssd1 vssd1 vccd1 vccd1 _20594_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_96_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19814_ _20172_/CLK _19814_/D vssd1 vssd1 vccd1 vccd1 _19814_/Q sky130_fd_sc_hd__dfxtp_1
X_12149_ _20953_/Q _12146_/Y _12073_/X _12147_/Y _12148_/X vssd1 vssd1 vccd1 vccd1
+ _12159_/A sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_143_HCLK_A clkbuf_4_3_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18130__S _18910_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19745_ _21121_/CLK _19745_/D vssd1 vssd1 vccd1 vccd1 _19745_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16957_ _19968_/Q vssd1 vssd1 vccd1 vccd1 _16957_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18938__A1 _21138_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15908_ _19580_/Q _15904_/X _15869_/X _15906_/X vssd1 vssd1 vccd1 vccd1 _19580_/D
+ sky130_fd_sc_hd__a22o_1
X_19676_ _19812_/CLK _19676_/D vssd1 vssd1 vccd1 vccd1 _19676_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12683__B1 _09636_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16888_ _19950_/Q vssd1 vssd1 vccd1 vccd1 _16889_/B sky130_fd_sc_hd__inv_2
XFILLER_92_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18627_ _18626_/X _21373_/Q _18841_/S vssd1 vssd1 vccd1 vccd1 _18627_/X sky130_fd_sc_hd__mux2_1
X_15839_ _19611_/Q _15834_/X _09824_/X _15836_/X vssd1 vssd1 vccd1 vccd1 _19611_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_53_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18558_ _17281_/X _17867_/Y _18835_/S vssd1 vssd1 vccd1 vccd1 _18558_/X sky130_fd_sc_hd__mux2_1
X_17509_ _19482_/Q vssd1 vssd1 vccd1 vccd1 _17509_/Y sky130_fd_sc_hd__inv_2
X_18489_ _18488_/X _14902_/Y _18907_/S vssd1 vssd1 vccd1 vccd1 _18489_/X sky130_fd_sc_hd__mux2_2
XFILLER_166_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20520_ _20937_/CLK _20520_/D repeater275/X vssd1 vssd1 vccd1 vccd1 _20520_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__20561__CLK _20592_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20451_ _20476_/CLK _20451_/D repeater183/X vssd1 vssd1 vccd1 vccd1 _20451_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_158_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18305__S _18907_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19210__S1 _20131_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21219__RESET_B repeater235/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20382_ _20480_/CLK _20382_/D repeater183/X vssd1 vssd1 vccd1 vccd1 _20382_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_134_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput120 _18113_/X vssd1 vssd1 vccd1 vccd1 IRQ[2] sky130_fd_sc_hd__clkbuf_2
XANTENNA__14134__A _20540_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput131 _20004_/Q vssd1 vssd1 vccd1 vccd1 RsTx_S1 sky130_fd_sc_hd__clkbuf_2
XFILLER_133_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput142 _18123_/LO vssd1 vssd1 vccd1 vccd1 sda_o_S4 sky130_fd_sc_hd__clkbuf_2
XFILLER_133_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21003_ _21009_/CLK _21003_/D repeater235/X vssd1 vssd1 vccd1 vccd1 _21003_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_153_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20854__RESET_B repeater243/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19277__S1 _20122_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15860__B1 _15793_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_65_HCLK_A clkbuf_4_11_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09627_ _21484_/Q _09620_/X _09626_/X _09624_/X vssd1 vssd1 vccd1 vccd1 _21484_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_16_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12977__A1 _20699_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14309__A _14309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11520_ _15354_/A vssd1 vssd1 vccd1 vccd1 _11520_/Y sky130_fd_sc_hd__inv_2
XPHY_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13213__A input50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20718_ _20724_/CLK _20718_/D repeater254/X vssd1 vssd1 vccd1 vccd1 _20718_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_8_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13926__B1 _20663_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11451_ _21163_/Q _11451_/B vssd1 vssd1 vccd1 vccd1 _11452_/B sky130_fd_sc_hd__or2_1
XPHY_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20649_ _21486_/CLK _20649_/D repeater198/X vssd1 vssd1 vccd1 vccd1 _20649_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_165_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19201__S1 _20133_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18215__S _18903_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10402_ _10402_/A vssd1 vssd1 vccd1 vccd1 _10405_/A sky130_fd_sc_hd__inv_2
X_14170_ _14170_/A _14170_/B _14170_/C _14170_/D vssd1 vssd1 vccd1 vccd1 _14171_/D
+ sky130_fd_sc_hd__and4_1
X_11382_ _21169_/Q vssd1 vssd1 vccd1 vccd1 _11385_/A sky130_fd_sc_hd__clkbuf_2
X_13121_ _13133_/A vssd1 vssd1 vccd1 vccd1 _13121_/X sky130_fd_sc_hd__buf_1
X_10333_ _20729_/Q vssd1 vssd1 vccd1 vccd1 _10333_/Y sky130_fd_sc_hd__inv_2
XFILLER_194_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input54_A HWDATA[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13052_ _13072_/A vssd1 vssd1 vccd1 vccd1 _13052_/X sky130_fd_sc_hd__buf_1
X_10264_ _10264_/A _10264_/B vssd1 vssd1 vccd1 vccd1 _10412_/A sky130_fd_sc_hd__or2_1
X_12003_ _20997_/Q _12003_/B vssd1 vssd1 vccd1 vccd1 _12003_/X sky130_fd_sc_hd__or2_2
XANTENNA__19046__S _19046_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18093__B2 _17861_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17860_ _18578_/X _17856_/X _18564_/X _17569_/X _17859_/X vssd1 vssd1 vccd1 vccd1
+ _17860_/X sky130_fd_sc_hd__o221a_1
X_10195_ _10151_/A _10151_/B _10185_/X _10193_/Y vssd1 vssd1 vccd1 vccd1 _21390_/D
+ sky130_fd_sc_hd__a211oi_2
X_16811_ _16815_/B _16810_/X _16803_/X vssd1 vssd1 vccd1 vccd1 _16811_/X sky130_fd_sc_hd__o21a_1
XANTENNA__20595__RESET_B repeater259/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17791_ _17789_/Y _17139_/A _17790_/Y _17136_/A vssd1 vssd1 vccd1 vccd1 _17791_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__18885__S _18885_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19268__S1 _20131_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19530_ _19784_/CLK _19530_/D vssd1 vssd1 vccd1 vccd1 _19530_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_235_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16742_ _16744_/A _16742_/B vssd1 vssd1 vccd1 vccd1 _19911_/D sky130_fd_sc_hd__nor2_1
XFILLER_143_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13954_ _20649_/Q vssd1 vssd1 vccd1 vccd1 _13954_/Y sky130_fd_sc_hd__inv_2
XFILLER_219_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12665__B1 _12663_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12905_ _20734_/Q _12901_/X _12651_/X _12904_/X vssd1 vssd1 vccd1 vccd1 _20734_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_246_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16673_ _21161_/Q _11449_/B _11450_/B vssd1 vssd1 vccd1 vccd1 _16673_/X sky130_fd_sc_hd__a21bo_1
X_19461_ _20136_/CLK _19461_/D vssd1 vssd1 vccd1 vccd1 _19461_/Q sky130_fd_sc_hd__dfxtp_1
X_13885_ _13972_/B _13885_/B vssd1 vssd1 vccd1 vccd1 _13996_/A sky130_fd_sc_hd__or2_1
XFILLER_35_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15603__A _15603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18412_ _18411_/X _13911_/Y _18849_/S vssd1 vssd1 vccd1 vccd1 _18412_/X sky130_fd_sc_hd__mux2_1
X_12836_ _12842_/A vssd1 vssd1 vccd1 vccd1 _12836_/X sky130_fd_sc_hd__buf_1
X_15624_ _15919_/A _15624_/B _16451_/C vssd1 vssd1 vccd1 vccd1 _15632_/A sky130_fd_sc_hd__or3_4
X_19392_ _21222_/CLK _19392_/D vssd1 vssd1 vccd1 vccd1 _19392_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18343_ _18342_/X _15148_/Y _18906_/S vssd1 vssd1 vccd1 vccd1 _18343_/X sky130_fd_sc_hd__mux2_1
X_15555_ _19745_/Q _15553_/X _15518_/X _15554_/X vssd1 vssd1 vccd1 vccd1 _19745_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_187_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12767_ _20800_/Q _12765_/X _12663_/X _12766_/X vssd1 vssd1 vccd1 vccd1 _20800_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13090__B1 _13030_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14506_ _14504_/A _14504_/B _14504_/Y _14488_/X vssd1 vssd1 vccd1 vccd1 _20219_/D
+ sky130_fd_sc_hd__a211oi_2
XPHY_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11718_ _21069_/Q _11713_/X _11686_/X _11715_/X vssd1 vssd1 vccd1 vccd1 _21069_/D
+ sky130_fd_sc_hd__a22o_1
X_18274_ _18273_/X _14910_/Y _18907_/S vssd1 vssd1 vccd1 vccd1 _18274_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15486_ _19775_/Q _15479_/X _15485_/X _15481_/X vssd1 vssd1 vccd1 vccd1 _19775_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_30_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12698_ _20820_/Q _12693_/X _12697_/X _12694_/X vssd1 vssd1 vccd1 vccd1 _20820_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_187_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14437_ _14414_/Y _20209_/Q _21477_/Q _14462_/B _14436_/X vssd1 vssd1 vccd1 vccd1
+ _14437_/X sky130_fd_sc_hd__a221o_1
X_17225_ _17320_/A vssd1 vssd1 vccd1 vccd1 _17226_/A sky130_fd_sc_hd__buf_1
XFILLER_238_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11649_ _18982_/X _11640_/A _21098_/Q _11646_/X vssd1 vssd1 vccd1 vccd1 _21098_/D
+ sky130_fd_sc_hd__a22o_1
Xinput11 HADDR[19] vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__clkbuf_1
Xinput22 HADDR[29] vssd1 vssd1 vccd1 vccd1 input22/X sky130_fd_sc_hd__buf_1
XANTENNA__18125__S _18902_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput33 HREADY vssd1 vssd1 vccd1 vccd1 input33/X sky130_fd_sc_hd__buf_1
X_17156_ _17145_/Y _17147_/X _17148_/Y _17150_/X _17155_/X vssd1 vssd1 vccd1 vccd1
+ _17156_/X sky130_fd_sc_hd__o221a_1
Xinput44 HWDATA[15] vssd1 vssd1 vccd1 vccd1 input44/X sky130_fd_sc_hd__buf_2
XFILLER_7_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14368_ _14461_/D _14368_/B vssd1 vssd1 vccd1 vccd1 _14486_/A sky130_fd_sc_hd__or2_1
Xinput55 HWDATA[25] vssd1 vssd1 vccd1 vccd1 input55/X sky130_fd_sc_hd__clkbuf_4
XFILLER_155_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput66 HWDATA[6] vssd1 vssd1 vccd1 vccd1 input66/X sky130_fd_sc_hd__clkbuf_4
Xinput77 sda_i_S4 vssd1 vssd1 vccd1 vccd1 input77/X sky130_fd_sc_hd__clkbuf_1
XFILLER_143_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16107_ _16247_/A _16107_/B _16261_/C vssd1 vssd1 vccd1 vccd1 _16119_/A sky130_fd_sc_hd__or3_4
X_13319_ _20535_/Q _13315_/X _13245_/X _13316_/X vssd1 vssd1 vccd1 vccd1 _20535_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_182_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17087_ _17087_/A vssd1 vssd1 vccd1 vccd1 _18899_/S sky130_fd_sc_hd__clkinv_8
X_14299_ _15490_/A vssd1 vssd1 vccd1 vccd1 _14315_/A sky130_fd_sc_hd__buf_1
XANTENNA__18608__A0 _17079_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16038_ _19517_/Q _16035_/X _15969_/X _16037_/X vssd1 vssd1 vccd1 vccd1 _19517_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_88_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19259__S1 _20131_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18795__S _18930_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17989_ _17989_/A _17989_/B _17989_/C _17989_/D vssd1 vssd1 vccd1 vccd1 _17989_/X
+ sky130_fd_sc_hd__or4_4
XFILLER_85_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_245_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19728_ _19784_/CLK _19728_/D vssd1 vssd1 vccd1 vccd1 _19728_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19659_ _19821_/CLK _19659_/D vssd1 vssd1 vccd1 vccd1 _19659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10131__A1 _10154_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15513__A input64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11150__A1_N _21004_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_241_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10419__C1 _10381_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_221_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20503_ _21375_/CLK _20503_/D repeater267/X vssd1 vssd1 vccd1 vccd1 _20503_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_138_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21483_ _21483_/CLK _21483_/D repeater200/X vssd1 vssd1 vccd1 vccd1 _21483_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__12872__A _13163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21053__RESET_B repeater225/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19195__S0 _19280_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20434_ _20937_/CLK _20434_/D repeater278/X vssd1 vssd1 vccd1 vccd1 _20434_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_174_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11488__A _20872_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20365_ _20951_/CLK _20365_/D repeater271/X vssd1 vssd1 vccd1 vccd1 _20365_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_106_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20296_ _20322_/CLK _20296_/D repeater262/X vssd1 vssd1 vccd1 vccd1 _20296_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17175__A _17177_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10370__A1 _21373_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10951_ _21203_/Q vssd1 vssd1 vccd1 vccd1 _10951_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17586__B1 _17572_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_243_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13670_ _20358_/Q _13667_/X _13553_/X _13668_/X vssd1 vssd1 vccd1 vccd1 _20358_/D
+ sky130_fd_sc_hd__a22o_1
X_10882_ _21259_/Q _10879_/X _09663_/X _10881_/X vssd1 vssd1 vccd1 vccd1 _21259_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_243_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12621_ input8/X _12619_/X _20859_/Q _12620_/X vssd1 vssd1 vccd1 vccd1 _20859_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_73_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15340_ _19837_/Q _15337_/X _14258_/X _15339_/X vssd1 vssd1 vccd1 vccd1 _19837_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12552_ _20897_/Q _12543_/X _11733_/X _12546_/X vssd1 vssd1 vccd1 vccd1 _20897_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11503_ _11502_/X _11487_/X _19111_/S _11500_/Y _21150_/Q vssd1 vssd1 vccd1 vccd1
+ _21150_/D sky130_fd_sc_hd__a32o_1
XPHY_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15271_ _20482_/Q vssd1 vssd1 vccd1 vccd1 _17938_/A sky130_fd_sc_hd__inv_2
XFILLER_129_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12483_ _12483_/A vssd1 vssd1 vccd1 vccd1 _12483_/Y sky130_fd_sc_hd__inv_2
XPHY_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17010_ _17008_/Y _17009_/X _16984_/X vssd1 vssd1 vccd1 vccd1 _17010_/X sky130_fd_sc_hd__o21a_1
XFILLER_184_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19186__S0 _20123_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14222_ _14222_/A vssd1 vssd1 vccd1 vccd1 _14222_/Y sky130_fd_sc_hd__inv_2
X_11434_ _11388_/A _11420_/X _11389_/C _11421_/X vssd1 vssd1 vccd1 vccd1 _21171_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_172_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14153_ _20552_/Q _14091_/A _18003_/A _20281_/Q vssd1 vssd1 vccd1 vccd1 _14153_/X
+ sky130_fd_sc_hd__o22a_1
X_11365_ _11365_/A _11364_/X vssd1 vssd1 vccd1 vccd1 _11410_/A sky130_fd_sc_hd__or2b_1
XFILLER_164_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13104_ _13108_/A _13104_/B vssd1 vssd1 vccd1 vccd1 _13105_/S sky130_fd_sc_hd__or2_1
XFILLER_125_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10316_ _20703_/Q vssd1 vssd1 vccd1 vccd1 _10316_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18961_ _16635_/X _21075_/Q _18962_/S vssd1 vssd1 vccd1 vccd1 _18961_/X sky130_fd_sc_hd__mux2_1
X_14084_ _14084_/A _14204_/A vssd1 vssd1 vccd1 vccd1 _14085_/B sky130_fd_sc_hd__or2_2
X_11296_ _20903_/Q vssd1 vssd1 vccd1 vccd1 _11306_/B sky130_fd_sc_hd__buf_1
XANTENNA__12006__B _19888_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13035_ _13041_/A vssd1 vssd1 vccd1 vccd1 _13035_/X sky130_fd_sc_hd__buf_1
X_17912_ _20826_/Q vssd1 vssd1 vccd1 vccd1 _17912_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10247_ _21356_/Q vssd1 vssd1 vccd1 vccd1 _10271_/A sky130_fd_sc_hd__inv_2
XANTENNA__20705__RESET_B repeater210/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18892_ _18891_/X _10754_/A _18898_/S vssd1 vssd1 vccd1 vccd1 _18892_/X sky130_fd_sc_hd__mux2_2
XANTENNA_repeater206_A repeater207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17843_ _18602_/X _17839_/X _18606_/X _17840_/X _17842_/X vssd1 vssd1 vccd1 vccd1
+ _17843_/X sky130_fd_sc_hd__o221a_4
X_10178_ _10161_/A _10161_/B _10177_/X _10175_/Y vssd1 vssd1 vccd1 vccd1 _21400_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_227_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17774_ _18675_/X _17774_/B vssd1 vssd1 vccd1 vccd1 _17774_/X sky130_fd_sc_hd__and2_1
XFILLER_93_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14986_ _14961_/A _14872_/B _14984_/Y _14975_/X vssd1 vssd1 vccd1 vccd1 _20094_/D
+ sky130_fd_sc_hd__a211oi_2
X_19513_ _21462_/CLK _19513_/D vssd1 vssd1 vccd1 vccd1 _19513_/Q sky130_fd_sc_hd__dfxtp_1
X_16725_ _20987_/Q _11993_/B _11994_/B vssd1 vssd1 vccd1 vccd1 _16725_/X sky130_fd_sc_hd__a21bo_1
XFILLER_235_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13937_ _20644_/Q _13875_/A _20656_/Q _13974_/B vssd1 vssd1 vccd1 vccd1 _13937_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_34_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12957__A _14264_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_235_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19444_ _19834_/CLK _19444_/D vssd1 vssd1 vccd1 vccd1 _19444_/Q sky130_fd_sc_hd__dfxtp_1
X_16656_ _19862_/Q _15296_/B _15297_/B vssd1 vssd1 vccd1 vccd1 _16656_/X sky130_fd_sc_hd__a21bo_1
X_13868_ _20296_/Q vssd1 vssd1 vccd1 vccd1 _14012_/A sky130_fd_sc_hd__inv_2
XFILLER_223_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15607_ _19719_/Q _15603_/X _15485_/X _15604_/X vssd1 vssd1 vccd1 vccd1 _19719_/D
+ sky130_fd_sc_hd__a22o_1
X_12819_ _17083_/A _12973_/A vssd1 vssd1 vccd1 vccd1 _12847_/A sky130_fd_sc_hd__or2_2
X_19375_ _19706_/CLK _19375_/D vssd1 vssd1 vccd1 vccd1 _19375_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13063__B1 _12999_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16587_ _16587_/A _16587_/B vssd1 vssd1 vccd1 vccd1 _16588_/A sky130_fd_sc_hd__or2_1
X_13799_ _20202_/Q vssd1 vssd1 vccd1 vccd1 _14591_/A sky130_fd_sc_hd__inv_2
XFILLER_231_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18326_ _18325_/X _14937_/Y _18907_/S vssd1 vssd1 vccd1 vccd1 _18326_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15538_ _19753_/Q _15536_/X _15518_/X _15537_/X vssd1 vssd1 vccd1 vccd1 _19753_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_30_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19959__RESET_B repeater184/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13788__A _20193_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18257_ _18256_/X _14446_/Y _18897_/S vssd1 vssd1 vccd1 vccd1 _18257_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15469_ _15758_/A vssd1 vssd1 vccd1 vccd1 _15469_/X sky130_fd_sc_hd__buf_1
XFILLER_175_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19177__S0 _19280_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14563__B1 _20133_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17208_ _18880_/X _17200_/X _18886_/X _17203_/X _17207_/X vssd1 vssd1 vccd1 vccd1
+ _17235_/B sky130_fd_sc_hd__o221a_1
XFILLER_128_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18188_ _18187_/X _10771_/A _18617_/S vssd1 vssd1 vccd1 vccd1 _18188_/X sky130_fd_sc_hd__mux2_1
XFILLER_116_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17139_ _17139_/A vssd1 vssd1 vccd1 vccd1 _17177_/B sky130_fd_sc_hd__buf_2
X_20150_ _21239_/CLK _20150_/D repeater250/X vssd1 vssd1 vccd1 vccd1 _20150_/Q sky130_fd_sc_hd__dfrtp_4
X_09961_ _21423_/Q _09957_/X _09698_/X _09958_/X vssd1 vssd1 vccd1 vccd1 _21423_/D
+ sky130_fd_sc_hd__a22o_1
X_20081_ _20590_/CLK _20081_/D repeater260/X vssd1 vssd1 vccd1 vccd1 _20081_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12877__B1 _12875_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09892_ _09890_/Y _17025_/A _09890_/Y _17025_/A vssd1 vssd1 vccd1 vccd1 _09916_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_69_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20983_ _21141_/CLK _20983_/D repeater191/X vssd1 vssd1 vccd1 vccd1 _20983_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_66_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__21234__RESET_B repeater270/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12801__B1 _12550_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19168__S0 _19280_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21466_ _21477_/CLK _21466_/D repeater204/X vssd1 vssd1 vccd1 vccd1 _21466_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_153_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20417_ _20957_/CLK _20417_/D repeater187/X vssd1 vssd1 vccd1 vccd1 _20417_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_175_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21397_ _21401_/CLK _21397_/D repeater253/X vssd1 vssd1 vccd1 vccd1 _21397_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__09981__B1 _09698_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11150_ _21004_/Q _11149_/Y _21004_/Q _11149_/Y vssd1 vssd1 vccd1 vccd1 _11926_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_20348_ _20476_/CLK _20348_/D repeater183/X vssd1 vssd1 vccd1 vccd1 _20348_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_122_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10101_ _21378_/Q _20775_/Q _10041_/B _10100_/Y vssd1 vssd1 vccd1 vccd1 _10101_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_1_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11081_ _21235_/Q _11081_/B vssd1 vssd1 vccd1 vccd1 _11081_/Y sky130_fd_sc_hd__nor2_1
XFILLER_88_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20279_ _20293_/CLK _20279_/D repeater263/X vssd1 vssd1 vccd1 vccd1 _20279_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_88_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10032_ _21404_/Q vssd1 vssd1 vccd1 vccd1 _10034_/A sky130_fd_sc_hd__inv_2
XFILLER_88_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14840_ _20094_/Q vssd1 vssd1 vccd1 vccd1 _14961_/A sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_60_HCLK clkbuf_4_14_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _21481_/CLK sky130_fd_sc_hd__clkbuf_16
X_14771_ _16451_/A vssd1 vssd1 vccd1 vccd1 _15448_/A sky130_fd_sc_hd__buf_1
XANTENNA_input17_A HADDR[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_217_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11983_ _11983_/A _11983_/B _11983_/C _19118_/X vssd1 vssd1 vccd1 vccd1 _11983_/X
+ sky130_fd_sc_hd__or4b_4
XFILLER_232_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16510_ _16510_/A vssd1 vssd1 vccd1 vccd1 _16510_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13722_ _20329_/Q vssd1 vssd1 vccd1 vccd1 _15764_/A sky130_fd_sc_hd__buf_1
X_10934_ _21024_/Q vssd1 vssd1 vccd1 vccd1 _10934_/X sky130_fd_sc_hd__buf_1
XFILLER_205_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17490_ _19394_/Q vssd1 vssd1 vccd1 vccd1 _17490_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13653_ _20367_/Q _13651_/X _13446_/X _13652_/X vssd1 vssd1 vccd1 vccd1 _20367_/D
+ sky130_fd_sc_hd__a22o_1
X_16441_ _16441_/A vssd1 vssd1 vccd1 vccd1 _16441_/X sky130_fd_sc_hd__buf_1
XANTENNA__13045__B1 _12884_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10865_ _10871_/A vssd1 vssd1 vccd1 vccd1 _10872_/A sky130_fd_sc_hd__inv_2
XFILLER_32_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_220_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12604_ _17060_/A _12600_/X _18222_/X _12601_/X vssd1 vssd1 vccd1 vccd1 _20870_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16372_ _19352_/Q _16370_/X _16207_/X _16371_/X vssd1 vssd1 vccd1 vccd1 _19352_/D
+ sky130_fd_sc_hd__a22o_1
X_19160_ _19660_/Q _19652_/Q _19636_/Q _19820_/Q _19285_/S0 _21017_/Q vssd1 vssd1
+ vccd1 vccd1 _19160_/X sky130_fd_sc_hd__mux4_2
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13584_ input69/X vssd1 vssd1 vccd1 vccd1 _13584_/X sky130_fd_sc_hd__clkbuf_4
X_10796_ _10779_/A _10779_/B _10795_/X _10793_/Y vssd1 vssd1 vccd1 vccd1 _21303_/D
+ sky130_fd_sc_hd__a211oi_2
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18111_ _17531_/Y _17630_/Y _17444_/Y _17530_/X _18110_/X vssd1 vssd1 vccd1 vccd1
+ _18112_/B sky130_fd_sc_hd__o221a_2
X_15323_ _15329_/A vssd1 vssd1 vccd1 vccd1 _15323_/X sky130_fd_sc_hd__buf_1
X_12535_ _11310_/C _12518_/A _12500_/A _12521_/X vssd1 vssd1 vccd1 vccd1 _20907_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19091_ _16679_/X _21087_/Q _19870_/D vssd1 vssd1 vccd1 vccd1 _19091_/X sky130_fd_sc_hd__mux2_1
XFILLER_185_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_repeater156_A _18667_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19159__S0 _19285_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15254_ _20492_/Q _20071_/Q _15253_/Y _15085_/A vssd1 vssd1 vccd1 vccd1 _15259_/B
+ sky130_fd_sc_hd__o22a_1
X_18042_ _18042_/A _18042_/B _18042_/C _18042_/D vssd1 vssd1 vccd1 vccd1 _18042_/X
+ sky130_fd_sc_hd__or4_4
XFILLER_129_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12466_ _20931_/Q _12465_/Y _12480_/A _12421_/B vssd1 vssd1 vccd1 vccd1 _20931_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_173_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20957__RESET_B repeater187/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14205_ _14205_/A vssd1 vssd1 vccd1 vccd1 _14205_/X sky130_fd_sc_hd__clkbuf_2
X_11417_ _21180_/Q vssd1 vssd1 vccd1 vccd1 _11783_/B sky130_fd_sc_hd__inv_2
X_15185_ _15185_/A vssd1 vssd1 vccd1 vccd1 _15185_/X sky130_fd_sc_hd__buf_1
X_12397_ _12473_/A _12472_/A _12471_/A _12468_/A vssd1 vssd1 vccd1 vccd1 _12399_/C
+ sky130_fd_sc_hd__or4_4
XANTENNA__18403__S _18910_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16712__A _16718_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output85_A _17919_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12571__A2 _12566_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14136_ _14134_/Y _20269_/Q _17977_/A _20279_/Q vssd1 vssd1 vccd1 vccd1 _14136_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09972__B1 _09666_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11348_ _21177_/Q _21176_/Q _11348_/C vssd1 vssd1 vccd1 vccd1 _11362_/B sky130_fd_sc_hd__or3_1
X_19993_ _21055_/CLK _19993_/D repeater221/X vssd1 vssd1 vccd1 vccd1 _19993_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_235_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10582__B2 _20764_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18039__A1 _18365_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18944_ _16695_/X _20897_/Q _18946_/S vssd1 vssd1 vccd1 vccd1 _18944_/X sky130_fd_sc_hd__mux2_1
XFILLER_141_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14067_ _20261_/Q vssd1 vssd1 vccd1 vccd1 _14072_/A sky130_fd_sc_hd__inv_2
X_11279_ _20906_/Q vssd1 vssd1 vccd1 vccd1 _11299_/A sky130_fd_sc_hd__buf_1
X_13018_ _13018_/A vssd1 vssd1 vccd1 vccd1 _13040_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_140_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21128__CLK _21134_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18875_ _18874_/X _16889_/B _18875_/S vssd1 vssd1 vccd1 vccd1 _18875_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11531__B1 _10886_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_239_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17826_ _18288_/X _17933_/A _18289_/X _17932_/A _17825_/Y vssd1 vssd1 vccd1 vccd1
+ _17827_/C sky130_fd_sc_hd__o221a_1
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17757_ _19485_/Q vssd1 vssd1 vccd1 vccd1 _17757_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14969_ _20103_/Q _14968_/Y _14881_/B _14968_/A _14958_/X vssd1 vssd1 vccd1 vccd1
+ _20103_/D sky130_fd_sc_hd__o221a_1
XFILLER_75_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16708_ _19898_/Q _14238_/B _14239_/B vssd1 vssd1 vccd1 vccd1 _16708_/X sky130_fd_sc_hd__a21bo_1
XFILLER_207_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17688_ _19323_/Q vssd1 vssd1 vccd1 vccd1 _17688_/Y sky130_fd_sc_hd__inv_2
X_19427_ _20331_/CLK _19427_/D vssd1 vssd1 vccd1 vccd1 _19427_/Q sky130_fd_sc_hd__dfxtp_1
X_16639_ _16643_/A _18960_/X vssd1 vssd1 vccd1 vccd1 _19854_/D sky130_fd_sc_hd__and2_1
XANTENNA__13036__B1 _12950_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19358_ _19521_/CLK _19358_/D vssd1 vssd1 vccd1 vccd1 _19358_/Q sky130_fd_sc_hd__dfxtp_1
X_18309_ _18845_/A0 _13744_/Y _18896_/S vssd1 vssd1 vccd1 vccd1 _18309_/X sky130_fd_sc_hd__mux2_1
XFILLER_175_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19289_ _21374_/CLK _20771_/Q vssd1 vssd1 vccd1 vccd1 _19289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21320_ _21321_/CLK _21320_/D repeater205/X vssd1 vssd1 vccd1 vccd1 _21320_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_190_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20698__RESET_B repeater205/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21251_ _21390_/CLK _21251_/D repeater239/X vssd1 vssd1 vccd1 vccd1 _21251_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_128_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20627__RESET_B repeater193/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18313__S _18897_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20202_ _20623_/CLK _20202_/D repeater194/X vssd1 vssd1 vccd1 vccd1 _20202_/Q sky130_fd_sc_hd__dfrtp_1
X_21182_ _21182_/CLK _21182_/D repeater216/X vssd1 vssd1 vccd1 vccd1 _21182_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_145_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20133_ _20136_/CLK _20133_/D repeater249/X vssd1 vssd1 vccd1 vccd1 _20133_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__20280__RESET_B repeater262/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09944_ _09931_/X _21430_/Q _09944_/S vssd1 vssd1 vccd1 vccd1 _21430_/D sky130_fd_sc_hd__mux2_1
XFILLER_89_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20064_ _20066_/CLK _20064_/D hold8/X vssd1 vssd1 vccd1 vccd1 _20064_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_38_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09875_ _09875_/A vssd1 vssd1 vccd1 vccd1 _21442_/D sky130_fd_sc_hd__inv_2
XANTENNA_input9_A HADDR[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_83_HCLK clkbuf_4_13_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _21486_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_246_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18450__A1 _10126_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrepeater250 repeater251/X vssd1 vssd1 vccd1 vccd1 repeater250/X sky130_fd_sc_hd__buf_8
XFILLER_234_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater261 repeater262/X vssd1 vssd1 vccd1 vccd1 repeater261/X sky130_fd_sc_hd__buf_6
XPHY_4404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater272 repeater278/X vssd1 vssd1 vccd1 vccd1 repeater272/X sky130_fd_sc_hd__buf_6
XANTENNA__13275__B1 _13274_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10628__A2 _20763_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_242_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20966_ _20981_/CLK _20966_/D repeater186/X vssd1 vssd1 vccd1 vccd1 _20966_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_4459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17900__B _17938_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20897_ _21147_/CLK _20897_/D repeater212/X vssd1 vssd1 vccd1 vccd1 _20897_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_198_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10650_ _10722_/A _10650_/B vssd1 vssd1 vccd1 vccd1 _10651_/B sky130_fd_sc_hd__or2_2
XFILLER_139_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10581_ _10723_/C _20739_/Q _10662_/A _20761_/Q vssd1 vssd1 vccd1 vccd1 _10581_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_10_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12320_ _12320_/A _12362_/A vssd1 vssd1 vccd1 vccd1 _12321_/B sky130_fd_sc_hd__or2_2
XANTENNA__13221__A input46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12251_ _20529_/Q vssd1 vssd1 vccd1 vccd1 _12251_/Y sky130_fd_sc_hd__inv_2
X_21449_ _21449_/CLK _21449_/D repeater248/X vssd1 vssd1 vccd1 vccd1 _21449_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_182_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18223__S _18236_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11202_ _15847_/A _17553_/A vssd1 vssd1 vccd1 vccd1 _16488_/A sky130_fd_sc_hd__or2_4
XANTENNA__09954__B1 _09676_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17477__C1 _17476_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12182_ _20963_/Q _12179_/Y _12316_/A _20345_/Q _12181_/X vssd1 vssd1 vccd1 vccd1
+ _12190_/B sky130_fd_sc_hd__o221a_1
XFILLER_123_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11133_ _11124_/Y _11132_/X _11124_/Y _11132_/X vssd1 vssd1 vccd1 vccd1 _11151_/A
+ sky130_fd_sc_hd__a2bb2o_1
Xclkbuf_3_2_0_HCLK clkbuf_3_3_0_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_5_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_79_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16990_ _16994_/B _16989_/X _16967_/X vssd1 vssd1 vccd1 vccd1 _16990_/X sky130_fd_sc_hd__o21a_1
XFILLER_150_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15941_ _16332_/A vssd1 vssd1 vccd1 vccd1 _15941_/X sky130_fd_sc_hd__clkbuf_2
X_11064_ _20138_/Q vssd1 vssd1 vccd1 vccd1 _11101_/A sky130_fd_sc_hd__buf_1
XFILLER_95_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19054__S _19058_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10015_ _21417_/Q _17034_/A _10006_/X _10011_/X _10014_/X vssd1 vssd1 vccd1 vccd1
+ _10015_/X sky130_fd_sc_hd__o2111a_1
XFILLER_236_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18660_ _18659_/X _17003_/Y _18875_/S vssd1 vssd1 vccd1 vccd1 _18660_/X sky130_fd_sc_hd__mux2_1
X_15872_ _19595_/Q _15864_/X _15871_/X _15867_/X vssd1 vssd1 vccd1 vccd1 _19595_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_218_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17611_ _19483_/Q vssd1 vssd1 vccd1 vccd1 _17611_/Y sky130_fd_sc_hd__inv_2
X_14823_ _20024_/Q _20109_/Q _14823_/S vssd1 vssd1 vccd1 vccd1 _20109_/D sky130_fd_sc_hd__mux2_1
X_18591_ _18845_/A0 _10423_/Y _18896_/S vssd1 vssd1 vccd1 vccd1 _18591_/X sky130_fd_sc_hd__mux2_1
XFILLER_63_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18893__S _18899_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output123_A _17078_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17542_ _17542_/A _17542_/B vssd1 vssd1 vccd1 vccd1 _17542_/Y sky130_fd_sc_hd__nor2_1
XFILLER_151_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14754_ _14754_/A vssd1 vssd1 vccd1 vccd1 _14754_/Y sky130_fd_sc_hd__inv_2
X_11966_ _21002_/Q _11961_/Y _13717_/C vssd1 vssd1 vccd1 vccd1 _11966_/X sky130_fd_sc_hd__a21o_1
XFILLER_232_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13705_ _20336_/Q _13699_/X _13704_/X _13700_/X vssd1 vssd1 vccd1 vccd1 _20336_/D
+ sky130_fd_sc_hd__a22o_1
X_10917_ _10917_/A _14680_/A _14679_/A vssd1 vssd1 vccd1 vccd1 _10918_/B sky130_fd_sc_hd__or3_4
XANTENNA__17810__B _17812_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14685_ _14685_/A vssd1 vssd1 vccd1 vccd1 _16490_/B sky130_fd_sc_hd__buf_1
X_17473_ _18789_/X vssd1 vssd1 vccd1 vccd1 _17473_/Y sky130_fd_sc_hd__inv_2
X_11897_ _11897_/A vssd1 vssd1 vccd1 vccd1 _11900_/A sky130_fd_sc_hd__inv_2
X_19212_ _17666_/Y _17667_/Y _17668_/Y _17669_/Y _19275_/S0 _21004_/Q vssd1 vssd1
+ vccd1 vccd1 _19212_/X sky130_fd_sc_hd__mux4_2
XFILLER_220_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16424_ _19323_/Q _16420_/X _15869_/A _16422_/X vssd1 vssd1 vccd1 vccd1 _19323_/D
+ sky130_fd_sc_hd__a22o_1
X_13636_ _20378_/Q _13632_/X _13422_/X _13634_/X vssd1 vssd1 vccd1 vccd1 _20378_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_60_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10848_ _19281_/X _15314_/A _10846_/X _21276_/Q _10847_/X vssd1 vssd1 vccd1 vccd1
+ _21276_/D sky130_fd_sc_hd__a32o_1
XFILLER_220_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19143_ _19761_/Q _19753_/Q _19745_/Q _19737_/Q _19285_/S0 _21017_/Q vssd1 vssd1
+ vccd1 vccd1 _19143_/X sky130_fd_sc_hd__mux4_2
XFILLER_158_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13567_ _13567_/A vssd1 vssd1 vccd1 vccd1 _13567_/X sky130_fd_sc_hd__buf_1
X_16355_ _19360_/Q _16352_/X _16291_/X _16353_/X vssd1 vssd1 vccd1 vccd1 _19360_/D
+ sky130_fd_sc_hd__a22o_1
X_10779_ _10779_/A _10779_/B vssd1 vssd1 vccd1 vccd1 _10793_/A sky130_fd_sc_hd__or2_1
XANTENNA__09788__A3 input74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15306_ _20040_/Q _15302_/X _19869_/Q _15305_/X vssd1 vssd1 vccd1 vccd1 _20040_/D
+ sky130_fd_sc_hd__a22o_1
X_12518_ _12518_/A vssd1 vssd1 vccd1 vccd1 _12518_/X sky130_fd_sc_hd__buf_1
XFILLER_145_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19074_ _16729_/X _21136_/Q _19908_/D vssd1 vssd1 vccd1 vccd1 _19074_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16286_ _19394_/Q _16276_/X _16285_/X _16279_/X vssd1 vssd1 vccd1 vccd1 _19394_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_172_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13498_ _20445_/Q _13492_/X _13426_/X _13494_/X vssd1 vssd1 vccd1 vccd1 _20445_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__20791__RESET_B repeater255/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18025_ _18350_/X _17963_/X _18318_/X _17996_/X vssd1 vssd1 vccd1 vccd1 _18025_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_246_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15237_ _20467_/Q vssd1 vssd1 vccd1 vccd1 _15237_/Y sky130_fd_sc_hd__inv_2
X_12449_ _20941_/Q _12447_/Y _12448_/X _12431_/B vssd1 vssd1 vccd1 vccd1 _20941_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__20720__RESET_B repeater264/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18133__S _18748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13741__B2 _20193_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15168_ _15086_/A _15086_/B _15165_/Y _15201_/B vssd1 vssd1 vccd1 vccd1 _20072_/D
+ sky130_fd_sc_hd__a211oi_4
XFILLER_99_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14119_ _14116_/Y _20266_/Q _20535_/Q _14075_/A _14118_/X vssd1 vssd1 vccd1 vccd1
+ _14120_/D sky130_fd_sc_hd__o221a_1
XFILLER_4_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17483__A2 _17461_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15099_ _15099_/A vssd1 vssd1 vccd1 vccd1 _15099_/X sky130_fd_sc_hd__buf_2
X_19976_ _20809_/CLK _19976_/D repeater188/X vssd1 vssd1 vccd1 vccd1 _19976_/Q sky130_fd_sc_hd__dfrtp_1
X_18927_ _18926_/X _18109_/A _18927_/S vssd1 vssd1 vccd1 vccd1 _18927_/X sky130_fd_sc_hd__mux2_1
XFILLER_228_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09660_ _09660_/A vssd1 vssd1 vccd1 vccd1 _09660_/X sky130_fd_sc_hd__buf_1
XANTENNA__18432__A1 _20447_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18858_ _18857_/X _21409_/Q _20869_/Q vssd1 vssd1 vccd1 vccd1 _18858_/X sky130_fd_sc_hd__mux2_1
XFILLER_216_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17809_ _17809_/A _17812_/B vssd1 vssd1 vccd1 vccd1 _17809_/Y sky130_fd_sc_hd__nor2_1
XFILLER_27_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18789_ _17449_/X _21415_/Q _20870_/Q vssd1 vssd1 vccd1 vccd1 _18789_/X sky130_fd_sc_hd__mux2_1
XFILLER_215_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20820_ _21374_/CLK _20820_/D repeater256/X vssd1 vssd1 vccd1 vccd1 _20820_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_224_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20751_ _21342_/CLK _20751_/D repeater210/X vssd1 vssd1 vccd1 vccd1 _20751_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13009__B1 _12918_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18308__S _18886_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15521__A _15588_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20682_ _21302_/CLK _20682_/D repeater208/X vssd1 vssd1 vccd1 vccd1 _20682_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13041__A _13041_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21303_ _21306_/CLK _21303_/D repeater207/X vssd1 vssd1 vccd1 vccd1 _21303_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_156_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21234_ _21234_/CLK _21234_/D repeater270/X vssd1 vssd1 vccd1 vccd1 _21234_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_172_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21165_ _21167_/CLK _21165_/D repeater225/X vssd1 vssd1 vccd1 vccd1 _21165_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_105_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20024__D input72/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20116_ _21419_/CLK _20116_/D repeater234/X vssd1 vssd1 vccd1 vccd1 _20116_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_104_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09927_ _21432_/Q _21433_/Q _09929_/S vssd1 vssd1 vccd1 vccd1 _21433_/D sky130_fd_sc_hd__mux2_1
X_21096_ _21120_/CLK _21096_/D repeater231/X vssd1 vssd1 vccd1 vccd1 _21096_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__13496__B1 _13422_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20047_ _20066_/CLK _20047_/D repeater281/X vssd1 vssd1 vccd1 vccd1 _20047_/Q sky130_fd_sc_hd__dfrtp_4
X_09858_ _09853_/X _09857_/A _21445_/Q _09840_/X _09849_/X vssd1 vssd1 vccd1 vccd1
+ _09859_/B sky130_fd_sc_hd__a41o_1
XFILLER_246_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09789_ _16619_/A _09787_/X _09788_/X vssd1 vssd1 vccd1 vccd1 _09789_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_45_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13216__A input48/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11820_ _11820_/A vssd1 vssd1 vccd1 vccd1 _21039_/D sky130_fd_sc_hd__inv_2
XPHY_4234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11751_ _21052_/Q vssd1 vssd1 vccd1 vccd1 _11761_/A sky130_fd_sc_hd__buf_1
XPHY_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20949_ _20949_/CLK _20949_/D repeater272/X vssd1 vssd1 vccd1 vccd1 _20949_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_4289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10702_ _10702_/A _10720_/A vssd1 vssd1 vccd1 vccd1 _10718_/A sky130_fd_sc_hd__or2_2
XANTENNA__15431__A _15592_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14470_ _14378_/A _14378_/B _14469_/X _14380_/C vssd1 vssd1 vccd1 vccd1 _20235_/D
+ sky130_fd_sc_hd__a211oi_2
XPHY_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11682_ _11690_/A vssd1 vssd1 vccd1 vccd1 _11682_/X sky130_fd_sc_hd__buf_1
XPHY_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13421_ _20480_/Q _13417_/X _13418_/X _13420_/X vssd1 vssd1 vccd1 vccd1 _20480_/D
+ sky130_fd_sc_hd__a22o_1
X_10633_ _21312_/Q _10629_/Y _21339_/Q _10630_/Y _10632_/X vssd1 vssd1 vccd1 vccd1
+ _10638_/C sky130_fd_sc_hd__o221a_1
XPHY_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16140_ _19466_/Q _16130_/X _16139_/X _16133_/X vssd1 vssd1 vccd1 vccd1 _19466_/D
+ sky130_fd_sc_hd__a22o_1
X_13352_ _13352_/A vssd1 vssd1 vccd1 vccd1 _13352_/X sky130_fd_sc_hd__buf_1
X_10564_ _21326_/Q vssd1 vssd1 vccd1 vccd1 _10655_/A sky130_fd_sc_hd__inv_2
XFILLER_154_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12303_ _12453_/A vssd1 vssd1 vccd1 vccd1 _12410_/A sky130_fd_sc_hd__inv_2
XFILLER_182_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16071_ _16071_/A vssd1 vssd1 vccd1 vccd1 _16071_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__19049__S _19058_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13283_ _20555_/Q _13276_/X _13282_/X _13278_/X vssd1 vssd1 vccd1 vccd1 _20555_/D
+ sky130_fd_sc_hd__a22o_1
X_10495_ _21287_/Q _10490_/Y _10758_/A _20670_/Q _10494_/X vssd1 vssd1 vccd1 vccd1
+ _10496_/D sky130_fd_sc_hd__o221a_1
X_15022_ _15022_/A vssd1 vssd1 vccd1 vccd1 _15025_/A sky130_fd_sc_hd__inv_2
X_12234_ _20511_/Q vssd1 vssd1 vccd1 vccd1 _12234_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20131__RESET_B repeater249/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18888__S _18910_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11734__B1 _11733_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19830_ _19834_/CLK _19830_/D vssd1 vssd1 vccd1 vccd1 _19830_/Q sky130_fd_sc_hd__dfxtp_1
X_12165_ _20350_/Q vssd1 vssd1 vccd1 vccd1 _12165_/Y sky130_fd_sc_hd__inv_2
XFILLER_122_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11116_ _11116_/A vssd1 vssd1 vccd1 vccd1 _21227_/D sky130_fd_sc_hd__inv_2
XFILLER_110_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19761_ _21011_/CLK _19761_/D vssd1 vssd1 vccd1 vccd1 _19761_/Q sky130_fd_sc_hd__dfxtp_1
X_16973_ _16970_/A _16965_/A _16972_/Y vssd1 vssd1 vccd1 vccd1 _16974_/B sky130_fd_sc_hd__a21oi_1
X_12096_ _20958_/Q vssd1 vssd1 vccd1 vccd1 _12312_/A sky130_fd_sc_hd__inv_2
XFILLER_49_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18712_ _18711_/X _16770_/A _18880_/S vssd1 vssd1 vccd1 vccd1 _18712_/X sky130_fd_sc_hd__mux2_1
XANTENNA__21337__RESET_B repeater204/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15924_ _19572_/Q _15920_/X _15891_/X _15922_/X vssd1 vssd1 vccd1 vccd1 _19572_/D
+ sky130_fd_sc_hd__a22o_1
X_11047_ _21241_/Q _11021_/B _11022_/X vssd1 vssd1 vccd1 vccd1 _21241_/D sky130_fd_sc_hd__o21a_1
X_19692_ _19776_/CLK _19692_/D vssd1 vssd1 vccd1 vccd1 _19692_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput9 HADDR[17] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__clkbuf_1
XFILLER_77_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18643_ _18848_/A0 _10312_/Y _18884_/S vssd1 vssd1 vccd1 vccd1 _18643_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09604__A _14304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15855_ _19602_/Q _15849_/X _15785_/X _15851_/X vssd1 vssd1 vccd1 vccd1 _19602_/D
+ sky130_fd_sc_hd__a22o_1
X_14806_ _20120_/Q _14805_/X _20120_/Q _14805_/X vssd1 vssd1 vccd1 vccd1 _20120_/D
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_80_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18574_ _18848_/A0 _14134_/Y _18902_/S vssd1 vssd1 vccd1 vccd1 _18574_/X sky130_fd_sc_hd__mux2_1
XFILLER_206_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15786_ _19634_/Q _15779_/X _15785_/X _15781_/X vssd1 vssd1 vccd1 vccd1 _19634_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_224_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12998_ _20693_/Q _12995_/X _12996_/X _12997_/X vssd1 vssd1 vccd1 vccd1 _20693_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17525_ _20117_/Q _17131_/Y _14795_/Y _19334_/Q vssd1 vssd1 vccd1 vccd1 _17525_/X
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__17540__B _17542_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14737_ _20140_/Q _14731_/X _13712_/X _14733_/X vssd1 vssd1 vccd1 vccd1 _20140_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18128__S _18908_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11949_ _11943_/X _11947_/A _11943_/X _11947_/A vssd1 vssd1 vccd1 vccd1 _21007_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_60_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17456_ _21088_/Q vssd1 vssd1 vccd1 vccd1 _17456_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20972__RESET_B repeater187/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14668_ _14665_/X _14664_/X _14665_/X _14664_/X vssd1 vssd1 vccd1 vccd1 _20174_/D
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_60_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_103_HCLK_A clkbuf_4_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16407_ _16413_/A vssd1 vssd1 vccd1 vccd1 _16414_/A sky130_fd_sc_hd__inv_2
X_13619_ _13625_/A vssd1 vssd1 vccd1 vccd1 _13619_/X sky130_fd_sc_hd__buf_1
XANTENNA__20901__RESET_B repeater217/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17387_ _17387_/A vssd1 vssd1 vccd1 vccd1 _17387_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_leaf_166_HCLK_A clkbuf_opt_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14599_ _14624_/A vssd1 vssd1 vccd1 vccd1 _14599_/X sky130_fd_sc_hd__clkbuf_2
X_19126_ _16481_/Y _14275_/Y _19126_/S vssd1 vssd1 vccd1 vccd1 _19126_/X sky130_fd_sc_hd__mux2_2
XANTENNA__20219__RESET_B repeater202/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16338_ _16338_/A vssd1 vssd1 vccd1 vccd1 _16338_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_119_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13796__A _20611_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19057_ _16754_/Y _20812_/Q _19058_/S vssd1 vssd1 vccd1 vccd1 _19919_/D sky130_fd_sc_hd__mux2_1
X_16269_ _16269_/A vssd1 vssd1 vccd1 vccd1 _16269_/X sky130_fd_sc_hd__buf_1
XFILLER_173_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18008_ _18085_/B vssd1 vssd1 vccd1 vccd1 _18084_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_173_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18798__S _18928_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19959_ _20408_/CLK _19959_/D repeater184/X vssd1 vssd1 vccd1 vccd1 _19959_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_228_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09712_ _21455_/Q vssd1 vssd1 vccd1 vccd1 _09792_/A sky130_fd_sc_hd__inv_2
XFILLER_19_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17208__A2 _17200_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09643_ _09657_/A vssd1 vssd1 vccd1 vccd1 _09643_/X sky130_fd_sc_hd__buf_1
XANTENNA__21007__RESET_B repeater235/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18169__A0 _18848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_113_HCLK clkbuf_opt_3_HCLK/A vssd1 vssd1 vccd1 vccd1 _20480_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_224_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20803_ _21407_/CLK _20803_/D repeater213/X vssd1 vssd1 vccd1 vccd1 _20803_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13650__B1 _13442_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17916__B1 _18471_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12875__A _13166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20734_ _21366_/CLK _20734_/D repeater257/X vssd1 vssd1 vccd1 vccd1 _20734_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19706__CLK _19706_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13402__B1 _13282_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20665_ _20665_/CLK _20665_/D repeater261/X vssd1 vssd1 vccd1 vccd1 _20665_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_167_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_25_HCLK_A clkbuf_4_9_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20596_ _20665_/CLK _20596_/D repeater261/X vssd1 vssd1 vccd1 vccd1 _20596_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_192_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17178__A _17178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_88_HCLK_A clkbuf_4_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10280_ _10280_/A _10385_/A vssd1 vssd1 vccd1 vccd1 _10281_/B sky130_fd_sc_hd__or2_1
XFILLER_3_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21217_ _21223_/CLK _21217_/D repeater241/X vssd1 vssd1 vccd1 vccd1 _21217_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18644__A1 _10119_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18501__S _18910_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21148_ _21151_/CLK _21148_/D repeater223/X vssd1 vssd1 vccd1 vccd1 _21148_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_132_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13469__B1 _13280_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_219_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21079_ _21087_/CLK _21079_/D repeater227/X vssd1 vssd1 vccd1 vccd1 _21079_/Q sky130_fd_sc_hd__dfstp_1
X_13970_ _20320_/Q _13896_/B _13969_/X _13897_/B vssd1 vssd1 vccd1 vccd1 _20320_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_247_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12921_ _20724_/Q _12915_/X _12920_/X _12916_/X vssd1 vssd1 vccd1 vccd1 _20724_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_246_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17641__A _21085_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15640_ _15647_/A vssd1 vssd1 vccd1 vccd1 _15640_/X sky130_fd_sc_hd__buf_1
XPHY_4020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12852_ _20753_/Q _12848_/X _12849_/X _12851_/X vssd1 vssd1 vccd1 vccd1 _20753_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_132_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11803_ _11827_/A vssd1 vssd1 vccd1 vccd1 _11803_/X sky130_fd_sc_hd__buf_1
XFILLER_221_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15571_ _19736_/Q _15568_/X _15521_/X _15569_/X vssd1 vssd1 vccd1 vccd1 _19736_/D
+ sky130_fd_sc_hd__a22o_1
X_12783_ _12783_/A vssd1 vssd1 vccd1 vccd1 _12803_/A sky130_fd_sc_hd__clkbuf_2
XPHY_4075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13641__B1 _13429_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17310_ _18860_/X vssd1 vssd1 vccd1 vccd1 _17310_/Y sky130_fd_sc_hd__inv_2
XFILLER_203_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14522_ _14351_/B _14521_/A _20211_/Q _14524_/A _14458_/X vssd1 vssd1 vccd1 vccd1
+ _20211_/D sky130_fd_sc_hd__o221a_1
X_11734_ _21060_/Q _11727_/X _11733_/X _11729_/X vssd1 vssd1 vccd1 vccd1 _21060_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_242_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_214_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18290_ _17830_/X _10920_/Y _18928_/S vssd1 vssd1 vccd1 vccd1 _18290_/X sky130_fd_sc_hd__mux2_1
XPHY_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17241_ _19423_/Q vssd1 vssd1 vccd1 vccd1 _17241_/Y sky130_fd_sc_hd__inv_2
XPHY_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14453_ _14477_/A vssd1 vssd1 vccd1 vccd1 _14453_/X sky130_fd_sc_hd__clkbuf_2
X_11665_ _21091_/Q vssd1 vssd1 vccd1 vccd1 _11665_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15394__B1 _15355_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10616_ _10575_/A _10615_/Y _21340_/Q _20768_/Q vssd1 vssd1 vccd1 vccd1 _10616_/X
+ sky130_fd_sc_hd__a22o_1
X_13404_ _13410_/A vssd1 vssd1 vccd1 vccd1 _13404_/X sky130_fd_sc_hd__buf_1
XPHY_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14384_ _20240_/Q vssd1 vssd1 vccd1 vccd1 _14384_/Y sky130_fd_sc_hd__inv_2
X_17172_ _20498_/Q vssd1 vssd1 vccd1 vccd1 _17172_/Y sky130_fd_sc_hd__inv_2
XPHY_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18332__A0 _18848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11596_ _11596_/A _11596_/B vssd1 vssd1 vccd1 vccd1 _11599_/A sky130_fd_sc_hd__or2_1
XPHY_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13335_ _20529_/Q _13331_/X _13265_/X _13334_/X vssd1 vssd1 vccd1 vccd1 _20529_/D
+ sky130_fd_sc_hd__a22o_1
X_16123_ _20326_/Q vssd1 vssd1 vccd1 vccd1 _16123_/X sky130_fd_sc_hd__clkbuf_2
X_10547_ _21319_/Q vssd1 vssd1 vccd1 vccd1 _10707_/A sky130_fd_sc_hd__inv_2
XFILLER_182_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13266_ _13299_/A vssd1 vssd1 vccd1 vccd1 _13301_/A sky130_fd_sc_hd__inv_2
X_16054_ _19507_/Q _16049_/X _15764_/X _16051_/X vssd1 vssd1 vccd1 vccd1 _19507_/D
+ sky130_fd_sc_hd__a22o_1
X_10478_ _21282_/Q vssd1 vssd1 vccd1 vccd1 _10759_/A sky130_fd_sc_hd__inv_2
X_12217_ _20941_/Q vssd1 vssd1 vccd1 vccd1 _12430_/A sky130_fd_sc_hd__inv_2
X_15005_ _15005_/A _15009_/A vssd1 vssd1 vccd1 vccd1 _15006_/B sky130_fd_sc_hd__or2_2
XANTENNA__18096__C1 _18095_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18411__S _18902_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13197_ _20595_/Q _13192_/X _12989_/X _13195_/X vssd1 vssd1 vccd1 vccd1 _20595_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16720__A _16720_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19813_ _19813_/CLK _19813_/D vssd1 vssd1 vccd1 vccd1 _19813_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12148_ _12320_/A _20349_/Q _12093_/X _20344_/Q vssd1 vssd1 vccd1 vccd1 _12148_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_96_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17843__C1 _17842_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__21171__RESET_B repeater216/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19744_ _19765_/CLK _19744_/D vssd1 vssd1 vccd1 vccd1 _19744_/Q sky130_fd_sc_hd__dfxtp_1
X_12079_ _12073_/X _12074_/Y _12309_/A _20369_/Q _12078_/X vssd1 vssd1 vccd1 vccd1
+ _12087_/C sky130_fd_sc_hd__o221a_1
X_16956_ _16956_/A _16956_/B vssd1 vssd1 vccd1 vccd1 _16956_/Y sky130_fd_sc_hd__nor2_1
XFILLER_2_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18399__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_136_HCLK clkbuf_4_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20841_/CLK sky130_fd_sc_hd__clkbuf_16
X_15907_ _19581_/Q _15904_/X _15865_/X _15906_/X vssd1 vssd1 vccd1 vccd1 _19581_/D
+ sky130_fd_sc_hd__a22o_1
X_19675_ _19811_/CLK _19675_/D vssd1 vssd1 vccd1 vccd1 _19675_/Q sky130_fd_sc_hd__dfxtp_1
X_16887_ _19951_/Q vssd1 vssd1 vccd1 vccd1 _16889_/A sky130_fd_sc_hd__inv_2
XFILLER_238_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17551__A _21084_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18626_ _18083_/Y _20802_/Q _18885_/S vssd1 vssd1 vccd1 vccd1 _18626_/X sky130_fd_sc_hd__mux2_1
X_15838_ _19612_/Q _15834_/X _09821_/X _15836_/X vssd1 vssd1 vccd1 vccd1 _19612_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_65_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18557_ _17830_/X _10935_/Y _18928_/S vssd1 vssd1 vccd1 vccd1 _18557_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15769_ _15769_/A vssd1 vssd1 vccd1 vccd1 _15769_/X sky130_fd_sc_hd__buf_1
XFILLER_206_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17508_ _19602_/Q _17533_/B vssd1 vssd1 vccd1 vccd1 _17508_/Y sky130_fd_sc_hd__nand2_1
XFILLER_33_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_221_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18488_ _18487_/X _15116_/Y _18784_/S vssd1 vssd1 vccd1 vccd1 _18488_/X sky130_fd_sc_hd__mux2_2
XANTENNA__18571__A0 _18848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17439_ _19352_/Q vssd1 vssd1 vccd1 vccd1 _17439_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20450_ _20476_/CLK _20450_/D repeater280/X vssd1 vssd1 vccd1 vccd1 _20450_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__20053__RESET_B repeater281/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19109_ _16616_/Y _11123_/Y _19117_/S vssd1 vssd1 vccd1 vccd1 _19109_/X sky130_fd_sc_hd__mux2_2
XFILLER_118_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20381_ _20971_/CLK _20381_/D repeater183/X vssd1 vssd1 vccd1 vccd1 _20381_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_174_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput110 _17847_/Y vssd1 vssd1 vccd1 vccd1 HRDATA[9] sky130_fd_sc_hd__clkbuf_2
Xoutput121 _18114_/X vssd1 vssd1 vccd1 vccd1 IRQ[3] sky130_fd_sc_hd__clkbuf_2
XFILLER_133_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput132 _21248_/Q vssd1 vssd1 vccd1 vccd1 SCLK_S2 sky130_fd_sc_hd__clkbuf_2
XFILLER_217_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput143 _18124_/LO vssd1 vssd1 vccd1 vccd1 sda_o_S5 sky130_fd_sc_hd__clkbuf_2
XANTENNA__18321__S _18910_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21002_ _21125_/CLK _21002_/D repeater190/X vssd1 vssd1 vccd1 vccd1 _21002_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_130_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10382__C1 _10381_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_248_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09626_ input51/X vssd1 vssd1 vccd1 vccd1 _09626_/X sky130_fd_sc_hd__buf_4
XFILLER_43_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17180__B _17187_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20823__RESET_B repeater251/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20717_ _20724_/CLK _20717_/D repeater254/X vssd1 vssd1 vccd1 vccd1 _20717_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_23_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11450_ _21162_/Q _11450_/B vssd1 vssd1 vccd1 vccd1 _11451_/B sky130_fd_sc_hd__or2_1
XPHY_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20648_ _21486_/CLK _20648_/D repeater199/X vssd1 vssd1 vccd1 vccd1 _20648_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_17_HCLK clkbuf_4_3_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19821_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_127_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10401_ _10271_/A _10271_/B _10399_/Y _10397_/X vssd1 vssd1 vccd1 vccd1 _21356_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_137_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11381_ _21168_/Q vssd1 vssd1 vccd1 vccd1 _11384_/B sky130_fd_sc_hd__inv_2
XFILLER_109_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20579_ _20946_/CLK _20579_/D repeater274/X vssd1 vssd1 vccd1 vccd1 _20579_/Q sky130_fd_sc_hd__dfrtp_4
X_13120_ _13132_/A vssd1 vssd1 vccd1 vccd1 _13120_/X sky130_fd_sc_hd__buf_1
XFILLER_125_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10332_ _10265_/A _20708_/Q _21347_/Q _10329_/Y _10331_/X vssd1 vssd1 vccd1 vccd1
+ _10340_/B sky130_fd_sc_hd__o221a_1
XFILLER_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13051_ _13078_/A vssd1 vssd1 vccd1 vccd1 _13072_/A sky130_fd_sc_hd__clkbuf_2
X_10263_ _10263_/A _10415_/A vssd1 vssd1 vccd1 vccd1 _10264_/B sky130_fd_sc_hd__or2_2
XANTENNA__18231__S _18236_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12002_ _20996_/Q _12002_/B vssd1 vssd1 vccd1 vccd1 _12003_/B sky130_fd_sc_hd__or2_1
XFILLER_79_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_159_HCLK clkbuf_opt_1_HCLK/A vssd1 vssd1 vccd1 vccd1 _19835_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__18093__A2 _17205_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input47_A HWDATA[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10194_ _21391_/Q _10193_/Y _10183_/X _10153_/B vssd1 vssd1 vccd1 vccd1 _21391_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_239_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11684__A _12548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16810_ _19932_/Q _16801_/A _19933_/Q vssd1 vssd1 vccd1 vccd1 _16810_/X sky130_fd_sc_hd__o21a_1
X_17790_ _20900_/Q vssd1 vssd1 vccd1 vccd1 _17790_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16741_ _16535_/X _16537_/Y _16561_/Y _16583_/A _16539_/X vssd1 vssd1 vccd1 vccd1
+ _16742_/B sky130_fd_sc_hd__o32a_1
X_13953_ _20635_/Q _14031_/C _13951_/Y _20296_/Q _13952_/X vssd1 vssd1 vccd1 vccd1
+ _13961_/B sky130_fd_sc_hd__o221a_1
XFILLER_235_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19062__S _19910_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19460_ _20241_/CLK _19460_/D vssd1 vssd1 vccd1 vccd1 _19460_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12904_ _12926_/A vssd1 vssd1 vccd1 vccd1 _12904_/X sky130_fd_sc_hd__buf_1
XFILLER_235_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16672_ _21160_/Q _11448_/B _11449_/B vssd1 vssd1 vccd1 vccd1 _16672_/X sky130_fd_sc_hd__a21bo_1
XFILLER_34_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13884_ _13884_/A _13999_/A vssd1 vssd1 vccd1 vccd1 _13885_/B sky130_fd_sc_hd__or2_2
XFILLER_47_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18411_ _18848_/A0 _14164_/Y _18902_/S vssd1 vssd1 vccd1 vccd1 _18411_/X sky130_fd_sc_hd__mux2_1
X_15623_ _19710_/Q _15618_/X _15487_/X _15619_/X vssd1 vssd1 vccd1 vccd1 _19710_/D
+ sky130_fd_sc_hd__a22o_1
X_12835_ _12841_/A vssd1 vssd1 vccd1 vccd1 _12835_/X sky130_fd_sc_hd__buf_1
XFILLER_61_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19391_ _21222_/CLK _19391_/D vssd1 vssd1 vccd1 vccd1 _19391_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__20564__RESET_B repeater264/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater186_A repeater187/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18342_ _17079_/Y _15233_/Y _18908_/S vssd1 vssd1 vccd1 vccd1 _18342_/X sky130_fd_sc_hd__mux2_1
XFILLER_188_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09601__B _10859_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15554_ _15554_/A vssd1 vssd1 vccd1 vccd1 _15554_/X sky130_fd_sc_hd__buf_1
XPHY_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18553__A0 _17079_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12766_ _12778_/A vssd1 vssd1 vccd1 vccd1 _12766_/X sky130_fd_sc_hd__buf_1
XFILLER_203_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14505_ _20220_/Q _14504_/Y _14477_/A _14364_/B vssd1 vssd1 vccd1 vccd1 _20220_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_15_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11717_ _21070_/Q _11713_/X _11684_/X _11715_/X vssd1 vssd1 vccd1 vccd1 _21070_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18273_ _18272_/X _15102_/Y _18906_/S vssd1 vssd1 vccd1 vccd1 _18273_/X sky130_fd_sc_hd__mux2_1
XFILLER_187_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15485_ _15774_/A vssd1 vssd1 vccd1 vccd1 _15485_/X sky130_fd_sc_hd__buf_1
X_12697_ _13311_/A vssd1 vssd1 vccd1 vccd1 _12697_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_203_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18406__S _18908_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17224_ _17932_/A vssd1 vssd1 vccd1 vccd1 _17224_/X sky130_fd_sc_hd__buf_1
XPHY_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14436_ _21474_/Q _20220_/Q _14435_/Y _14361_/C vssd1 vssd1 vccd1 vccd1 _14436_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_187_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11648_ _18981_/X _11640_/A _21099_/Q _11646_/X vssd1 vssd1 vccd1 vccd1 _21099_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_128_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput12 HADDR[1] vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__buf_1
XFILLER_11_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput23 HADDR[2] vssd1 vssd1 vccd1 vccd1 input23/X sky130_fd_sc_hd__buf_1
XPHY_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput34 HRESETn vssd1 vssd1 vccd1 vccd1 hold8/A sky130_fd_sc_hd__clkbuf_2
XPHY_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17155_ _17046_/A _17151_/X _17152_/Y _17154_/X vssd1 vssd1 vccd1 vccd1 _17155_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_155_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput45 HWDATA[16] vssd1 vssd1 vccd1 vccd1 input45/X sky130_fd_sc_hd__clkbuf_4
X_11579_ _16541_/A vssd1 vssd1 vccd1 vccd1 _16545_/A sky130_fd_sc_hd__inv_2
X_14367_ _14462_/A _14490_/A vssd1 vssd1 vccd1 vccd1 _14368_/B sky130_fd_sc_hd__or2_1
XFILLER_156_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput56 HWDATA[26] vssd1 vssd1 vccd1 vccd1 input56/X sky130_fd_sc_hd__clkbuf_4
XFILLER_128_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput67 HWDATA[7] vssd1 vssd1 vccd1 vccd1 input67/X sky130_fd_sc_hd__clkbuf_4
Xinput78 sda_i_S5 vssd1 vssd1 vccd1 vccd1 input78/X sky130_fd_sc_hd__clkbuf_1
X_16106_ _19478_/Q _16101_/X _15916_/X _16102_/X vssd1 vssd1 vccd1 vccd1 _19478_/D
+ sky130_fd_sc_hd__a22o_1
X_13318_ _20536_/Q _13315_/X _13243_/X _13316_/X vssd1 vssd1 vccd1 vccd1 _20536_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_128_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_71_HCLK_A clkbuf_opt_6_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14298_ _15335_/A _15357_/B vssd1 vssd1 vccd1 vccd1 _15490_/A sky130_fd_sc_hd__or2_1
X_17086_ _20564_/Q _20108_/Q vssd1 vssd1 vccd1 vccd1 _17086_/X sky130_fd_sc_hd__and2_1
XFILLER_115_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19401__CLK _19813_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16037_ _16043_/A vssd1 vssd1 vccd1 vccd1 _16037_/X sky130_fd_sc_hd__buf_1
XANTENNA__21352__RESET_B repeater252/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18141__S _18748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13249_ _13249_/A vssd1 vssd1 vccd1 vccd1 _13249_/X sky130_fd_sc_hd__buf_1
XFILLER_130_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17988_ _18294_/X _17954_/X _18376_/X _17955_/X vssd1 vssd1 vccd1 vccd1 _17989_/D
+ sky130_fd_sc_hd__a22o_2
XANTENNA__19551__CLK _19706_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19727_ _19828_/CLK _19727_/D vssd1 vssd1 vccd1 vccd1 _19727_/Q sky130_fd_sc_hd__dfxtp_1
X_16939_ _16984_/A vssd1 vssd1 vccd1 vccd1 _16939_/X sky130_fd_sc_hd__buf_1
XFILLER_37_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17281__A _18901_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19658_ _19820_/CLK _19658_/D vssd1 vssd1 vccd1 vccd1 _19658_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10131__A2 _20790_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18609_ _18608_/X _15091_/Y _18906_/S vssd1 vssd1 vccd1 vccd1 _18609_/X sky130_fd_sc_hd__mux2_1
XFILLER_53_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19589_ _20142_/CLK _19589_/D vssd1 vssd1 vccd1 vccd1 _19589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20234__RESET_B repeater203/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18544__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18316__S _18907_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20502_ _21375_/CLK _20502_/D repeater257/X vssd1 vssd1 vccd1 vccd1 _20502_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_165_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21482_ _21485_/CLK _21482_/D repeater200/X vssd1 vssd1 vccd1 vccd1 _21482_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_147_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20433_ _20937_/CLK _20433_/D repeater278/X vssd1 vssd1 vccd1 vccd1 _20433_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__19195__S1 _20122_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20364_ _20951_/CLK _20364_/D repeater271/X vssd1 vssd1 vccd1 vccd1 _20364_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__21093__RESET_B repeater226/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17456__A _21088_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20295_ _20661_/CLK _20295_/D repeater262/X vssd1 vssd1 vccd1 vccd1 _20295_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_115_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__21022__RESET_B repeater238/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17903__B _17944_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_217_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10950_ _21198_/Q _11863_/A _21200_/Q _11804_/D _10949_/X vssd1 vssd1 vccd1 vccd1
+ _10969_/A sky130_fd_sc_hd__o221a_1
XFILLER_217_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18783__A0 _17079_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17586__A1 _18741_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09609_ _20874_/Q _20873_/Q vssd1 vssd1 vccd1 vccd1 _13383_/A sky130_fd_sc_hd__or2_4
XFILLER_243_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10881_ _10890_/A vssd1 vssd1 vccd1 vccd1 _10881_/X sky130_fd_sc_hd__buf_1
XFILLER_32_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_243_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12620_ _12620_/A vssd1 vssd1 vccd1 vccd1 _12620_/X sky130_fd_sc_hd__buf_1
XFILLER_231_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18535__A0 _18848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12551_ _20898_/Q _12543_/X _12550_/X _12546_/X vssd1 vssd1 vccd1 vccd1 _20898_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18226__S _18236_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11502_ _15382_/A vssd1 vssd1 vccd1 vccd1 _11502_/X sky130_fd_sc_hd__buf_4
XPHY_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15270_ _20470_/Q vssd1 vssd1 vccd1 vccd1 _15270_/Y sky130_fd_sc_hd__inv_2
X_12482_ _12474_/A _12474_/B _12479_/Y _12445_/X vssd1 vssd1 vccd1 vccd1 _20926_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_200_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11433_ _11390_/C _11401_/X _11389_/A _11404_/X vssd1 vssd1 vccd1 vccd1 _21172_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19186__S1 _20124_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14221_ _14076_/A _14076_/B _14219_/Y _14207_/X vssd1 vssd1 vccd1 vccd1 _20265_/D
+ sky130_fd_sc_hd__a211oi_4
XPHY_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14152_ _20552_/Q vssd1 vssd1 vccd1 vccd1 _18003_/A sky130_fd_sc_hd__inv_2
X_11364_ _11364_/A _21178_/Q _11363_/A vssd1 vssd1 vccd1 vccd1 _11364_/X sky130_fd_sc_hd__or3b_1
XFILLER_164_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19057__S _19058_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10315_ _10289_/A _20733_/Q _21374_/Q _10312_/Y _10314_/X vssd1 vssd1 vccd1 vccd1
+ _10323_/B sky130_fd_sc_hd__o221a_1
X_13103_ _20634_/Q _13098_/X _12884_/X _13099_/X vssd1 vssd1 vccd1 vccd1 _20634_/D
+ sky130_fd_sc_hd__a22o_1
X_18960_ _16638_/X _21076_/Q _18962_/S vssd1 vssd1 vccd1 vccd1 _18960_/X sky130_fd_sc_hd__mux2_1
X_14083_ _14083_/A _14083_/B vssd1 vssd1 vccd1 vccd1 _14204_/A sky130_fd_sc_hd__or2_1
X_11295_ _20917_/Q _20902_/Q _11307_/C _11306_/C vssd1 vssd1 vccd1 vccd1 _11311_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_152_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13034_ _13040_/A vssd1 vssd1 vccd1 vccd1 _13034_/X sky130_fd_sc_hd__buf_1
X_17911_ _17852_/X _17904_/X _17906_/X _17910_/Y vssd1 vssd1 vccd1 vccd1 _17911_/Y
+ sky130_fd_sc_hd__o211ai_4
X_10246_ _21357_/Q vssd1 vssd1 vccd1 vccd1 _10272_/A sky130_fd_sc_hd__inv_2
X_18891_ _18890_/X _17183_/Y _18891_/S vssd1 vssd1 vccd1 vccd1 _18891_/X sky130_fd_sc_hd__mux2_1
XANTENNA__18896__S _18896_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17842_ _18590_/X _18024_/A _18610_/X _18019_/A vssd1 vssd1 vccd1 vccd1 _17842_/X
+ sky130_fd_sc_hd__o22a_2
XANTENNA__10897__B1 _10896_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10177_ _10177_/A vssd1 vssd1 vccd1 vccd1 _10177_/X sky130_fd_sc_hd__buf_2
XFILLER_66_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17773_ _19316_/Q _17773_/B vssd1 vssd1 vccd1 vccd1 _17773_/X sky130_fd_sc_hd__or2_1
XANTENNA__17813__B _18666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14985_ _20095_/Q _14984_/Y _14973_/X _14874_/B vssd1 vssd1 vccd1 vccd1 _20095_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_19_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19512_ _19784_/CLK _19512_/D vssd1 vssd1 vccd1 vccd1 _19512_/Q sky130_fd_sc_hd__dfxtp_1
X_16724_ _20986_/Q _11992_/B _11993_/B vssd1 vssd1 vccd1 vccd1 _16724_/X sky130_fd_sc_hd__a21bo_1
X_13936_ _20638_/Q vssd1 vssd1 vccd1 vccd1 _13936_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18774__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10113__A2 _20777_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19443_ _19834_/CLK _19443_/D vssd1 vssd1 vccd1 vccd1 _19443_/Q sky130_fd_sc_hd__dfxtp_1
X_16655_ _16661_/A _18953_/X vssd1 vssd1 vccd1 vccd1 _19861_/D sky130_fd_sc_hd__and2_1
XFILLER_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13867_ _20297_/Q vssd1 vssd1 vccd1 vccd1 _14013_/A sky130_fd_sc_hd__inv_2
XFILLER_62_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15606_ _19720_/Q _15603_/X _15483_/X _15604_/X vssd1 vssd1 vccd1 vccd1 _19720_/D
+ sky130_fd_sc_hd__a22o_1
X_19374_ _19706_/CLK _19374_/D vssd1 vssd1 vccd1 vccd1 _19374_/Q sky130_fd_sc_hd__dfxtp_1
X_12818_ _13048_/A _17212_/A vssd1 vssd1 vccd1 vccd1 _12973_/A sky130_fd_sc_hd__or2_1
X_16586_ _21151_/Q _19879_/D _16566_/C _16551_/Y _11577_/A vssd1 vssd1 vccd1 vccd1
+ _16587_/B sky130_fd_sc_hd__o32a_1
XFILLER_90_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13798_ _13793_/Y _20181_/Q _20602_/Q _14569_/A _13797_/X vssd1 vssd1 vccd1 vccd1
+ _13811_/B sky130_fd_sc_hd__o221a_1
XFILLER_203_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18325_ _18324_/X _15137_/Y _18784_/S vssd1 vssd1 vccd1 vccd1 _18325_/X sky130_fd_sc_hd__mux2_1
X_15537_ _15537_/A vssd1 vssd1 vccd1 vccd1 _15537_/X sky130_fd_sc_hd__buf_1
X_12749_ _12734_/A _12748_/X _12745_/X vssd1 vssd1 vccd1 vccd1 _20806_/D sky130_fd_sc_hd__a21boi_1
XFILLER_231_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18136__S _18908_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18256_ _18845_/A0 _13749_/Y _18896_/S vssd1 vssd1 vccd1 vccd1 _18256_/X sky130_fd_sc_hd__mux2_1
XFILLER_147_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15468_ _15479_/A vssd1 vssd1 vccd1 vccd1 _15468_/X sky130_fd_sc_hd__buf_1
XANTENNA__16552__A2 _16550_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17207_ _18898_/X _17205_/X _17206_/Y _17157_/D vssd1 vssd1 vccd1 vccd1 _17207_/X
+ sky130_fd_sc_hd__o22a_1
X_14419_ _14414_/Y _20209_/Q _14415_/Y _20224_/Q _14418_/X vssd1 vssd1 vccd1 vccd1
+ _14420_/D sky130_fd_sc_hd__o221a_1
XANTENNA__19177__S1 _20122_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18829__A1 _19251_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18187_ _18186_/X _10626_/Y _18891_/S vssd1 vssd1 vccd1 vccd1 _18187_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15399_ _15405_/A vssd1 vssd1 vccd1 vccd1 _15406_/A sky130_fd_sc_hd__inv_2
XANTENNA__19999__RESET_B repeater225/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17138_ _17387_/A vssd1 vssd1 vccd1 vccd1 _17139_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17069_ _20258_/Q _20256_/Q vssd1 vssd1 vccd1 vccd1 _17069_/X sky130_fd_sc_hd__or2_1
X_09960_ _21424_/Q _09957_/X _09693_/X _09958_/X vssd1 vssd1 vccd1 vccd1 _21424_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__15512__B1 _15456_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20080_ _20088_/CLK _20080_/D repeater259/X vssd1 vssd1 vccd1 vccd1 _20080_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_98_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09891_ _20011_/Q _09885_/B _09886_/A vssd1 vssd1 vccd1 vccd1 _17025_/A sky130_fd_sc_hd__o21ai_1
XFILLER_69_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_214_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_238_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20982_ _20982_/CLK _20982_/D repeater187/X vssd1 vssd1 vccd1 vccd1 _20982_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__20415__RESET_B repeater185/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17568__A1 _16550_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15579__B1 _15544_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_225_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12883__A _15354_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19168__S1 _20122_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21274__RESET_B repeater245/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14554__A1 _20131_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_239_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21465_ _21477_/CLK _21465_/D repeater205/X vssd1 vssd1 vccd1 vccd1 _21465_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_193_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20416_ _20957_/CLK _20416_/D repeater185/X vssd1 vssd1 vccd1 vccd1 _20416_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_4_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21396_ _21401_/CLK _21396_/D repeater253/X vssd1 vssd1 vccd1 vccd1 _21396_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_190_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20347_ _20949_/CLK _20347_/D repeater269/X vssd1 vssd1 vccd1 vccd1 _20347_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_161_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10100_ _20775_/Q vssd1 vssd1 vccd1 vccd1 _10100_/Y sky130_fd_sc_hd__inv_2
XFILLER_122_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11080_ _11080_/A vssd1 vssd1 vccd1 vccd1 _11081_/B sky130_fd_sc_hd__inv_2
XFILLER_122_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20278_ _20286_/CLK _20278_/D repeater262/X vssd1 vssd1 vccd1 vccd1 _20278_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_248_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10031_ _21402_/Q vssd1 vssd1 vccd1 vccd1 _10162_/C sky130_fd_sc_hd__inv_2
XANTENNA__13219__A input47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_1_1_0_HCLK_A clkbuf_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14770_ _20129_/Q _14769_/Y _14763_/Y _14534_/X vssd1 vssd1 vccd1 vccd1 _20129_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_44_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11982_ _10988_/X _11981_/X _21018_/Q _11981_/X vssd1 vssd1 vccd1 vccd1 _11983_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_217_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13721_ _15758_/A _15762_/A _13725_/S vssd1 vssd1 vccd1 vccd1 _20330_/D sky130_fd_sc_hd__mux2_1
XFILLER_232_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10933_ _21197_/Q vssd1 vssd1 vccd1 vccd1 _10933_/Y sky130_fd_sc_hd__inv_2
XFILLER_217_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16440_ _19313_/Q _16434_/X _16332_/X _16436_/X vssd1 vssd1 vccd1 vccd1 _19313_/D
+ sky130_fd_sc_hd__a22o_1
X_10864_ _10871_/A vssd1 vssd1 vccd1 vccd1 _10864_/X sky130_fd_sc_hd__buf_1
X_13652_ _13652_/A vssd1 vssd1 vccd1 vccd1 _13652_/X sky130_fd_sc_hd__buf_1
XFILLER_220_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18508__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12603_ _17060_/C _12600_/X _18223_/X _12601_/X vssd1 vssd1 vccd1 vccd1 _20871_/D
+ sky130_fd_sc_hd__a22o_1
X_16371_ _16371_/A vssd1 vssd1 vccd1 vccd1 _16371_/X sky130_fd_sc_hd__buf_1
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10795_ _10827_/A vssd1 vssd1 vccd1 vccd1 _10795_/X sky130_fd_sc_hd__buf_2
X_13583_ _20407_/Q _13580_/X _13432_/X _13581_/X vssd1 vssd1 vccd1 vccd1 _20407_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18110_ _17366_/Y _20129_/Q _20241_/Q _17275_/Y vssd1 vssd1 vccd1 vccd1 _18110_/X
+ sky130_fd_sc_hd__o22a_1
X_15322_ _20032_/Q _09690_/X _13538_/X _09694_/X vssd1 vssd1 vccd1 vccd1 _20032_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12534_ _11310_/B _12527_/X _11301_/B _12528_/X vssd1 vssd1 vccd1 vccd1 _20908_/D
+ sky130_fd_sc_hd__o22ai_1
X_19090_ _19308_/Q _21056_/Q _19872_/Q vssd1 vssd1 vccd1 vccd1 _19090_/X sky130_fd_sc_hd__mux2_1
XPHY_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19159__S1 _21017_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18041_ _18335_/X _17954_/X _18341_/X _17955_/X vssd1 vssd1 vccd1 vccd1 _18042_/D
+ sky130_fd_sc_hd__a22o_2
X_15253_ _20492_/Q vssd1 vssd1 vccd1 vccd1 _15253_/Y sky130_fd_sc_hd__inv_2
XFILLER_149_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12465_ _12465_/A vssd1 vssd1 vccd1 vccd1 _12465_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_repeater149_A _17281_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14204_ _14204_/A vssd1 vssd1 vccd1 vccd1 _14204_/Y sky130_fd_sc_hd__inv_2
X_11416_ _11416_/A vssd1 vssd1 vccd1 vccd1 _21181_/D sky130_fd_sc_hd__inv_2
XFILLER_138_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15184_ _15184_/A vssd1 vssd1 vccd1 vccd1 _15184_/Y sky130_fd_sc_hd__inv_2
X_12396_ _12396_/A _12396_/B _12490_/C vssd1 vssd1 vccd1 vccd1 _12469_/C sky130_fd_sc_hd__or3_1
XFILLER_126_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11347_ _21177_/Q _11347_/B _11373_/C vssd1 vssd1 vccd1 vccd1 _11410_/C sky130_fd_sc_hd__nor3_4
X_14135_ _20550_/Q vssd1 vssd1 vccd1 vccd1 _17977_/A sky130_fd_sc_hd__inv_2
X_19992_ _21055_/CLK _19992_/D repeater221/X vssd1 vssd1 vccd1 vccd1 _19992_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_140_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10582__A2 _20744_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11278_ _11541_/C _11541_/A _11541_/B _11280_/A vssd1 vssd1 vccd1 vccd1 _12502_/A
+ sky130_fd_sc_hd__and4b_1
X_18943_ _16697_/X _20898_/Q _18946_/S vssd1 vssd1 vccd1 vccd1 _18943_/X sky130_fd_sc_hd__mux2_1
X_14066_ _20262_/Q vssd1 vssd1 vccd1 vccd1 _14073_/A sky130_fd_sc_hd__inv_2
XFILLER_113_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13017_ _20682_/Q _13012_/X _12932_/X _13013_/X vssd1 vssd1 vccd1 vccd1 _20682_/D
+ sky130_fd_sc_hd__a22o_1
X_10229_ _21374_/Q vssd1 vssd1 vccd1 vccd1 _10289_/A sky130_fd_sc_hd__inv_2
X_18874_ _18873_/X _17191_/Y _18874_/S vssd1 vssd1 vccd1 vccd1 _18874_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11531__A1 _21142_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17825_ _18271_/X _17574_/A _18328_/X _17576_/A vssd1 vssd1 vccd1 vccd1 _17825_/Y
+ sky130_fd_sc_hd__a22oi_4
XFILLER_239_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12968__A _12968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17756_ _18677_/X _17775_/B vssd1 vssd1 vccd1 vccd1 _17756_/Y sky130_fd_sc_hd__nand2_1
XFILLER_47_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14968_ _14968_/A vssd1 vssd1 vccd1 vccd1 _14968_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16707_ _16709_/A _18939_/X vssd1 vssd1 vccd1 vccd1 _19897_/D sky130_fd_sc_hd__and2_1
XFILLER_207_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13919_ _20641_/Q vssd1 vssd1 vccd1 vccd1 _13919_/Y sky130_fd_sc_hd__inv_2
XFILLER_208_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17687_ _19452_/Q vssd1 vssd1 vccd1 vccd1 _17687_/Y sky130_fd_sc_hd__inv_2
X_14899_ _14895_/Y _20092_/Q _14896_/Y _20086_/Q _14898_/X vssd1 vssd1 vccd1 vccd1
+ _14901_/C sky130_fd_sc_hd__a221o_1
XANTENNA__20257__SET_B repeater217/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19426_ _20331_/CLK _19426_/D vssd1 vssd1 vccd1 vccd1 _19426_/Q sky130_fd_sc_hd__dfxtp_1
X_16638_ _19854_/Q _15288_/B _15289_/B vssd1 vssd1 vccd1 vccd1 _16638_/X sky130_fd_sc_hd__a21bo_1
XFILLER_35_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17970__A1 _18207_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19357_ _21338_/CLK _19357_/D vssd1 vssd1 vccd1 vccd1 _19357_/Q sky130_fd_sc_hd__dfxtp_1
X_16569_ _16569_/A _16569_/B _16569_/C _16569_/D vssd1 vssd1 vccd1 vccd1 _16569_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_200_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18308_ _18307_/X _10284_/A _18886_/S vssd1 vssd1 vccd1 vccd1 _18308_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12795__B1 _12697_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19288_ _21338_/CLK _21185_/Q vssd1 vssd1 vccd1 vccd1 _19288_/Q sky130_fd_sc_hd__dfxtp_1
X_18239_ _20863_/Q input13/X _18242_/S vssd1 vssd1 vccd1 vccd1 _18239_/X sky130_fd_sc_hd__mux2_1
XFILLER_175_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12547__B1 _12544_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21250_ _21390_/CLK _21250_/D repeater239/X vssd1 vssd1 vccd1 vccd1 _21250_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_172_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20201_ _20626_/CLK _20201_/D repeater193/X vssd1 vssd1 vccd1 vccd1 _20201_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_132_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21181_ _21183_/CLK _21181_/D repeater216/X vssd1 vssd1 vccd1 vccd1 _21181_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_116_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20132_ _20136_/CLK _20132_/D repeater249/X vssd1 vssd1 vccd1 vccd1 _20132_/Q sky130_fd_sc_hd__dfrtp_2
X_09943_ _10908_/A _10026_/B _17370_/A vssd1 vssd1 vccd1 vccd1 _09944_/S sky130_fd_sc_hd__or3_1
XFILLER_131_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20667__RESET_B repeater207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_225_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20063_ _20066_/CLK _20063_/D repeater281/X vssd1 vssd1 vccd1 vccd1 _20063_/Q sky130_fd_sc_hd__dfrtp_1
X_09874_ _21442_/Q _09871_/A _09870_/X _09847_/A _09873_/X vssd1 vssd1 vccd1 vccd1
+ _09875_/A sky130_fd_sc_hd__o32a_1
XFILLER_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12878__A _16338_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater240 repeater241/X vssd1 vssd1 vccd1 vccd1 repeater240/X sky130_fd_sc_hd__buf_6
Xrepeater251 repeater256/X vssd1 vssd1 vccd1 vccd1 repeater251/X sky130_fd_sc_hd__buf_8
Xrepeater262 repeater263/X vssd1 vssd1 vccd1 vccd1 repeater262/X sky130_fd_sc_hd__buf_8
Xrepeater273 repeater274/X vssd1 vssd1 vccd1 vccd1 repeater273/X sky130_fd_sc_hd__buf_6
XPHY_4405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20965_ _20981_/CLK _20965_/D repeater186/X vssd1 vssd1 vccd1 vccd1 _20965_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_241_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_199_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_202_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20896_ _21141_/CLK _20896_/D repeater192/X vssd1 vssd1 vccd1 vccd1 _20896_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_241_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21455__RESET_B repeater245/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10580_ _21313_/Q _10578_/Y _10534_/A _20766_/Q _10579_/Y vssd1 vssd1 vccd1 vccd1
+ _10591_/A sky130_fd_sc_hd__o221a_1
XFILLER_110_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18910__A0 _18909_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18504__S _18617_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12250_ _20933_/Q vssd1 vssd1 vccd1 vccd1 _12422_/A sky130_fd_sc_hd__inv_2
X_21448_ _21449_/CLK _21448_/D repeater248/X vssd1 vssd1 vccd1 vccd1 _21448_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_119_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11201_ _12898_/B vssd1 vssd1 vccd1 vccd1 _17553_/A sky130_fd_sc_hd__buf_2
XANTENNA__11210__B1 _09645_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12181_ _12320_/A _20349_/Q _20955_/Q _12180_/Y vssd1 vssd1 vccd1 vccd1 _12181_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__15429__A _15429_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21379_ _21379_/CLK _21379_/D repeater213/X vssd1 vssd1 vccd1 vccd1 _21379_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_135_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11132_ _21005_/Q _11128_/X _16465_/A _15756_/A _11951_/B vssd1 vssd1 vccd1 vccd1
+ _11132_/X sky130_fd_sc_hd__a32o_1
XFILLER_135_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15940_ _19563_/Q _15935_/X _15893_/X _15937_/X vssd1 vssd1 vccd1 vccd1 _19563_/D
+ sky130_fd_sc_hd__a22o_1
X_11063_ _11063_/A _11063_/B vssd1 vssd1 vccd1 vccd1 _11066_/A sky130_fd_sc_hd__or2_1
XFILLER_103_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10014_ _21418_/Q _17035_/A _21418_/Q _17035_/A vssd1 vssd1 vccd1 vccd1 _10014_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_15871_ _15871_/A vssd1 vssd1 vccd1 vccd1 _15871_/X sky130_fd_sc_hd__buf_1
XFILLER_95_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17610_ _18740_/X _17703_/B vssd1 vssd1 vccd1 vccd1 _17610_/Y sky130_fd_sc_hd__nand2_1
X_14822_ _20109_/Q _20110_/Q _14823_/S vssd1 vssd1 vccd1 vccd1 _20110_/D sky130_fd_sc_hd__mux2_1
X_18590_ _18589_/X _12236_/Y _18907_/S vssd1 vssd1 vccd1 vccd1 _18590_/X sky130_fd_sc_hd__mux2_1
XFILLER_236_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17541_ _17541_/A _17542_/B vssd1 vssd1 vccd1 vccd1 _17541_/Y sky130_fd_sc_hd__nor2_1
X_14753_ _14753_/A _14753_/B vssd1 vssd1 vccd1 vccd1 _14754_/A sky130_fd_sc_hd__or2_1
X_11965_ _18975_/S _16525_/C vssd1 vssd1 vccd1 vccd1 _13717_/C sky130_fd_sc_hd__or2_1
XFILLER_151_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19070__S _19908_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13704_ _15421_/A vssd1 vssd1 vccd1 vccd1 _13704_/X sky130_fd_sc_hd__buf_4
XANTENNA__10739__C _16777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10916_ _20168_/Q vssd1 vssd1 vccd1 vccd1 _14679_/A sky130_fd_sc_hd__inv_2
X_17472_ _17472_/A vssd1 vssd1 vccd1 vccd1 _17472_/X sky130_fd_sc_hd__buf_1
XFILLER_232_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14684_ _20168_/Q _14673_/A _14682_/A vssd1 vssd1 vccd1 vccd1 _20168_/D sky130_fd_sc_hd__o21a_1
XANTENNA__19762__CLK _21009_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11896_ _11896_/A _11896_/B vssd1 vssd1 vccd1 vccd1 _11897_/A sky130_fd_sc_hd__or2_1
X_19211_ _19207_/X _19208_/X _19209_/X _19210_/X _20132_/Q _20133_/Q vssd1 vssd1 vccd1
+ vccd1 _19211_/X sky130_fd_sc_hd__mux4_2
X_16423_ _19324_/Q _16420_/X _15865_/A _16422_/X vssd1 vssd1 vccd1 vccd1 _19324_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_232_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21196__RESET_B repeater218/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13635_ _20379_/Q _13632_/X _13418_/X _13634_/X vssd1 vssd1 vccd1 vccd1 _20379_/D
+ sky130_fd_sc_hd__a22o_1
X_10847_ _10853_/A vssd1 vssd1 vccd1 vccd1 _10847_/X sky130_fd_sc_hd__buf_1
XFILLER_220_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_repeater266_A repeater267/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19142_ _19681_/Q _19809_/Q _19801_/Q _19793_/Q _19285_/S0 _21017_/Q vssd1 vssd1
+ vccd1 vccd1 _19142_/X sky130_fd_sc_hd__mux4_2
X_16354_ _19361_/Q _16352_/X _16288_/X _16353_/X vssd1 vssd1 vccd1 vccd1 _19361_/D
+ sky130_fd_sc_hd__a22o_1
X_13566_ _13566_/A vssd1 vssd1 vccd1 vccd1 _13566_/X sky130_fd_sc_hd__buf_1
XFILLER_81_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09642__B1 _09641_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10778_ _10778_/A _10797_/A vssd1 vssd1 vccd1 vccd1 _10779_/B sky130_fd_sc_hd__or2_2
XFILLER_8_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15305_ _15305_/A vssd1 vssd1 vccd1 vccd1 _15305_/X sky130_fd_sc_hd__buf_1
XFILLER_158_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12517_ _12520_/A vssd1 vssd1 vccd1 vccd1 _12518_/A sky130_fd_sc_hd__buf_1
XFILLER_185_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19073_ _16730_/X _21137_/Q _19908_/D vssd1 vssd1 vccd1 vccd1 _19073_/X sky130_fd_sc_hd__mux2_1
XFILLER_200_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16285_ _20328_/Q vssd1 vssd1 vccd1 vccd1 _16285_/X sky130_fd_sc_hd__buf_1
X_13497_ _20446_/Q _13492_/X _13424_/X _13494_/X vssd1 vssd1 vccd1 vccd1 _20446_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18414__S _18835_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18024_ _18024_/A vssd1 vssd1 vccd1 vccd1 _18024_/X sky130_fd_sc_hd__buf_1
X_15236_ _20483_/Q _15076_/A _20493_/Q _15086_/A _15235_/X vssd1 vssd1 vccd1 vccd1
+ _15250_/A sky130_fd_sc_hd__o221a_1
XFILLER_60_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12448_ _12462_/A vssd1 vssd1 vccd1 vccd1 _12448_/X sky130_fd_sc_hd__buf_1
XFILLER_154_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15167_ _15029_/A _15165_/Y _15166_/X _15088_/B vssd1 vssd1 vccd1 vccd1 _20073_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_99_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12379_ _12097_/X _12312_/B _12364_/X _12377_/Y vssd1 vssd1 vccd1 vccd1 _20958_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_114_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14118_ _18080_/A _20288_/Q _20537_/Q _14077_/A vssd1 vssd1 vccd1 vccd1 _14118_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_125_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19975_ _20422_/CLK _19975_/D repeater188/X vssd1 vssd1 vccd1 vccd1 _19975_/Q sky130_fd_sc_hd__dfrtp_1
X_15098_ _20063_/Q vssd1 vssd1 vccd1 vccd1 _15098_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_101_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20078__RESET_B repeater259/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18926_ _17113_/Y _17110_/Y _18926_/S vssd1 vssd1 vccd1 vccd1 _18926_/X sky130_fd_sc_hd__mux2_1
X_14049_ _20279_/Q vssd1 vssd1 vccd1 vccd1 _14089_/A sky130_fd_sc_hd__inv_2
XFILLER_141_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_126_HCLK_A clkbuf_4_4_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20007__RESET_B repeater238/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18857_ _17280_/X _21413_/Q _20870_/Q vssd1 vssd1 vccd1 vccd1 _18857_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17808_ _17808_/A vssd1 vssd1 vccd1 vccd1 _17812_/B sky130_fd_sc_hd__buf_2
X_18788_ _18787_/X _12209_/Y _18910_/S vssd1 vssd1 vccd1 vccd1 _18788_/X sky130_fd_sc_hd__mux2_1
XANTENNA__15505__C _15505_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_224_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17739_ _19645_/Q vssd1 vssd1 vccd1 vccd1 _17739_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18196__A1 _10606_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20750_ _21294_/CLK _20750_/D repeater210/X vssd1 vssd1 vccd1 vccd1 _20750_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_23_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19409_ _21222_/CLK _19409_/D vssd1 vssd1 vccd1 vccd1 _19409_/Q sky130_fd_sc_hd__dfxtp_1
X_20681_ _21357_/CLK _20681_/D repeater199/X vssd1 vssd1 vccd1 vccd1 _20681_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_189_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12768__B1 _12666_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19240__S0 _20130_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18324__S _18908_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21302_ _21302_/CLK _21302_/D repeater208/X vssd1 vssd1 vccd1 vccd1 _21302_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_164_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_50_HCLK clkbuf_4_9_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _21134_/CLK sky130_fd_sc_hd__clkbuf_16
X_21233_ _21234_/CLK _21233_/D repeater270/X vssd1 vssd1 vccd1 vccd1 _21233_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_116_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12940__B1 _12855_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21164_ _21164_/CLK _21164_/D repeater226/X vssd1 vssd1 vccd1 vccd1 _21164_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_49_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20115_ _21419_/CLK _20115_/D repeater234/X vssd1 vssd1 vccd1 vccd1 _20115_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_120_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09926_ _21433_/Q _21434_/Q _09929_/S vssd1 vssd1 vccd1 vccd1 _21434_/D sky130_fd_sc_hd__mux2_1
X_21095_ _21151_/CLK _21095_/D repeater226/X vssd1 vssd1 vccd1 vccd1 _21095_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__13496__A1 _20447_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20430__RESET_B repeater190/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20046_ _20066_/CLK _20046_/D repeater281/X vssd1 vssd1 vccd1 vccd1 _20046_/Q sky130_fd_sc_hd__dfrtp_4
X_09857_ _09857_/A vssd1 vssd1 vccd1 vccd1 _09859_/A sky130_fd_sc_hd__inv_2
XFILLER_100_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09788_ _09780_/A _16619_/B input74/X _18963_/X vssd1 vssd1 vccd1 vccd1 _09788_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA_clkbuf_leaf_48_HCLK_A clkbuf_opt_4_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18187__A1 _10626_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ _21055_/Q _11749_/Y _19308_/Q _11749_/A _11327_/X vssd1 vssd1 vccd1 vccd1
+ _21055_/D sky130_fd_sc_hd__o221a_1
XPHY_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_242_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20762__CLK _21342_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20948_ _20949_/CLK _20948_/D repeater269/X vssd1 vssd1 vccd1 vccd1 _20948_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10701_ _10723_/A _10722_/A _10701_/C vssd1 vssd1 vccd1 vccd1 _10720_/A sky130_fd_sc_hd__or3_1
XFILLER_42_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11681_ _11689_/A vssd1 vssd1 vccd1 vccd1 _11690_/A sky130_fd_sc_hd__inv_2
XPHY_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20879_ _21459_/CLK _20879_/D repeater244/X vssd1 vssd1 vccd1 vccd1 _20879_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13420_ _13447_/A vssd1 vssd1 vccd1 vccd1 _13420_/X sky130_fd_sc_hd__buf_1
X_10632_ _21338_/Q _10631_/Y _10703_/A _20743_/Q vssd1 vssd1 vccd1 vccd1 _10632_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19231__S0 _20132_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10563_ _21329_/Q vssd1 vssd1 vccd1 vccd1 _10658_/A sky130_fd_sc_hd__inv_2
XANTENNA__17639__A _17639_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13351_ _13351_/A vssd1 vssd1 vccd1 vccd1 _13351_/X sky130_fd_sc_hd__buf_1
XANTENNA__18234__S _18236_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12302_ _12302_/A _12302_/B _12302_/C _12302_/D vssd1 vssd1 vccd1 vccd1 _12453_/A
+ sky130_fd_sc_hd__and4_2
X_16070_ _19498_/Q _16064_/X _15766_/X _16066_/X vssd1 vssd1 vccd1 vccd1 _19498_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_input77_A sda_i_S4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13282_ input55/X vssd1 vssd1 vccd1 vccd1 _13282_/X sky130_fd_sc_hd__clkbuf_2
X_10494_ _21299_/Q _18005_/A _10775_/A _20688_/Q vssd1 vssd1 vccd1 vccd1 _10494_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_136_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15021_ _15021_/A _15021_/B _15025_/C vssd1 vssd1 vccd1 vccd1 _20079_/D sky130_fd_sc_hd__nor3_1
XFILLER_154_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12233_ _20931_/Q vssd1 vssd1 vccd1 vccd1 _12420_/A sky130_fd_sc_hd__inv_2
XANTENNA__12931__B1 _12930_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12164_ _20347_/Q vssd1 vssd1 vccd1 vccd1 _12164_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19065__S _19910_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11115_ _11109_/B _11114_/X _11051_/X _11101_/X _11052_/D vssd1 vssd1 vccd1 vccd1
+ _11116_/A sky130_fd_sc_hd__o32a_1
X_16972_ _19970_/Q _16979_/B vssd1 vssd1 vccd1 vccd1 _16972_/Y sky130_fd_sc_hd__nor2_1
X_12095_ _20962_/Q _20376_/Q _12093_/X _12094_/Y vssd1 vssd1 vccd1 vccd1 _12103_/B
+ sky130_fd_sc_hd__o22a_1
X_19760_ _19765_/CLK _19760_/D vssd1 vssd1 vccd1 vccd1 _19760_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__20171__RESET_B repeater190/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18711_ _18845_/A0 _17635_/Y _18879_/S vssd1 vssd1 vccd1 vccd1 _18711_/X sky130_fd_sc_hd__mux2_1
X_11046_ _21242_/Q _11045_/X _11024_/Y vssd1 vssd1 vccd1 vccd1 _21242_/D sky130_fd_sc_hd__o21a_1
X_15923_ _19573_/Q _15920_/X _15887_/X _15922_/X vssd1 vssd1 vccd1 vccd1 _19573_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_39_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20100__RESET_B repeater259/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19691_ _19813_/CLK _19691_/D vssd1 vssd1 vccd1 vccd1 _19691_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15228__A2 _15099_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18642_ _18641_/X _14891_/Y _18907_/S vssd1 vssd1 vccd1 vccd1 _18642_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15854_ _19603_/Q _15849_/X _15733_/X _15851_/X vssd1 vssd1 vccd1 vccd1 _19603_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_37_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14436__B1 _14435_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14805_ _14791_/Y _14807_/B _14804_/A _19125_/S _14804_/Y vssd1 vssd1 vccd1 vccd1
+ _14805_/X sky130_fd_sc_hd__a32o_1
XFILLER_206_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18573_ _17830_/X _09721_/Y _18928_/S vssd1 vssd1 vccd1 vccd1 _18573_/X sky130_fd_sc_hd__mux2_1
X_15785_ _15785_/A vssd1 vssd1 vccd1 vccd1 _15785_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__18409__S _18669_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12997_ _13013_/A vssd1 vssd1 vccd1 vccd1 _12997_/X sky130_fd_sc_hd__buf_1
XFILLER_17_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16718__A _16718_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12998__B1 _12996_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17524_ _19466_/Q vssd1 vssd1 vccd1 vccd1 _17524_/Y sky130_fd_sc_hd__inv_2
XFILLER_91_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14736_ _20141_/Q _14731_/X _13710_/X _14733_/X vssd1 vssd1 vccd1 vccd1 _20141_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_45_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11948_ _11917_/X _11934_/Y _11947_/X _11943_/X _11932_/X vssd1 vssd1 vccd1 vccd1
+ _21008_/D sky130_fd_sc_hd__a32o_1
XFILLER_221_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17455_ _21059_/Q vssd1 vssd1 vccd1 vccd1 _17455_/Y sky130_fd_sc_hd__inv_2
X_14667_ _20175_/Q _14666_/X _20175_/Q _14666_/X vssd1 vssd1 vccd1 vccd1 _20175_/D
+ sky130_fd_sc_hd__o2bb2a_1
X_11879_ _21020_/Q vssd1 vssd1 vccd1 vccd1 _11881_/A sky130_fd_sc_hd__buf_1
XFILLER_232_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16406_ _16413_/A vssd1 vssd1 vccd1 vccd1 _16406_/X sky130_fd_sc_hd__buf_1
X_13618_ _20388_/Q _13613_/X _13557_/X _13614_/X vssd1 vssd1 vccd1 vccd1 _20388_/D
+ sky130_fd_sc_hd__a22o_1
X_17386_ _21129_/Q vssd1 vssd1 vccd1 vccd1 _17386_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19222__S0 _19275_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14598_ _14642_/A vssd1 vssd1 vccd1 vccd1 _14624_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_158_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_73_HCLK clkbuf_opt_7_HCLK/X vssd1 vssd1 vccd1 vccd1 _20626_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_146_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19125_ _16481_/Y _14313_/Y _19125_/S vssd1 vssd1 vccd1 vccd1 _19125_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16337_ _19369_/Q _16334_/X _16335_/X _16336_/X vssd1 vssd1 vccd1 vccd1 _19369_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_146_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13549_ _13566_/A vssd1 vssd1 vccd1 vccd1 _13549_/X sky130_fd_sc_hd__buf_1
XANTENNA__18144__S _18748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16453__A _16459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19056_ _16758_/Y _20813_/Q _19058_/S vssd1 vssd1 vccd1 vccd1 _19920_/D sky130_fd_sc_hd__mux2_1
XFILLER_9_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16268_ _19402_/Q _16262_/X _16117_/X _16264_/X vssd1 vssd1 vccd1 vccd1 _19402_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_134_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18007_ _20833_/Q _18007_/B vssd1 vssd1 vccd1 vccd1 _18007_/Y sky130_fd_sc_hd__nand2_1
X_15219_ _20471_/Q _15065_/A _15218_/Y _20044_/Q vssd1 vssd1 vccd1 vccd1 _15219_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__18090__D _18090_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16199_ _19437_/Q _16195_/X _16196_/X _16198_/X vssd1 vssd1 vccd1 vccd1 _19437_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18102__A1 _18649_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20259__RESET_B repeater262/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10528__A2 _10375_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19958_ _20422_/CLK _19958_/D repeater184/X vssd1 vssd1 vccd1 vccd1 _19958_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_113_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09711_ _18965_/X vssd1 vssd1 vccd1 vccd1 _09812_/A sky130_fd_sc_hd__inv_2
X_18909_ _18908_/X _12201_/Y _18909_/S vssd1 vssd1 vccd1 vccd1 _18909_/X sky130_fd_sc_hd__mux2_1
X_19889_ _21338_/CLK _19889_/D repeater221/X vssd1 vssd1 vccd1 vccd1 _19889_/Q sky130_fd_sc_hd__dfstp_1
X_09642_ _21478_/Q _09632_/X _09641_/X _09634_/X vssd1 vssd1 vccd1 vccd1 _21478_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_110_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18319__S _18908_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__21047__RESET_B repeater226/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20802_ _21407_/CLK _20802_/D repeater252/X vssd1 vssd1 vccd1 vccd1 _20802_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_42_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20733_ _21375_/CLK _20733_/D repeater257/X vssd1 vssd1 vccd1 vccd1 _20733_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14148__A _20541_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13052__A _13072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20664_ _20665_/CLK _20664_/D repeater261/X vssd1 vssd1 vccd1 vccd1 _20664_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_51_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19213__S0 _19275_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20595_ _20665_/CLK _20595_/D repeater259/X vssd1 vssd1 vccd1 vccd1 _20595_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12891__A _13600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20682__RESET_B repeater208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_247_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11716__A1 _16663_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12913__B1 _12668_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21216_ _21223_/CLK _21216_/D repeater238/X vssd1 vssd1 vccd1 vccd1 _21216_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_116_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21147_ _21147_/CLK _21147_/D repeater212/X vssd1 vssd1 vccd1 vccd1 _21147_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_120_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09909_ _21253_/Q _17020_/A vssd1 vssd1 vccd1 vccd1 _09909_/Y sky130_fd_sc_hd__nand2_1
X_21078_ _21087_/CLK _21078_/D repeater227/X vssd1 vssd1 vccd1 vccd1 _21078_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_47_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12920_ input51/X vssd1 vssd1 vccd1 vccd1 _12920_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__17604__B1 _21007_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20029_ _21357_/CLK _20029_/D repeater199/X vssd1 vssd1 vccd1 vccd1 _20029_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_46_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21470__RESET_B repeater204/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12851_ _12876_/A vssd1 vssd1 vccd1 vccd1 _12851_/X sky130_fd_sc_hd__buf_1
XFILLER_46_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18229__S _18236_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11802_ _11816_/A vssd1 vssd1 vccd1 vccd1 _11827_/A sky130_fd_sc_hd__buf_1
XPHY_4054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15570_ _19737_/Q _15568_/X _15518_/X _15569_/X vssd1 vssd1 vccd1 vccd1 _19737_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12782_ _20789_/Q _12777_/X _09638_/X _12778_/X vssd1 vssd1 vccd1 vccd1 _20789_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_203_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_96_HCLK clkbuf_4_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20286_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_4087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19865__RESET_B repeater225/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14521_ _14521_/A vssd1 vssd1 vccd1 vccd1 _14524_/A sky130_fd_sc_hd__inv_2
XPHY_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11733_ _13163_/A vssd1 vssd1 vccd1 vccd1 _11733_/X sky130_fd_sc_hd__clkbuf_2
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_214_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18580__A1 _14435_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17240_ _19359_/Q vssd1 vssd1 vccd1 vccd1 _17240_/Y sky130_fd_sc_hd__inv_2
X_14452_ _14566_/B vssd1 vssd1 vccd1 vccd1 _14477_/A sky130_fd_sc_hd__buf_1
XFILLER_186_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11664_ _21071_/Q vssd1 vssd1 vccd1 vccd1 _16654_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__19204__S0 _19275_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13403_ _20489_/Q _13398_/X _13284_/X _13399_/X vssd1 vssd1 vccd1 vccd1 _20489_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10615_ _20768_/Q vssd1 vssd1 vccd1 vccd1 _10615_/Y sky130_fd_sc_hd__inv_2
XPHY_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17171_ _17163_/X _17168_/X _17170_/X vssd1 vssd1 vccd1 vccd1 _17171_/Y sky130_fd_sc_hd__a21oi_1
X_14383_ _14383_/A vssd1 vssd1 vccd1 vccd1 _14383_/Y sky130_fd_sc_hd__inv_2
XFILLER_195_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11595_ _11591_/A _11591_/B _11583_/B _11586_/A vssd1 vssd1 vccd1 vccd1 _21121_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16122_ _19473_/Q _16119_/X _16120_/X _16121_/X vssd1 vssd1 vccd1 vccd1 _19473_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13334_ _13352_/A vssd1 vssd1 vccd1 vccd1 _13334_/X sky130_fd_sc_hd__buf_1
X_10546_ _10705_/A _10704_/A _10703_/A _10700_/A vssd1 vssd1 vccd1 vccd1 _10552_/C
+ sky130_fd_sc_hd__or4_4
XFILLER_116_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18899__S _18899_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_2_HCLK clkbuf_opt_0_HCLK/A vssd1 vssd1 vccd1 vccd1 _19706_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_127_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13157__B1 _13032_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16053_ _19508_/Q _16049_/X _15762_/X _16051_/X vssd1 vssd1 vccd1 vccd1 _19508_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_157_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13265_ input62/X vssd1 vssd1 vccd1 vccd1 _13265_/X sky130_fd_sc_hd__clkbuf_2
X_10477_ _21298_/Q _10472_/Y _21294_/Q _17942_/A _10476_/X vssd1 vssd1 vccd1 vccd1
+ _10496_/A sky130_fd_sc_hd__o221a_1
XFILLER_182_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15004_ _15004_/A _15004_/B vssd1 vssd1 vccd1 vccd1 _15009_/A sky130_fd_sc_hd__or2_1
XFILLER_124_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12216_ _20919_/Q vssd1 vssd1 vccd1 vccd1 _12490_/C sky130_fd_sc_hd__inv_2
XANTENNA__17816__B _17944_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13196_ _20596_/Q _13192_/X _12984_/X _13195_/X vssd1 vssd1 vccd1 vccd1 _20596_/D
+ sky130_fd_sc_hd__a22o_1
X_19812_ _19812_/CLK _19812_/D vssd1 vssd1 vccd1 vccd1 _19812_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_0_HCLK_A HCLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12147_ _20333_/Q vssd1 vssd1 vccd1 vccd1 _12147_/Y sky130_fd_sc_hd__inv_2
XFILLER_173_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19743_ _21121_/CLK _19743_/D vssd1 vssd1 vccd1 vccd1 _19743_/Q sky130_fd_sc_hd__dfxtp_1
X_12078_ _20972_/Q _18000_/A _12333_/A _20394_/Q vssd1 vssd1 vccd1 vccd1 _12078_/X
+ sky130_fd_sc_hd__o22a_1
X_16955_ _16958_/A _16958_/C _16954_/Y _16950_/Y vssd1 vssd1 vccd1 vccd1 _16956_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11029_ _19955_/Q _16901_/A vssd1 vssd1 vccd1 vccd1 _16905_/A sky130_fd_sc_hd__or2_1
X_15906_ _15912_/A vssd1 vssd1 vccd1 vccd1 _15906_/X sky130_fd_sc_hd__buf_1
XFILLER_238_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16886_ _16886_/A vssd1 vssd1 vccd1 vccd1 _16892_/A sky130_fd_sc_hd__buf_1
X_19674_ _19812_/CLK _19674_/D vssd1 vssd1 vccd1 vccd1 _19674_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15837_ _19613_/Q _15834_/X _09818_/X _15836_/X vssd1 vssd1 vccd1 vccd1 _19613_/D
+ sky130_fd_sc_hd__a22o_1
X_18625_ _18084_/Y _16871_/Y _18667_/S vssd1 vssd1 vccd1 vccd1 _18625_/X sky130_fd_sc_hd__mux2_1
XANTENNA__18139__S _18896_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_31_HCLK_A clkbuf_opt_4_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15352__A _15429_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18556_ _17830_/X _10941_/Y _18928_/S vssd1 vssd1 vccd1 vccd1 _18556_/X sky130_fd_sc_hd__mux2_1
X_15768_ _15768_/A vssd1 vssd1 vccd1 vccd1 _15768_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_45_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_94_HCLK_A clkbuf_4_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_221_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11643__B1 _21103_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14719_ _20151_/Q _14717_/X _14258_/X _14718_/X vssd1 vssd1 vccd1 vccd1 _20151_/D
+ sky130_fd_sc_hd__a22o_1
X_17507_ _19586_/Q vssd1 vssd1 vccd1 vccd1 _17507_/Y sky130_fd_sc_hd__inv_2
X_18487_ _17079_/Y _15278_/Y _18908_/S vssd1 vssd1 vccd1 vccd1 _18487_/X sky130_fd_sc_hd__mux2_1
X_15699_ _19673_/Q _15696_/X _15697_/X _15698_/X vssd1 vssd1 vccd1 vccd1 _19673_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_221_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17438_ _19617_/Q vssd1 vssd1 vccd1 vccd1 _17438_/Y sky130_fd_sc_hd__inv_2
XFILLER_159_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13396__B1 _13272_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17369_ _19311_/Q _17369_/B vssd1 vssd1 vccd1 vccd1 _17369_/Y sky130_fd_sc_hd__nor2_1
X_19108_ _19118_/S _11986_/Y _19115_/S vssd1 vssd1 vccd1 vccd1 _19108_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13600__A _13600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20380_ _20480_/CLK _20380_/D repeater183/X vssd1 vssd1 vccd1 vccd1 _20380_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_174_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19039_ _16832_/X _20830_/Q _19046_/S vssd1 vssd1 vccd1 vccd1 _19937_/D sky130_fd_sc_hd__mux2_1
XFILLER_174_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput100 _18090_/X vssd1 vssd1 vccd1 vccd1 HRDATA[29] sky130_fd_sc_hd__clkbuf_2
XANTENNA__18602__S _18904_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput111 _19985_/Q vssd1 vssd1 vccd1 vccd1 HREADYOUT sky130_fd_sc_hd__clkbuf_2
Xoutput122 _17061_/X vssd1 vssd1 vccd1 vccd1 IRQ[4] sky130_fd_sc_hd__clkbuf_2
Xoutput133 _21410_/Q vssd1 vssd1 vccd1 vccd1 SCLK_S3 sky130_fd_sc_hd__clkbuf_2
Xoutput144 _21042_/Q vssd1 vssd1 vccd1 vccd1 sda_oen_o_S4 sky130_fd_sc_hd__clkbuf_2
X_21001_ _21001_/CLK _21001_/D repeater190/X vssd1 vssd1 vccd1 vccd1 _21001_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_233_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13320__B1 _13163_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__21228__RESET_B repeater249/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09625_ _21485_/Q _09620_/X _09621_/X _09624_/X vssd1 vssd1 vccd1 vccd1 _21485_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_56_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12886__A _13104_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_243_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16358__A _19888_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19823__CLK _21452_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20716_ _21357_/CLK _20716_/D repeater199/X vssd1 vssd1 vccd1 vccd1 _20716_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_211_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13387__A0 _13254_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20647_ _21486_/CLK _20647_/D repeater198/X vssd1 vssd1 vccd1 vccd1 _20647_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_183_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10400_ _21357_/Q _10399_/Y _10395_/X _10273_/B vssd1 vssd1 vccd1 vccd1 _21357_/D
+ sky130_fd_sc_hd__o211a_1
X_11380_ _11388_/A _11386_/B _21184_/Q _11385_/D vssd1 vssd1 vccd1 vccd1 _11384_/C
+ sky130_fd_sc_hd__or4_4
X_20578_ _20946_/CLK _20578_/D repeater274/X vssd1 vssd1 vccd1 vccd1 _20578_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_137_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10331_ _21367_/Q _10330_/Y _10271_/A _20715_/Q vssd1 vssd1 vccd1 vccd1 _10331_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_125_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18512__S _18875_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13050_ _13657_/A _13259_/B vssd1 vssd1 vccd1 vccd1 _13078_/A sky130_fd_sc_hd__or2_2
X_10262_ _10262_/A _10262_/B vssd1 vssd1 vccd1 vccd1 _10415_/A sky130_fd_sc_hd__or2_1
XFILLER_117_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12001_ _20995_/Q _12001_/B vssd1 vssd1 vccd1 vccd1 _12002_/B sky130_fd_sc_hd__or2_1
XFILLER_105_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10193_ _10193_/A vssd1 vssd1 vccd1 vccd1 _10193_/Y sky130_fd_sc_hd__inv_2
XFILLER_120_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16740_ _16740_/A _18931_/X vssd1 vssd1 vccd1 vccd1 _19912_/D sky130_fd_sc_hd__and2_1
XFILLER_19_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13952_ _20651_/Q _13884_/A _20639_/Q _14012_/A vssd1 vssd1 vccd1 vccd1 _13952_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_235_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12903_ _12936_/A vssd1 vssd1 vccd1 vccd1 _12926_/A sky130_fd_sc_hd__buf_1
X_16671_ _21159_/Q _11447_/B _11448_/B vssd1 vssd1 vccd1 vccd1 _16671_/X sky130_fd_sc_hd__a21bo_1
XFILLER_74_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13883_ _13883_/A _13883_/B vssd1 vssd1 vccd1 vccd1 _13999_/A sky130_fd_sc_hd__or2_1
XFILLER_19_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18410_ _18409_/X _20190_/Q _18748_/S vssd1 vssd1 vccd1 vccd1 _18410_/X sky130_fd_sc_hd__mux2_2
X_15622_ _19711_/Q _15618_/X _15485_/X _15619_/X vssd1 vssd1 vccd1 vccd1 _19711_/D
+ sky130_fd_sc_hd__a22o_1
X_12834_ _20762_/Q _12829_/X _12670_/X _12830_/X vssd1 vssd1 vccd1 vccd1 _20762_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19390_ _19813_/CLK _19390_/D vssd1 vssd1 vccd1 vccd1 _19390_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_234_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18341_ _18340_/X _20200_/Q _18748_/S vssd1 vssd1 vccd1 vccd1 _18341_/X sky130_fd_sc_hd__mux2_1
XFILLER_187_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15553_ _15553_/A vssd1 vssd1 vccd1 vccd1 _15553_/X sky130_fd_sc_hd__buf_1
XPHY_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12765_ _12777_/A vssd1 vssd1 vccd1 vccd1 _12765_/X sky130_fd_sc_hd__buf_1
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_repeater179_A _18242_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_230_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14504_ _14504_/A _14504_/B vssd1 vssd1 vccd1 vccd1 _14504_/Y sky130_fd_sc_hd__nor2_2
XPHY_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11716_ _16663_/A _11713_/X _11680_/X _11715_/X vssd1 vssd1 vccd1 vccd1 _21071_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18272_ _17079_/Y _15253_/Y _18908_/S vssd1 vssd1 vccd1 vccd1 _18272_/X sky130_fd_sc_hd__mux2_1
XFILLER_187_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15484_ _19776_/Q _15479_/X _15483_/X _15481_/X vssd1 vssd1 vccd1 vccd1 _19776_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_14_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12696_ _20821_/Q _12693_/X _09659_/X _12694_/X vssd1 vssd1 vccd1 vccd1 _20821_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17223_ _17223_/A vssd1 vssd1 vccd1 vccd1 _17932_/A sky130_fd_sc_hd__clkbuf_2
XPHY_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14435_ _21474_/Q vssd1 vssd1 vccd1 vccd1 _14435_/Y sky130_fd_sc_hd__inv_2
XFILLER_175_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11647_ _18980_/X _11640_/X _21100_/Q _11646_/X vssd1 vssd1 vccd1 vccd1 _21100_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput13 HADDR[20] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__clkbuf_1
XPHY_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13420__A _13447_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17154_ _17390_/A vssd1 vssd1 vccd1 vccd1 _17154_/X sky130_fd_sc_hd__clkbuf_2
Xinput24 HADDR[30] vssd1 vssd1 vccd1 vccd1 input24/X sky130_fd_sc_hd__buf_1
X_14366_ _14462_/B _14366_/B vssd1 vssd1 vccd1 vccd1 _14490_/A sky130_fd_sc_hd__or2_1
XFILLER_11_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput35 HSEL vssd1 vssd1 vccd1 vccd1 hold9/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__16316__B1 _16235_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11578_ _12515_/A vssd1 vssd1 vccd1 vccd1 _16541_/A sky130_fd_sc_hd__buf_1
XFILLER_10_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput46 HWDATA[17] vssd1 vssd1 vccd1 vccd1 input46/X sky130_fd_sc_hd__clkbuf_4
Xinput57 HWDATA[27] vssd1 vssd1 vccd1 vccd1 input57/X sky130_fd_sc_hd__clkbuf_4
X_16105_ _19479_/Q _16101_/X _15881_/X _16102_/X vssd1 vssd1 vccd1 vccd1 _19479_/D
+ sky130_fd_sc_hd__a22o_1
Xinput68 HWDATA[8] vssd1 vssd1 vccd1 vccd1 input68/X sky130_fd_sc_hd__buf_2
XFILLER_156_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13317_ _20537_/Q _13315_/X _13240_/X _13316_/X vssd1 vssd1 vccd1 vccd1 _20537_/D
+ sky130_fd_sc_hd__a22o_1
X_10529_ _21340_/Q vssd1 vssd1 vccd1 vccd1 _10575_/A sky130_fd_sc_hd__inv_2
X_17085_ _17085_/A vssd1 vssd1 vccd1 vccd1 _18910_/S sky130_fd_sc_hd__inv_16
XFILLER_183_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14297_ _20126_/Q vssd1 vssd1 vccd1 vccd1 _15335_/A sky130_fd_sc_hd__inv_2
XANTENNA__18422__S _18667_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16036_ _16042_/A vssd1 vssd1 vccd1 vccd1 _16043_/A sky130_fd_sc_hd__inv_2
XFILLER_6_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_103_HCLK clkbuf_4_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20088_/CLK sky130_fd_sc_hd__clkbuf_16
X_13248_ _13248_/A vssd1 vssd1 vccd1 vccd1 _13248_/X sky130_fd_sc_hd__buf_1
XANTENNA__17546__B _18879_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13179_ _13182_/A _13179_/B input73/X vssd1 vssd1 vccd1 vccd1 _13521_/A sky130_fd_sc_hd__and3_1
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17987_ _18292_/X _17951_/X _18251_/X _17952_/X vssd1 vssd1 vccd1 vccd1 _17989_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_85_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__21321__RESET_B repeater205/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19726_ _19828_/CLK _19726_/D vssd1 vssd1 vccd1 vccd1 _19726_/Q sky130_fd_sc_hd__dfxtp_1
X_16938_ _19962_/Q _16930_/A _19963_/Q vssd1 vssd1 vccd1 vccd1 _16938_/X sky130_fd_sc_hd__o21a_1
XFILLER_96_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17281__B _18899_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19657_ _21021_/CLK _19657_/D vssd1 vssd1 vccd1 vccd1 _19657_/Q sky130_fd_sc_hd__dfxtp_1
X_16869_ _19946_/Q _16868_/A _16867_/Y _16868_/Y vssd1 vssd1 vccd1 vccd1 _16870_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_38_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18608_ _17079_/Y _15257_/Y _18908_/S vssd1 vssd1 vccd1 vccd1 _18608_/X sky130_fd_sc_hd__mux2_1
XFILLER_92_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19588_ _21218_/CLK _19588_/D vssd1 vssd1 vccd1 vccd1 _19588_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14802__B1 _20119_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_240_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18539_ _17281_/X _17922_/Y _18835_/S vssd1 vssd1 vccd1 vccd1 _18539_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13369__B1 _13311_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_221_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20501_ _20929_/CLK _20501_/D repeater265/X vssd1 vssd1 vccd1 vccd1 _20501_/Q sky130_fd_sc_hd__dfrtp_2
X_21481_ _21481_/CLK _21481_/D repeater200/X vssd1 vssd1 vccd1 vccd1 _21481_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20274__RESET_B repeater263/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13330__A _13357_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20432_ _20432_/CLK _20432_/D repeater235/X vssd1 vssd1 vccd1 vccd1 _20432_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_147_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20203__RESET_B repeater193/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20363_ _20951_/CLK _20363_/D repeater272/X vssd1 vssd1 vccd1 vccd1 _20363_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_174_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18332__S _18666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20294_ _20661_/CLK _20294_/D repeater262/X vssd1 vssd1 vccd1 vccd1 _20294_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__15257__A _20474_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21409__RESET_B repeater233/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19376__CLK _19706_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_7_0_HCLK_A clkbuf_3_7_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09608_ _20870_/Q _11187_/A vssd1 vssd1 vccd1 vccd1 _11489_/C sky130_fd_sc_hd__or2_1
X_10880_ _10880_/A vssd1 vssd1 vccd1 vccd1 _10890_/A sky130_fd_sc_hd__inv_2
XFILLER_244_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18507__S _18886_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12550_ _12550_/A vssd1 vssd1 vccd1 vccd1 _12550_/X sky130_fd_sc_hd__clkbuf_2
XPHY_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11501_ _11486_/X _11487_/X _19111_/S _16548_/A _11500_/Y vssd1 vssd1 vccd1 vccd1
+ _21151_/D sky130_fd_sc_hd__a32o_1
XPHY_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12481_ _20927_/Q _12479_/Y _12476_/B _12480_/X vssd1 vssd1 vccd1 vccd1 _20927_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18299__A0 _17281_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13240__A _14258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14220_ _20266_/Q _14219_/Y _14205_/X _14078_/B vssd1 vssd1 vccd1 vccd1 _20266_/D
+ sky130_fd_sc_hd__o211a_1
X_11432_ _11432_/A vssd1 vssd1 vccd1 vccd1 _21173_/D sky130_fd_sc_hd__inv_2
XPHY_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_126_HCLK clkbuf_4_4_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20408_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_153_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14151_ _20534_/Q vssd1 vssd1 vccd1 vccd1 _17541_/A sky130_fd_sc_hd__inv_2
XFILLER_138_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11363_ _11363_/A _11363_/B _11364_/A vssd1 vssd1 vccd1 vccd1 _11365_/A sky130_fd_sc_hd__nor3_2
XANTENNA__18242__S _18242_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13102_ _20635_/Q _13098_/X _12881_/X _13099_/X vssd1 vssd1 vccd1 vccd1 _20635_/D
+ sky130_fd_sc_hd__a22o_1
X_10314_ _10285_/A _20729_/Q _21355_/Q _10313_/Y vssd1 vssd1 vccd1 vccd1 _10314_/X
+ sky130_fd_sc_hd__o22a_1
X_14082_ _14082_/A _14209_/A vssd1 vssd1 vccd1 vccd1 _14083_/B sky130_fd_sc_hd__or2_1
X_11294_ _11294_/A _11299_/D vssd1 vssd1 vccd1 vccd1 _11306_/C sky130_fd_sc_hd__or2_1
XFILLER_3_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13033_ _20674_/Q _13026_/X _13032_/X _13027_/X vssd1 vssd1 vccd1 vccd1 _20674_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11695__A _12715_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17910_ _18465_/X _17907_/X _18456_/X _17908_/X _17909_/X vssd1 vssd1 vccd1 vccd1
+ _17910_/Y sky130_fd_sc_hd__a221oi_2
X_10245_ _21358_/Q vssd1 vssd1 vccd1 vccd1 _10273_/A sky130_fd_sc_hd__inv_2
X_18890_ _18889_/X _10459_/Y _18896_/S vssd1 vssd1 vccd1 vccd1 _18890_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17841_ _17857_/A vssd1 vssd1 vccd1 vccd1 _18024_/A sky130_fd_sc_hd__clkbuf_2
X_10176_ _10162_/A _10175_/A _21401_/Q _10175_/Y _10166_/X vssd1 vssd1 vccd1 vccd1
+ _21401_/D sky130_fd_sc_hd__o221a_1
XFILLER_120_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19073__S _19908_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17772_ _19469_/Q vssd1 vssd1 vccd1 vccd1 _17772_/Y sky130_fd_sc_hd__inv_2
X_14984_ _14984_/A vssd1 vssd1 vccd1 vccd1 _14984_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19880__RESET_B repeater212/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19511_ _21462_/CLK _19511_/D vssd1 vssd1 vccd1 vccd1 _19511_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_247_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16723_ _20985_/Q _11991_/B _11992_/B vssd1 vssd1 vccd1 vccd1 _16723_/X sky130_fd_sc_hd__a21bo_1
XFILLER_47_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13935_ _20662_/Q vssd1 vssd1 vccd1 vccd1 _13935_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16654_ _16654_/A vssd1 vssd1 vccd1 vccd1 _16661_/A sky130_fd_sc_hd__buf_1
X_19442_ _20136_/CLK _19442_/D vssd1 vssd1 vccd1 vccd1 _19442_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_235_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13866_ _20298_/Q vssd1 vssd1 vccd1 vccd1 _14014_/A sky130_fd_sc_hd__inv_2
XFILLER_222_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13599__B1 _13454_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15605_ _19721_/Q _15603_/X _15480_/X _15604_/X vssd1 vssd1 vccd1 vccd1 _19721_/D
+ sky130_fd_sc_hd__a22o_1
X_12817_ _13047_/A _13047_/B _13327_/C vssd1 vssd1 vccd1 vccd1 _17212_/A sky130_fd_sc_hd__or3_4
X_16585_ _16585_/A _16744_/B _16585_/C vssd1 vssd1 vccd1 vccd1 _19991_/D sky130_fd_sc_hd__nand3_1
X_19373_ _19777_/CLK _19373_/D vssd1 vssd1 vccd1 vccd1 _19373_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13797_ _20622_/Q _14588_/A _13796_/Y _20188_/Q vssd1 vssd1 vccd1 vccd1 _13797_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_15_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18417__S _18874_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20714__RESET_B repeater254/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17329__A2 _17298_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18324_ _17079_/Y _15246_/Y _18908_/S vssd1 vssd1 vccd1 vccd1 _18324_/X sky130_fd_sc_hd__mux2_1
X_15536_ _15536_/A vssd1 vssd1 vccd1 vccd1 _15536_/X sky130_fd_sc_hd__buf_1
XFILLER_203_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12748_ _12748_/A _12751_/B vssd1 vssd1 vccd1 vccd1 _12748_/X sky130_fd_sc_hd__or2_1
XFILLER_187_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18255_ _18254_/X _10780_/A _18898_/S vssd1 vssd1 vccd1 vccd1 _18255_/X sky130_fd_sc_hd__mux2_1
X_15467_ _15610_/A _16215_/B _16297_/C vssd1 vssd1 vccd1 vccd1 _15479_/A sky130_fd_sc_hd__or3_4
XANTENNA__14246__A _14246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12679_ _12679_/A vssd1 vssd1 vccd1 vccd1 _12679_/X sky130_fd_sc_hd__buf_1
XFILLER_175_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17206_ _18912_/X vssd1 vssd1 vccd1 vccd1 _17206_/Y sky130_fd_sc_hd__inv_2
X_14418_ _20240_/Q _14416_/Y _20232_/Q _14417_/Y vssd1 vssd1 vccd1 vccd1 _14418_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_30_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18186_ _18845_/A0 _10428_/Y _18896_/S vssd1 vssd1 vccd1 vccd1 _18186_/X sky130_fd_sc_hd__mux2_1
X_15398_ _15405_/A vssd1 vssd1 vccd1 vccd1 _15398_/X sky130_fd_sc_hd__buf_1
X_17137_ _21056_/Q vssd1 vssd1 vccd1 vccd1 _17137_/Y sky130_fd_sc_hd__inv_2
XFILLER_116_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14349_ _20211_/Q vssd1 vssd1 vccd1 vccd1 _14351_/B sky130_fd_sc_hd__inv_2
XANTENNA__18152__S _18784_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17068_ _20255_/Q _20253_/Q _20254_/Q _17067_/X vssd1 vssd1 vccd1 vccd1 _19886_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_6_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16019_ _21221_/Q vssd1 vssd1 vccd1 vccd1 _16107_/B sky130_fd_sc_hd__buf_1
XFILLER_98_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09890_ _21258_/Q vssd1 vssd1 vccd1 vccd1 _09890_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19968__RESET_B repeater185/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_214_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18214__A0 _18848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19709_ _19777_/CLK _19709_/D vssd1 vssd1 vccd1 vccd1 _19709_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_4609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20981_ _20981_/CLK _20981_/D repeater187/X vssd1 vssd1 vccd1 vccd1 _20981_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_65_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16636__A _16663_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18327__S _18885_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_149_HCLK clkbuf_4_4_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _21234_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_159_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13060__A _13072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21464_ _21481_/CLK _21464_/D repeater206/X vssd1 vssd1 vccd1 vccd1 _21464_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_119_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20415_ _20957_/CLK _20415_/D repeater185/X vssd1 vssd1 vccd1 vccd1 _20415_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_162_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21395_ _21401_/CLK _21395_/D repeater253/X vssd1 vssd1 vccd1 vccd1 _21395_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_135_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20346_ _20930_/CLK _20346_/D repeater269/X vssd1 vssd1 vccd1 vccd1 _20346_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_107_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18997__S _19026_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20277_ _20286_/CLK _20277_/D repeater265/X vssd1 vssd1 vccd1 vccd1 _20277_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_108_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21243__RESET_B repeater190/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10030_ _20736_/Q vssd1 vssd1 vccd1 vccd1 _10220_/A sky130_fd_sc_hd__inv_2
XFILLER_76_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13817__A1 _20603_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18205__A0 _17079_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11981_ _15559_/A _15374_/B _11910_/B vssd1 vssd1 vccd1 vccd1 _11981_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__10859__A _13188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13720_ _20330_/Q vssd1 vssd1 vccd1 vccd1 _15762_/A sky130_fd_sc_hd__buf_1
XFILLER_217_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10932_ _21024_/Q vssd1 vssd1 vccd1 vccd1 _11864_/A sky130_fd_sc_hd__inv_2
XFILLER_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13651_ _13651_/A vssd1 vssd1 vccd1 vccd1 _13651_/X sky130_fd_sc_hd__buf_1
XFILLER_232_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20196__RESET_B repeater193/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10863_ _13384_/C _10908_/B vssd1 vssd1 vccd1 vccd1 _10871_/A sky130_fd_sc_hd__or2_2
XANTENNA__18237__S _18242_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12602_ _20872_/Q _12600_/X _18224_/X _12601_/X vssd1 vssd1 vccd1 vccd1 _20872_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_71_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15450__A _15657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16370_ _16370_/A vssd1 vssd1 vccd1 vccd1 _16370_/X sky130_fd_sc_hd__buf_1
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20125__RESET_B repeater247/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13582_ _20408_/Q _13580_/X _13429_/X _13581_/X vssd1 vssd1 vccd1 vccd1 _20408_/D
+ sky130_fd_sc_hd__a22o_1
X_10794_ _21304_/Q _10793_/Y _10787_/X _10781_/B vssd1 vssd1 vccd1 vccd1 _21304_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15321_ _09851_/X _15320_/Y _10842_/A _15320_/B vssd1 vssd1 vccd1 vccd1 _20033_/D
+ sky130_fd_sc_hd__o22a_1
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12533_ _11313_/B _12518_/A _12503_/B _12521_/X vssd1 vssd1 vccd1 vccd1 _20909_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_185_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18040_ _18372_/X _17951_/X _18316_/X _17952_/X vssd1 vssd1 vccd1 vccd1 _18042_/C
+ sky130_fd_sc_hd__a22o_1
X_15252_ _20496_/Q _20075_/Q _15251_/Y _15090_/Y vssd1 vssd1 vccd1 vccd1 _15259_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_157_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12464_ _12421_/A _12421_/B _12453_/X _12461_/Y vssd1 vssd1 vccd1 vccd1 _20932_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_149_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14203_ _14085_/A _14085_/B _14201_/Y _14193_/X vssd1 vssd1 vccd1 vccd1 _20275_/D
+ sky130_fd_sc_hd__a211oi_4
X_11415_ _11407_/Y _11408_/X _11413_/X _11357_/C _11414_/X vssd1 vssd1 vccd1 vccd1
+ _11416_/A sky130_fd_sc_hd__o32a_1
XANTENNA__19068__S _19908_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11202__B _17553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15183_ _15112_/X _15078_/B _15181_/Y _15179_/X vssd1 vssd1 vccd1 vccd1 _20064_/D
+ sky130_fd_sc_hd__a211oi_2
X_12395_ _12395_/A _12395_/B vssd1 vssd1 vccd1 vccd1 _12433_/A sky130_fd_sc_hd__or2_1
XFILLER_125_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18692__A0 _18848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14134_ _20540_/Q vssd1 vssd1 vccd1 vccd1 _14134_/Y sky130_fd_sc_hd__inv_2
X_11346_ _11390_/A _11348_/C _11346_/C vssd1 vssd1 vccd1 vccd1 _11373_/C sky130_fd_sc_hd__or3_4
X_19991_ _21055_/CLK _19991_/D repeater220/X vssd1 vssd1 vccd1 vccd1 _19991_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_125_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19691__CLK _19813_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18942_ _16699_/X _20899_/Q _18946_/S vssd1 vssd1 vccd1 vccd1 _18942_/X sky130_fd_sc_hd__mux2_1
XFILLER_165_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_repeater211_A repeater212/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14065_ _20263_/Q vssd1 vssd1 vccd1 vccd1 _14074_/A sky130_fd_sc_hd__inv_2
X_11277_ _11304_/D vssd1 vssd1 vccd1 vccd1 _11280_/A sky130_fd_sc_hd__buf_1
XANTENNA__18700__S _18910_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13016_ _20683_/Q _13012_/X _12930_/X _13013_/X vssd1 vssd1 vccd1 vccd1 _20683_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18444__A0 _18443_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10228_ _10221_/A _10221_/B _21376_/Q _10145_/A _10170_/X vssd1 vssd1 vccd1 vccd1
+ _21376_/D sky130_fd_sc_hd__o221a_1
X_18873_ _18872_/X _17192_/Y _18901_/S vssd1 vssd1 vccd1 vccd1 _18873_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15625__A _15632_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17824_ _18185_/X _17954_/A _18183_/X _17572_/B vssd1 vssd1 vccd1 vccd1 _17827_/B
+ sky130_fd_sc_hd__a22oi_4
XFILLER_0_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10159_ _10159_/A _10159_/B vssd1 vssd1 vccd1 vccd1 _10179_/A sky130_fd_sc_hd__or2_1
XANTENNA__20966__RESET_B repeater186/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17755_ _18678_/X _17774_/B vssd1 vssd1 vccd1 vccd1 _17755_/X sky130_fd_sc_hd__and2_1
X_14967_ _14967_/A _15025_/C _14967_/C vssd1 vssd1 vccd1 vccd1 _20104_/D sky130_fd_sc_hd__nor3_1
XANTENNA__18747__A1 _21467_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16706_ _19897_/Q _14237_/B _14238_/B vssd1 vssd1 vccd1 vccd1 _16706_/X sky130_fd_sc_hd__a21bo_1
XFILLER_81_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17840__A _17928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13918_ _20653_/Q _20310_/Q _13917_/Y _13972_/A vssd1 vssd1 vccd1 vccd1 _13922_/B
+ sky130_fd_sc_hd__o22a_1
X_17686_ _19484_/Q vssd1 vssd1 vccd1 vccd1 _17686_/Y sky130_fd_sc_hd__inv_2
X_14898_ _20587_/Q _14963_/D _14897_/Y _20077_/Q vssd1 vssd1 vccd1 vccd1 _14898_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_63_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19425_ _21222_/CLK _19425_/D vssd1 vssd1 vccd1 vccd1 _19425_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16637_ _16643_/A _18961_/X vssd1 vssd1 vccd1 vccd1 _19853_/D sky130_fd_sc_hd__and2_1
X_13849_ _20312_/Q vssd1 vssd1 vccd1 vccd1 _13971_/A sky130_fd_sc_hd__inv_2
XFILLER_62_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12984__A input62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18147__S _18886_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19356_ _21453_/CLK _19356_/D vssd1 vssd1 vccd1 vccd1 _19356_/Q sky130_fd_sc_hd__dfxtp_1
X_16568_ _16568_/A _16568_/B _16568_/C vssd1 vssd1 vccd1 vccd1 _16569_/B sky130_fd_sc_hd__or3_2
XFILLER_176_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18307_ _18306_/X _10082_/Y _18644_/S vssd1 vssd1 vccd1 vccd1 _18307_/X sky130_fd_sc_hd__mux2_1
X_15519_ _15519_/A vssd1 vssd1 vccd1 vccd1 _15519_/X sky130_fd_sc_hd__buf_1
X_19287_ _20042_/CLK _21043_/Q vssd1 vssd1 vccd1 vccd1 _19287_/Q sky130_fd_sc_hd__dfxtp_1
X_16499_ _16495_/Y _19997_/Q _16496_/Y _16498_/Y vssd1 vssd1 vccd1 vccd1 _16499_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_200_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18238_ _20862_/Q input11/X _18242_/S vssd1 vssd1 vccd1 vccd1 _18238_/X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_149_HCLK_A clkbuf_4_4_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12547__A1 _20900_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17287__A _21057_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18169_ _18848_/A0 _10356_/Y _18884_/S vssd1 vssd1 vccd1 vccd1 _18169_/X sky130_fd_sc_hd__mux2_1
XFILLER_190_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20200_ _20623_/CLK _20200_/D repeater194/X vssd1 vssd1 vccd1 vccd1 _20200_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__18683__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21180_ _21183_/CLK _21180_/D repeater216/X vssd1 vssd1 vccd1 vccd1 _21180_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__15497__B1 _15456_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20131_ _21235_/CLK _20131_/D repeater249/X vssd1 vssd1 vccd1 vccd1 _20131_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_89_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09942_ _17133_/A vssd1 vssd1 vccd1 vccd1 _17370_/A sky130_fd_sc_hd__buf_1
XFILLER_143_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18610__S _18907_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18435__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20062_ _20066_/CLK _20062_/D repeater281/X vssd1 vssd1 vccd1 vccd1 _20062_/Q sky130_fd_sc_hd__dfrtp_2
X_09873_ _14307_/B _09870_/A _09878_/B vssd1 vssd1 vccd1 vccd1 _09873_/X sky130_fd_sc_hd__o21ba_1
XFILLER_100_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater230 repeater231/X vssd1 vssd1 vccd1 vccd1 repeater230/X sky130_fd_sc_hd__clkbuf_8
Xrepeater241 repeater242/X vssd1 vssd1 vccd1 vccd1 repeater241/X sky130_fd_sc_hd__buf_8
XFILLER_239_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrepeater252 repeater255/X vssd1 vssd1 vccd1 vccd1 repeater252/X sky130_fd_sc_hd__buf_8
Xrepeater263 repeater264/X vssd1 vssd1 vccd1 vccd1 repeater263/X sky130_fd_sc_hd__buf_6
Xrepeater274 repeater277/X vssd1 vssd1 vccd1 vccd1 repeater274/X sky130_fd_sc_hd__buf_8
XFILLER_241_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13055__A _13073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20964_ _20981_/CLK _20964_/D repeater186/X vssd1 vssd1 vccd1 vccd1 _20964_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_38_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_242_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_214_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20895_ _21141_/CLK _20895_/D repeater192/X vssd1 vssd1 vccd1 vccd1 _20895_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_80_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19564__CLK _19706_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20541__CLK _20592_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21447_ _21449_/CLK _21447_/D repeater248/X vssd1 vssd1 vccd1 vccd1 _21447_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_182_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11200_ _11200_/A _17838_/A vssd1 vssd1 vccd1 vccd1 _12898_/B sky130_fd_sc_hd__or2_1
X_12180_ _20337_/Q vssd1 vssd1 vccd1 vccd1 _12180_/Y sky130_fd_sc_hd__inv_2
XFILLER_135_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21378_ _21379_/CLK _21378_/D repeater213/X vssd1 vssd1 vccd1 vccd1 _21378_/Q sky130_fd_sc_hd__dfrtp_1
X_11131_ _21005_/Q _11131_/B vssd1 vssd1 vccd1 vccd1 _11951_/B sky130_fd_sc_hd__nand2_1
X_20329_ _20331_/CLK _20329_/D repeater190/X vssd1 vssd1 vccd1 vccd1 _20329_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18520__S _18850_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11062_ _11062_/A _11071_/A vssd1 vssd1 vccd1 vccd1 _11063_/B sky130_fd_sc_hd__or2_1
XFILLER_77_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10013_ _10013_/A _10013_/B vssd1 vssd1 vccd1 vccd1 _17035_/A sky130_fd_sc_hd__or2_1
X_15870_ _19596_/Q _15864_/X _15869_/X _15867_/X vssd1 vssd1 vccd1 vccd1 _19596_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_103_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input22_A HADDR[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14821_ _20110_/Q _20111_/Q _14823_/S vssd1 vssd1 vccd1 vccd1 _20111_/D sky130_fd_sc_hd__mux2_1
XFILLER_236_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20377__RESET_B repeater186/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17540_ _17540_/A _17542_/B vssd1 vssd1 vccd1 vccd1 _17540_/Y sky130_fd_sc_hd__nor2_1
X_14752_ _20132_/Q _14757_/A vssd1 vssd1 vccd1 vccd1 _14753_/B sky130_fd_sc_hd__nand2_1
XFILLER_63_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11964_ _11964_/A vssd1 vssd1 vccd1 vccd1 _18975_/S sky130_fd_sc_hd__buf_2
XFILLER_244_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13703_ _20337_/Q _13699_/X _13511_/X _13700_/X vssd1 vssd1 vccd1 vccd1 _20337_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_189_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17471_ _18790_/X vssd1 vssd1 vccd1 vccd1 _17471_/Y sky130_fd_sc_hd__inv_2
X_10915_ _20169_/Q vssd1 vssd1 vccd1 vccd1 _14680_/A sky130_fd_sc_hd__inv_2
XFILLER_204_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14683_ _10985_/A _14674_/X _20169_/Q _14682_/Y _14680_/X vssd1 vssd1 vccd1 vccd1
+ _20169_/D sky130_fd_sc_hd__o221a_1
XFILLER_189_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11895_ _19114_/X vssd1 vssd1 vccd1 vccd1 _11896_/A sky130_fd_sc_hd__inv_2
XFILLER_189_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output109_A _17828_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19210_ _17698_/Y _17699_/Y _17700_/Y _17701_/Y _20130_/Q _20131_/Q vssd1 vssd1 vccd1
+ vccd1 _19210_/X sky130_fd_sc_hd__mux4_2
XFILLER_71_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16422_ _16428_/A vssd1 vssd1 vccd1 vccd1 _16422_/X sky130_fd_sc_hd__buf_1
X_13634_ _13652_/A vssd1 vssd1 vccd1 vccd1 _13634_/X sky130_fd_sc_hd__buf_1
XFILLER_177_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10846_ _10849_/A vssd1 vssd1 vccd1 vccd1 _10846_/X sky130_fd_sc_hd__buf_1
XFILLER_60_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19141_ _19137_/X _19138_/X _19139_/X _19140_/X _21018_/Q _21019_/Q vssd1 vssd1 vccd1
+ vccd1 _19141_/X sky130_fd_sc_hd__mux4_2
X_16353_ _16353_/A vssd1 vssd1 vccd1 vccd1 _16353_/X sky130_fd_sc_hd__buf_1
XFILLER_158_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13565_ _20417_/Q _13559_/X _13479_/X _13561_/X vssd1 vssd1 vccd1 vccd1 _20417_/D
+ sky130_fd_sc_hd__a22o_1
X_10777_ _10777_/A _10777_/B vssd1 vssd1 vccd1 vccd1 _10797_/A sky130_fd_sc_hd__or2_1
XANTENNA_repeater161_A _18617_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15304_ _20041_/Q _15302_/X _20040_/Q _18962_/S vssd1 vssd1 vccd1 vccd1 _20041_/D
+ sky130_fd_sc_hd__a22o_1
X_12516_ _12528_/A vssd1 vssd1 vccd1 vccd1 _12521_/A sky130_fd_sc_hd__inv_2
X_19072_ _16731_/X _21138_/Q _19908_/D vssd1 vssd1 vccd1 vccd1 _19072_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16284_ _19395_/Q _16276_/X _16283_/X _16279_/X vssd1 vssd1 vccd1 vccd1 _19395_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_9_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13496_ _20447_/Q _13492_/X _13422_/X _13494_/X vssd1 vssd1 vccd1 vccd1 _20447_/D
+ sky130_fd_sc_hd__a22o_1
X_15235_ _15233_/Y _20065_/Q _15234_/Y _20045_/Q vssd1 vssd1 vccd1 vccd1 _15235_/X
+ sky130_fd_sc_hd__o22a_1
X_18023_ _18305_/X _18019_/X _18357_/X _18020_/X _18022_/X vssd1 vssd1 vccd1 vccd1
+ _18027_/B sky130_fd_sc_hd__o221a_2
XANTENNA__21165__RESET_B repeater225/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12447_ _12447_/A vssd1 vssd1 vccd1 vccd1 _12447_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output90_A _17329_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18665__A0 _18848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15166_ _15185_/A vssd1 vssd1 vccd1 vccd1 _15166_/X sky130_fd_sc_hd__buf_1
X_12378_ _12139_/X _12377_/A _20959_/Q _12377_/Y _12206_/X vssd1 vssd1 vccd1 vccd1
+ _20959_/D sky130_fd_sc_hd__o221a_1
XFILLER_125_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14117_ _20559_/Q vssd1 vssd1 vccd1 vccd1 _18080_/A sky130_fd_sc_hd__inv_2
X_11329_ _11390_/A vssd1 vssd1 vccd1 vccd1 _11375_/A sky130_fd_sc_hd__buf_1
X_19974_ _20809_/CLK _19974_/D repeater188/X vssd1 vssd1 vccd1 vccd1 _19974_/Q sky130_fd_sc_hd__dfrtp_1
X_15097_ _20452_/Q vssd1 vssd1 vccd1 vccd1 _15097_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18430__S _18885_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18417__A0 _18848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18925_ _18924_/X _19271_/X _18930_/S vssd1 vssd1 vccd1 vccd1 _18925_/X sky130_fd_sc_hd__mux2_1
X_14048_ _20280_/Q vssd1 vssd1 vccd1 vccd1 _14090_/A sky130_fd_sc_hd__inv_2
XFILLER_122_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_228_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19090__A0 _19308_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15355__A _15592_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18856_ _18855_/X _12265_/Y _18910_/S vssd1 vssd1 vccd1 vccd1 _18856_/X sky130_fd_sc_hd__mux2_1
XFILLER_228_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17807_ _17807_/A _17807_/B vssd1 vssd1 vccd1 vccd1 _17807_/Y sky130_fd_sc_hd__nor2_1
XFILLER_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_4_0_HCLK clkbuf_4_5_0_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_4_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_18787_ _18786_/X _12146_/Y _18787_/S vssd1 vssd1 vccd1 vccd1 _18787_/X sky130_fd_sc_hd__mux2_1
X_15999_ _16034_/A _16229_/B _15999_/C vssd1 vssd1 vccd1 vccd1 _16008_/A sky130_fd_sc_hd__or3_4
XFILLER_48_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_236_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17738_ _19501_/Q vssd1 vssd1 vccd1 vccd1 _17738_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20047__RESET_B repeater281/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_224_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17669_ _19476_/Q vssd1 vssd1 vccd1 vccd1 _17669_/Y sky130_fd_sc_hd__inv_2
XFILLER_196_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13603__A _17080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19408_ _19813_/CLK _19408_/D vssd1 vssd1 vccd1 vccd1 _19408_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20680_ _21357_/CLK _20680_/D repeater199/X vssd1 vssd1 vccd1 vccd1 _20680_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_223_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19339_ _20142_/CLK _19339_/D vssd1 vssd1 vccd1 vccd1 _19339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18605__S _18669_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19240__S1 _20131_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21301_ _21480_/CLK _21301_/D repeater208/X vssd1 vssd1 vccd1 vccd1 _21301_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_117_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19983__RESET_B repeater185/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21232_ _21234_/CLK _21232_/D repeater249/X vssd1 vssd1 vccd1 vccd1 _21232_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_160_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21163_ _21164_/CLK _21163_/D repeater226/X vssd1 vssd1 vccd1 vccd1 _21163_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18340__S _18669_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20888__RESET_B repeater247/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18408__A0 _18407_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09925_ _09925_/A vssd1 vssd1 vccd1 vccd1 _09929_/S sky130_fd_sc_hd__clkbuf_2
X_20114_ _21419_/CLK _20114_/D repeater234/X vssd1 vssd1 vccd1 vccd1 _20114_/Q sky130_fd_sc_hd__dfrtp_1
X_21094_ _21164_/CLK _21094_/D repeater226/X vssd1 vssd1 vccd1 vccd1 _21094_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_59_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20817__RESET_B repeater212/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15890__B1 _15887_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20045_ _20070_/CLK _20045_/D repeater276/X vssd1 vssd1 vccd1 vccd1 _20045_/Q sky130_fd_sc_hd__dfrtp_2
X_09856_ _09840_/X _09849_/X _09855_/X vssd1 vssd1 vccd1 vccd1 _21445_/D sky130_fd_sc_hd__o21a_1
XFILLER_86_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09787_ _09787_/A _09787_/B _18976_/S vssd1 vssd1 vccd1 vccd1 _09787_/X sky130_fd_sc_hd__or3_1
XFILLER_45_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17480__A _17928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17919__C1 _17918_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20947_ _20947_/CLK _20947_/D repeater275/X vssd1 vssd1 vccd1 vccd1 _20947_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_4269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17934__A2 _17203_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10700_ _10700_/A vssd1 vssd1 vccd1 vccd1 _10723_/A sky130_fd_sc_hd__buf_1
XPHY_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ _12544_/A vssd1 vssd1 vccd1 vccd1 _11680_/X sky130_fd_sc_hd__buf_1
XPHY_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20878_ _21459_/CLK _20878_/D repeater243/X vssd1 vssd1 vccd1 vccd1 _20878_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_42_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10631_ _20766_/Q vssd1 vssd1 vccd1 vccd1 _10631_/Y sky130_fd_sc_hd__inv_2
XPHY_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18515__S _18850_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19231__S1 _20133_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13350_ _20518_/Q _13345_/X _13213_/X _13346_/X vssd1 vssd1 vccd1 vccd1 _20518_/D
+ sky130_fd_sc_hd__a22o_1
X_10562_ _21327_/Q vssd1 vssd1 vccd1 vccd1 _10656_/A sky130_fd_sc_hd__inv_2
XFILLER_14_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12301_ _12282_/X _12301_/B _12301_/C _12301_/D vssd1 vssd1 vccd1 vccd1 _12302_/D
+ sky130_fd_sc_hd__and4b_1
XFILLER_154_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_132_HCLK_A clkbuf_4_4_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13281_ _20556_/Q _13276_/X _13280_/X _13278_/X vssd1 vssd1 vccd1 vccd1 _20556_/D
+ sky130_fd_sc_hd__a22o_1
X_10493_ _21299_/Q vssd1 vssd1 vccd1 vccd1 _10775_/A sky130_fd_sc_hd__inv_2
X_15020_ _14853_/B _15022_/A _14853_/A vssd1 vssd1 vccd1 vccd1 _15021_/B sky130_fd_sc_hd__o21a_1
XFILLER_154_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18647__A0 _17079_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12232_ _12232_/A _12232_/B _12232_/C _12232_/D vssd1 vssd1 vccd1 vccd1 _12302_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__11195__B1 _10894_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12163_ _12325_/A _20354_/Q _20972_/Q _12160_/Y _12162_/X vssd1 vssd1 vccd1 vccd1
+ _12175_/A sky130_fd_sc_hd__a221o_1
XFILLER_123_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18250__S _18784_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11114_ _11112_/X _11113_/X _09739_/X _11052_/D vssd1 vssd1 vccd1 vccd1 _11114_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_122_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16971_ _16971_/A vssd1 vssd1 vccd1 vccd1 _17013_/A sky130_fd_sc_hd__clkbuf_2
X_12094_ _20376_/Q vssd1 vssd1 vccd1 vccd1 _12094_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18710_ _18709_/X _16906_/A _18875_/S vssd1 vssd1 vccd1 vccd1 _18710_/X sky130_fd_sc_hd__mux2_2
X_11045_ _19290_/Q _11045_/B vssd1 vssd1 vccd1 vccd1 _11045_/X sky130_fd_sc_hd__and2_1
X_15922_ _15928_/A vssd1 vssd1 vccd1 vccd1 _15922_/X sky130_fd_sc_hd__buf_1
X_19690_ _19813_/CLK _19690_/D vssd1 vssd1 vccd1 vccd1 _19690_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12695__B1 _09655_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18641_ _18640_/X _15122_/Y _18906_/S vssd1 vssd1 vccd1 vccd1 _18641_/X sky130_fd_sc_hd__mux2_2
XFILLER_92_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15853_ _19604_/Q _15849_/X _15730_/X _15851_/X vssd1 vssd1 vccd1 vccd1 _19604_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_65_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19081__S _19908_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14804_ _14804_/A vssd1 vssd1 vccd1 vccd1 _14804_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18572_ _18571_/X _16795_/A _18667_/S vssd1 vssd1 vccd1 vccd1 _18572_/X sky130_fd_sc_hd__mux2_1
XANTENNA__20140__RESET_B repeater250/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15784_ _19635_/Q _15779_/X _15733_/X _15781_/X vssd1 vssd1 vccd1 vccd1 _19635_/D
+ sky130_fd_sc_hd__a22o_1
X_12996_ input57/X vssd1 vssd1 vccd1 vccd1 _12996_/X sky130_fd_sc_hd__buf_2
XFILLER_206_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12998__A1 _20693_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17523_ _19458_/Q vssd1 vssd1 vccd1 vccd1 _17523_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14735_ _20142_/Q _14731_/X _13707_/X _14733_/X vssd1 vssd1 vccd1 vccd1 _20142_/D
+ sky130_fd_sc_hd__a22o_1
X_11947_ _11947_/A _11947_/B vssd1 vssd1 vccd1 vccd1 _11947_/X sky130_fd_sc_hd__or2_1
XFILLER_221_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17454_ _21083_/Q vssd1 vssd1 vccd1 vccd1 _17454_/Y sky130_fd_sc_hd__inv_2
X_14666_ _14534_/X _14660_/Y _19124_/S _14664_/X _14665_/X vssd1 vssd1 vccd1 vccd1
+ _14666_/X sky130_fd_sc_hd__o221a_1
X_11878_ _21021_/Q vssd1 vssd1 vccd1 vccd1 _11878_/Y sky130_fd_sc_hd__inv_2
X_16405_ _16405_/A _16405_/B _16405_/C vssd1 vssd1 vccd1 vccd1 _16413_/A sky130_fd_sc_hd__or3_4
X_13617_ _20389_/Q _13613_/X _13555_/X _13614_/X vssd1 vssd1 vccd1 vccd1 _20389_/D
+ sky130_fd_sc_hd__a22o_1
X_10829_ _10829_/A vssd1 vssd1 vccd1 vccd1 _10829_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21346__RESET_B repeater210/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_12_0_HCLK clkbuf_3_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_12_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_14597_ _14597_/A vssd1 vssd1 vccd1 vccd1 _14642_/A sky130_fd_sc_hd__inv_2
X_17385_ _21138_/Q vssd1 vssd1 vccd1 vccd1 _17385_/Y sky130_fd_sc_hd__inv_2
XFILLER_186_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18425__S _18907_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19222__S1 _21004_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19124_ _19123_/S _14526_/Y _19124_/S vssd1 vssd1 vccd1 vccd1 _19124_/X sky130_fd_sc_hd__mux2_1
X_13548_ _20425_/Q _13537_/X _13547_/X _13541_/X vssd1 vssd1 vccd1 vccd1 _20425_/D
+ sky130_fd_sc_hd__a22o_1
X_16336_ _16336_/A vssd1 vssd1 vccd1 vccd1 _16336_/X sky130_fd_sc_hd__buf_1
XANTENNA__12981__B _13261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19055_ _16763_/X _20814_/Q _19058_/S vssd1 vssd1 vccd1 vccd1 _19921_/D sky130_fd_sc_hd__mux2_1
X_16267_ _19403_/Q _16262_/X _16115_/X _16264_/X vssd1 vssd1 vccd1 vccd1 _19403_/D
+ sky130_fd_sc_hd__a22o_1
X_13479_ input50/X vssd1 vssd1 vccd1 vccd1 _13479_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15218_ _20465_/Q vssd1 vssd1 vccd1 vccd1 _15218_/Y sky130_fd_sc_hd__inv_2
X_18006_ _18006_/A _18006_/B vssd1 vssd1 vccd1 vccd1 _18006_/Y sky130_fd_sc_hd__nor2_1
X_16198_ _16208_/A vssd1 vssd1 vccd1 vccd1 _16198_/X sky130_fd_sc_hd__buf_1
XANTENNA__11186__A0 _11179_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_54_HCLK_A clkbuf_4_12_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15149_ _20434_/Q _15060_/A _20460_/Q _15085_/A vssd1 vssd1 vccd1 vccd1 _15149_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_141_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18160__S _18667_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20981__RESET_B repeater187/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19957_ _20408_/CLK _19957_/D repeater184/X vssd1 vssd1 vccd1 vccd1 _19957_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__20910__RESET_B repeater218/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14675__A1 _10985_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09710_ _16617_/A _09770_/B vssd1 vssd1 vccd1 vccd1 _09787_/A sky130_fd_sc_hd__nor2_1
X_18908_ _17173_/Y _12055_/Y _18908_/S vssd1 vssd1 vccd1 vccd1 _18908_/X sky130_fd_sc_hd__mux2_1
XFILLER_206_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19888_ _21338_/CLK _19888_/D repeater221/X vssd1 vssd1 vccd1 vccd1 _19888_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__20228__RESET_B repeater200/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09641_ _12849_/A vssd1 vssd1 vccd1 vccd1 _09641_/X sky130_fd_sc_hd__buf_4
X_18839_ _18845_/A0 _10347_/Y _18884_/S vssd1 vssd1 vccd1 vccd1 _18839_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20801_ _21407_/CLK _20801_/D repeater252/X vssd1 vssd1 vccd1 vccd1 _20801_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_35_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17916__A2 _17200_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11661__A1 _11502_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20732_ _21366_/CLK _20732_/D repeater257/X vssd1 vssd1 vccd1 vccd1 _20732_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19118__A1 _10985_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20663_ _20665_/CLK _20663_/D repeater261/X vssd1 vssd1 vccd1 vccd1 _20663_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__18335__S _18904_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19213__S1 _21004_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__21016__RESET_B repeater238/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20594_ _20665_/CLK _20594_/D repeater261/X vssd1 vssd1 vccd1 vccd1 _20594_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_167_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21215_ _21223_/CLK _21215_/D repeater240/X vssd1 vssd1 vccd1 vccd1 _21215_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_2_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19752__CLK _19765_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21146_ _21147_/CLK _21146_/D repeater215/X vssd1 vssd1 vccd1 vccd1 _21146_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_132_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09908_ _17022_/A vssd1 vssd1 vccd1 vccd1 _09908_/Y sky130_fd_sc_hd__inv_2
X_21077_ _21087_/CLK _21077_/D repeater227/X vssd1 vssd1 vccd1 vccd1 _21077_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__12677__B1 _09626_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18801__A0 _17281_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17604__A1 _11932_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09839_ _16163_/A _09827_/X _09838_/X _09829_/X vssd1 vssd1 vccd1 vccd1 _21446_/D
+ sky130_fd_sc_hd__a22o_1
X_20028_ _21486_/CLK _20028_/D repeater199/X vssd1 vssd1 vccd1 vccd1 _20028_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_47_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12850_ _12850_/A vssd1 vssd1 vccd1 vccd1 _12876_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_132_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11801_ _11817_/A _12968_/A vssd1 vssd1 vccd1 vccd1 _11816_/A sky130_fd_sc_hd__or2_1
XPHY_4044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12781_ _20790_/Q _12777_/X _09636_/X _12778_/X vssd1 vssd1 vccd1 vccd1 _20790_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14520_ _14520_/A _14520_/B _14524_/C vssd1 vssd1 vccd1 vccd1 _20212_/D sky130_fd_sc_hd__nor3_1
XPHY_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13243__A _14262_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11732_ _21061_/Q _11727_/X _11686_/X _11729_/X vssd1 vssd1 vccd1 vccd1 _21061_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19109__A1 _11123_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14451_ _14464_/B vssd1 vssd1 vccd1 vccd1 _14566_/B sky130_fd_sc_hd__inv_2
XPHY_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11663_ _10892_/A _11652_/X _11658_/A _11659_/Y _21092_/Q vssd1 vssd1 vccd1 vccd1
+ _21092_/D sky130_fd_sc_hd__a32o_1
XPHY_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19204__S1 _21004_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13402_ _20490_/Q _13398_/X _13282_/X _13399_/X vssd1 vssd1 vccd1 vccd1 _20490_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10614_ _20764_/Q vssd1 vssd1 vccd1 vccd1 _10614_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17170_ _17560_/A vssd1 vssd1 vccd1 vccd1 _17170_/X sky130_fd_sc_hd__clkbuf_4
XPHY_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14382_ _14382_/A _14382_/B vssd1 vssd1 vccd1 vccd1 _14383_/A sky130_fd_sc_hd__or2_1
XPHY_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11594_ _21122_/Q _11592_/B _11583_/B _11592_/Y vssd1 vssd1 vccd1 vccd1 _21122_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19287__D _21043_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16121_ _16121_/A vssd1 vssd1 vccd1 vccd1 _16121_/X sky130_fd_sc_hd__buf_1
XFILLER_195_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13333_ _13359_/A vssd1 vssd1 vccd1 vccd1 _13352_/A sky130_fd_sc_hd__clkbuf_2
XPHY_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10545_ _21310_/Q vssd1 vssd1 vccd1 vccd1 _10700_/A sky130_fd_sc_hd__inv_2
XFILLER_6_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_143_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16052_ _19509_/Q _16049_/X _15758_/X _16051_/X vssd1 vssd1 vccd1 vccd1 _19509_/D
+ sky130_fd_sc_hd__a22o_1
X_13264_ _13293_/A vssd1 vssd1 vccd1 vccd1 _13264_/X sky130_fd_sc_hd__buf_1
X_10476_ _10768_/A _20681_/Q _21292_/Q _10475_/Y vssd1 vssd1 vccd1 vccd1 _10476_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__20739__RESET_B repeater205/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15003_ _15003_/A _15012_/A vssd1 vssd1 vccd1 vccd1 _15004_/B sky130_fd_sc_hd__or2_2
XFILLER_124_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19076__S _19908_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12215_ _20924_/Q vssd1 vssd1 vccd1 vccd1 _12256_/A sky130_fd_sc_hd__inv_2
XANTENNA__17385__A _21138_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13195_ _13217_/A vssd1 vssd1 vccd1 vccd1 _13195_/X sky130_fd_sc_hd__buf_1
XFILLER_151_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19811_ _19811_/CLK _19811_/D vssd1 vssd1 vccd1 vccd1 _19811_/Q sky130_fd_sc_hd__dfxtp_1
X_12146_ _20335_/Q vssd1 vssd1 vccd1 vccd1 _12146_/Y sky130_fd_sc_hd__inv_2
XFILLER_173_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13418__A input44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19742_ _21121_/CLK _19742_/D vssd1 vssd1 vccd1 vccd1 _19742_/Q sky130_fd_sc_hd__dfxtp_1
X_12077_ _20980_/Q vssd1 vssd1 vccd1 vccd1 _12333_/A sky130_fd_sc_hd__inv_2
X_16954_ _16958_/A vssd1 vssd1 vccd1 vccd1 _16954_/Y sky130_fd_sc_hd__inv_2
XFILLER_237_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19140__S0 _19285_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15905_ _15911_/A vssd1 vssd1 vccd1 vccd1 _15912_/A sky130_fd_sc_hd__inv_2
X_11028_ _19954_/Q _16896_/A vssd1 vssd1 vccd1 vccd1 _16901_/A sky130_fd_sc_hd__or2_1
X_19673_ _19811_/CLK _19673_/D vssd1 vssd1 vccd1 vccd1 _19673_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_237_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16885_ _16894_/A _16885_/B vssd1 vssd1 vccd1 vccd1 _19026_/S sky130_fd_sc_hd__nor2_8
X_18624_ _18623_/X _16867_/Y _18667_/S vssd1 vssd1 vccd1 vccd1 _18624_/X sky130_fd_sc_hd__mux2_1
X_15836_ _15842_/A vssd1 vssd1 vccd1 vccd1 _15836_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_92_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_225_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_40_HCLK clkbuf_4_11_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _21182_/CLK sky130_fd_sc_hd__clkbuf_16
X_18555_ _18554_/X _12280_/Y _18910_/S vssd1 vssd1 vccd1 vccd1 _18555_/X sky130_fd_sc_hd__mux2_1
XFILLER_206_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15767_ _19642_/Q _15757_/X _15766_/X _15760_/X vssd1 vssd1 vccd1 vccd1 _19642_/D
+ sky130_fd_sc_hd__a22o_1
X_12979_ _17085_/A _12981_/A vssd1 vssd1 vccd1 vccd1 _12980_/S sky130_fd_sc_hd__or2_2
XFILLER_45_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17506_ _21217_/Q vssd1 vssd1 vccd1 vccd1 _17506_/Y sky130_fd_sc_hd__inv_2
XFILLER_233_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14718_ _14724_/A vssd1 vssd1 vccd1 vccd1 _14718_/X sky130_fd_sc_hd__buf_1
XANTENNA__12840__B1 _09628_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18486_ _18485_/X _14915_/Y _18907_/S vssd1 vssd1 vccd1 vccd1 _18486_/X sky130_fd_sc_hd__mux2_1
XFILLER_221_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15698_ _15698_/A vssd1 vssd1 vccd1 vccd1 _15698_/X sky130_fd_sc_hd__buf_1
XANTENNA__21180__RESET_B repeater216/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17437_ _19433_/Q vssd1 vssd1 vccd1 vccd1 _17437_/Y sky130_fd_sc_hd__inv_2
XFILLER_221_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14649_ _20179_/Q _14648_/Y _14642_/X _14570_/B vssd1 vssd1 vccd1 vccd1 _20179_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__18155__S _18775_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_221_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17368_ _17368_/A vssd1 vssd1 vccd1 vccd1 _17368_/X sky130_fd_sc_hd__buf_1
X_19107_ _19126_/S _14313_/Y _19125_/S vssd1 vssd1 vccd1 vccd1 _19107_/X sky130_fd_sc_hd__mux2_1
X_16319_ _16319_/A vssd1 vssd1 vccd1 vccd1 _16319_/X sky130_fd_sc_hd__buf_1
X_17299_ _20894_/Q vssd1 vssd1 vccd1 vccd1 _17299_/Y sky130_fd_sc_hd__inv_2
XFILLER_174_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19038_ _16838_/Y _20831_/Q _19046_/S vssd1 vssd1 vccd1 vccd1 _19938_/D sky130_fd_sc_hd__mux2_1
Xoutput101 _17406_/Y vssd1 vssd1 vccd1 vccd1 HRDATA[2] sky130_fd_sc_hd__clkbuf_2
XFILLER_115_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput112 _18109_/Y vssd1 vssd1 vccd1 vccd1 IRQ[0] sky130_fd_sc_hd__clkbuf_2
Xoutput123 _17078_/X vssd1 vssd1 vccd1 vccd1 IRQ[5] sky130_fd_sc_hd__clkbuf_2
XANTENNA__18087__A1 _18617_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput134 _17042_/Y vssd1 vssd1 vccd1 vccd1 SSn_S2 sky130_fd_sc_hd__clkbuf_2
Xoutput145 _21135_/Q vssd1 vssd1 vccd1 vccd1 sda_oen_o_S5 sky130_fd_sc_hd__clkbuf_2
XANTENNA__20409__RESET_B repeater185/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21000_ _21001_/CLK _21000_/D repeater190/X vssd1 vssd1 vccd1 vccd1 _21000_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_141_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12659__B1 _12658_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20062__RESET_B repeater281/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09624_ _09660_/A vssd1 vssd1 vccd1 vccd1 _09624_/X sky130_fd_sc_hd__buf_1
XFILLER_28_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11790__B hold9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13084__B1 _12855_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14159__A _20551_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12831__B1 _12663_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20715_ _21357_/CLK _20715_/D repeater254/X vssd1 vssd1 vccd1 vccd1 _20715_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19198__S0 _20130_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13387__A1 _20497_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20646_ _21486_/CLK _20646_/D repeater199/X vssd1 vssd1 vccd1 vccd1 _20646_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_211_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20577_ _20946_/CLK _20577_/D repeater258/X vssd1 vssd1 vccd1 vccd1 _20577_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_194_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10330_ _20726_/Q vssd1 vssd1 vccd1 vccd1 _10330_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10261_ _10261_/A _10418_/A vssd1 vssd1 vccd1 vccd1 _10262_/B sky130_fd_sc_hd__or2_2
XFILLER_11_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12000_ _20994_/Q _12000_/B vssd1 vssd1 vccd1 vccd1 _12001_/B sky130_fd_sc_hd__or2_1
XFILLER_127_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17825__A1 _18271_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10192_ _10153_/A _10153_/B _10185_/X _10190_/Y vssd1 vssd1 vccd1 vccd1 _21392_/D
+ sky130_fd_sc_hd__a211oi_4
XFILLER_239_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21129_ _21134_/CLK _21129_/D repeater192/X vssd1 vssd1 vccd1 vccd1 _21129_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_78_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_63_HCLK clkbuf_4_14_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _21341_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_247_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13951_ _20639_/Q vssd1 vssd1 vccd1 vccd1 _13951_/Y sky130_fd_sc_hd__inv_2
XFILLER_87_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12902_ _12934_/A vssd1 vssd1 vccd1 vccd1 _12936_/A sky130_fd_sc_hd__inv_2
X_16670_ _21158_/Q _11446_/B _11447_/B vssd1 vssd1 vccd1 vccd1 _16670_/X sky130_fd_sc_hd__a21bo_1
X_13882_ _13882_/A _14002_/A vssd1 vssd1 vccd1 vccd1 _13883_/B sky130_fd_sc_hd__or2_1
XFILLER_46_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12833_ _20763_/Q _12829_/X _12668_/X _12830_/X vssd1 vssd1 vccd1 vccd1 _20763_/D
+ sky130_fd_sc_hd__a22o_1
X_15621_ _19712_/Q _15618_/X _15483_/X _15619_/X vssd1 vssd1 vccd1 vccd1 _19712_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13075__B1 _12928_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_243_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18340_ _18032_/Y _20025_/Q _18669_/S vssd1 vssd1 vccd1 vccd1 _18340_/X sky130_fd_sc_hd__mux2_1
X_15552_ _19746_/Q _15543_/X _15514_/X _15546_/X vssd1 vssd1 vccd1 vccd1 _19746_/D
+ sky130_fd_sc_hd__a22o_1
X_12764_ _20801_/Q _12757_/X _12660_/X _12760_/X vssd1 vssd1 vccd1 vccd1 _20801_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16013__B1 _16012_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14503_ _14503_/A _14507_/A vssd1 vssd1 vccd1 vccd1 _14504_/B sky130_fd_sc_hd__or2_2
X_11715_ _11721_/A vssd1 vssd1 vccd1 vccd1 _11715_/X sky130_fd_sc_hd__buf_1
XPHY_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18271_ _18270_/X _21285_/Q _18880_/S vssd1 vssd1 vccd1 vccd1 _18271_/X sky130_fd_sc_hd__mux2_2
X_15483_ _15772_/A vssd1 vssd1 vccd1 vccd1 _15483_/X sky130_fd_sc_hd__buf_1
XFILLER_203_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12695_ _20822_/Q _12693_/X _09655_/X _12694_/X vssd1 vssd1 vccd1 vccd1 _20822_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19189__S0 _19280_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17222_ _17316_/A vssd1 vssd1 vccd1 vccd1 _17223_/A sky130_fd_sc_hd__buf_1
XPHY_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14434_ _14434_/A _14434_/B _14434_/C _14434_/D vssd1 vssd1 vccd1 vccd1 _14450_/C
+ sky130_fd_sc_hd__and4_1
X_11646_ _11646_/A vssd1 vssd1 vccd1 vccd1 _11646_/X sky130_fd_sc_hd__buf_1
XPHY_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput14 HADDR[21] vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__clkbuf_1
XPHY_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14365_ _14460_/C _14493_/A vssd1 vssd1 vccd1 vccd1 _14366_/B sky130_fd_sc_hd__or2_2
X_17153_ _17153_/A vssd1 vssd1 vccd1 vccd1 _17390_/A sky130_fd_sc_hd__buf_1
Xinput25 HADDR[31] vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__buf_1
XPHY_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11577_ _11577_/A vssd1 vssd1 vccd1 vccd1 _11577_/Y sky130_fd_sc_hd__inv_2
Xinput36 HTRANS[0] vssd1 vssd1 vccd1 vccd1 input36/X sky130_fd_sc_hd__buf_1
XPHY_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_repeater241_A repeater242/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18703__S _18930_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput47 HWDATA[18] vssd1 vssd1 vccd1 vccd1 input47/X sky130_fd_sc_hd__clkbuf_4
X_16104_ _19480_/Q _16101_/X _15879_/X _16102_/X vssd1 vssd1 vccd1 vccd1 _19480_/D
+ sky130_fd_sc_hd__a22o_1
Xinput58 HWDATA[28] vssd1 vssd1 vccd1 vccd1 input58/X sky130_fd_sc_hd__clkbuf_4
X_13316_ _13322_/A vssd1 vssd1 vccd1 vccd1 _13316_/X sky130_fd_sc_hd__buf_1
XFILLER_183_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10528_ _21342_/Q _10375_/X _10527_/Y vssd1 vssd1 vccd1 vccd1 _21342_/D sky130_fd_sc_hd__o21a_1
Xinput69 HWDATA[9] vssd1 vssd1 vccd1 vccd1 input69/X sky130_fd_sc_hd__buf_2
X_17084_ _17814_/A vssd1 vssd1 vccd1 vccd1 _18874_/S sky130_fd_sc_hd__buf_6
X_14296_ _20126_/Q vssd1 vssd1 vccd1 vccd1 _15574_/A sky130_fd_sc_hd__buf_1
XANTENNA__17827__B _17827_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12889__A0 _12809_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16035_ _16042_/A vssd1 vssd1 vccd1 vccd1 _16035_/X sky130_fd_sc_hd__buf_1
X_13247_ _20569_/Q _13239_/X _13163_/X _13241_/X vssd1 vssd1 vccd1 vccd1 _20569_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_171_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10459_ _20666_/Q vssd1 vssd1 vccd1 vccd1 _10459_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20502__RESET_B repeater257/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09626__A input51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13178_ _11973_/A _16525_/B _13177_/Y vssd1 vssd1 vccd1 vccd1 _13178_/X sky130_fd_sc_hd__a21o_1
X_12129_ _20961_/Q _12127_/Y _20976_/Q _12128_/Y vssd1 vssd1 vccd1 vccd1 _12129_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__13148__A input41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17986_ _18368_/X _17907_/X _18370_/X _17908_/X vssd1 vssd1 vccd1 vccd1 _17989_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19725_ _20327_/CLK _19725_/D vssd1 vssd1 vccd1 vccd1 _19725_/Q sky130_fd_sc_hd__dfxtp_1
X_16937_ _16937_/A vssd1 vssd1 vccd1 vccd1 _16937_/Y sky130_fd_sc_hd__inv_2
XFILLER_96_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12987__A _13013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16459__A _16459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10116__B2 _20795_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_237_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19656_ _19821_/CLK _19656_/D vssd1 vssd1 vccd1 vccd1 _19656_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17281__C _18910_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16868_ _16868_/A vssd1 vssd1 vccd1 vccd1 _16868_/Y sky130_fd_sc_hd__inv_2
XFILLER_237_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18607_ _17830_/X _10947_/Y _18928_/S vssd1 vssd1 vccd1 vccd1 _18607_/X sky130_fd_sc_hd__mux2_1
X_15819_ _15825_/A vssd1 vssd1 vccd1 vccd1 _15819_/X sky130_fd_sc_hd__clkbuf_2
X_19587_ _21218_/CLK _19587_/D vssd1 vssd1 vccd1 vccd1 _19587_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__21361__RESET_B repeater254/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16799_ _16820_/A _16799_/B vssd1 vssd1 vccd1 vccd1 _16799_/Y sky130_fd_sc_hd__nor2_1
XFILLER_240_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18538_ _18537_/X _20515_/Q _18910_/S vssd1 vssd1 vccd1 vccd1 _18538_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10300__A _20732_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18469_ _18468_/X _14578_/A _18898_/S vssd1 vssd1 vccd1 vccd1 _18469_/X sky130_fd_sc_hd__mux2_2
XFILLER_33_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20500_ _20929_/CLK _20500_/D repeater265/X vssd1 vssd1 vccd1 vccd1 _20500_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_20_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21480_ _21480_/CLK _21480_/D repeater206/X vssd1 vssd1 vccd1 vccd1 _21480_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_165_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12041__A1 _12036_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20431_ _21009_/CLK _20431_/D repeater235/X vssd1 vssd1 vccd1 vccd1 _20431_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_158_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18613__S _18666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11131__A _21005_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20362_ _20951_/CLK _20362_/D repeater272/X vssd1 vssd1 vccd1 vccd1 _20362_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_161_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14442__A _20029_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20293_ _20293_/CLK _20293_/D repeater263/X vssd1 vssd1 vccd1 vccd1 _20293_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_103_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_86_HCLK clkbuf_4_12_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _21349_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_115_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_229_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__21449__RESET_B repeater248/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16243__B1 _16012_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09607_ _20869_/Q vssd1 vssd1 vccd1 vccd1 _11187_/A sky130_fd_sc_hd__inv_2
XANTENNA__13057__B1 _12989_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__21031__RESET_B repeater242/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11500_ _19111_/X vssd1 vssd1 vccd1 vccd1 _11500_/Y sky130_fd_sc_hd__inv_2
XPHY_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12480_ _12480_/A vssd1 vssd1 vccd1 vccd1 _12480_/X sky130_fd_sc_hd__buf_1
XFILLER_185_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11431_ _11430_/Y _11408_/X _11413_/X _11390_/B _11414_/X vssd1 vssd1 vccd1 vccd1
+ _11432_/A sky130_fd_sc_hd__o32a_1
XPHY_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20629_ _20697_/CLK _20629_/D repeater193/X vssd1 vssd1 vccd1 vccd1 _20629_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17928__A _17928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18523__S _18787_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14150_ _20556_/Q _14095_/A _14146_/Y _20259_/Q _14149_/X vssd1 vssd1 vccd1 vccd1
+ _14155_/C sky130_fd_sc_hd__o221a_1
X_11362_ _11390_/A _11362_/B _11362_/C vssd1 vssd1 vccd1 vccd1 _11364_/A sky130_fd_sc_hd__or3_1
XFILLER_192_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13101_ _20636_/Q _13098_/X _12879_/X _13099_/X vssd1 vssd1 vccd1 vccd1 _20636_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_137_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10313_ _20714_/Q vssd1 vssd1 vccd1 vccd1 _10313_/Y sky130_fd_sc_hd__inv_2
XFILLER_153_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14081_ _14081_/A _14081_/B vssd1 vssd1 vccd1 vccd1 _14209_/A sky130_fd_sc_hd__or2_1
X_11293_ _20901_/Q vssd1 vssd1 vccd1 vccd1 _11307_/C sky130_fd_sc_hd__buf_1
XFILLER_4_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13032_ _13313_/A vssd1 vssd1 vccd1 vccd1 _13032_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_180_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input52_A HWDATA[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10244_ _21359_/Q vssd1 vssd1 vccd1 vccd1 _10274_/A sky130_fd_sc_hd__inv_2
XFILLER_121_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17840_ _17928_/A vssd1 vssd1 vccd1 vccd1 _17840_/X sky130_fd_sc_hd__buf_1
X_10175_ _10175_/A vssd1 vssd1 vccd1 vccd1 _10175_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17771_ _19461_/Q vssd1 vssd1 vccd1 vccd1 _17771_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12099__B2 _17806_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14983_ _14960_/B _14874_/B _14981_/Y _14975_/X vssd1 vssd1 vccd1 vccd1 _20096_/D
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__13296__B1 _13219_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_219_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19510_ _19784_/CLK _19510_/D vssd1 vssd1 vccd1 vccd1 _19510_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16722_ _20984_/Q _20983_/Q _11991_/B vssd1 vssd1 vccd1 vccd1 _16722_/X sky130_fd_sc_hd__a21bo_1
X_13934_ _13931_/Y _20317_/Q _13932_/Y _20311_/Q _13933_/X vssd1 vssd1 vccd1 vccd1
+ _13947_/A sky130_fd_sc_hd__o221a_1
XFILLER_219_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16234__B1 _16231_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19441_ _20137_/CLK _19441_/D vssd1 vssd1 vccd1 vccd1 _19441_/Q sky130_fd_sc_hd__dfxtp_1
X_16653_ _19861_/Q _15295_/B _15296_/B vssd1 vssd1 vccd1 vccd1 _16653_/X sky130_fd_sc_hd__a21bo_1
XANTENNA_repeater191_A repeater212/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13865_ _13865_/A _13865_/B _14031_/C vssd1 vssd1 vccd1 vccd1 _14010_/C sky130_fd_sc_hd__or3_1
X_15604_ _15604_/A vssd1 vssd1 vccd1 vccd1 _15604_/X sky130_fd_sc_hd__buf_1
XFILLER_90_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19372_ _19777_/CLK _19372_/D vssd1 vssd1 vccd1 vccd1 _19372_/Q sky130_fd_sc_hd__dfxtp_1
X_12816_ _12809_/X _20770_/Q _12816_/S vssd1 vssd1 vccd1 vccd1 _20770_/D sky130_fd_sc_hd__mux2_1
X_16584_ _19991_/Q _16584_/B vssd1 vssd1 vccd1 vccd1 _16585_/C sky130_fd_sc_hd__nand2_1
X_13796_ _20611_/Q vssd1 vssd1 vccd1 vccd1 _13796_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18323_ _18322_/X _16983_/Y _18680_/S vssd1 vssd1 vccd1 vccd1 _18323_/X sky130_fd_sc_hd__mux2_1
XFILLER_187_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15535_ _19754_/Q _15529_/X _15514_/X _15531_/X vssd1 vssd1 vccd1 vccd1 _19754_/D
+ sky130_fd_sc_hd__a22o_1
X_12747_ _20807_/Q _12745_/X _12746_/X vssd1 vssd1 vccd1 vccd1 _20807_/D sky130_fd_sc_hd__a21bo_1
XANTENNA__14527__A _17169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18254_ _18253_/X _10634_/Y _18891_/S vssd1 vssd1 vccd1 vccd1 _18254_/X sky130_fd_sc_hd__mux2_1
XFILLER_147_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12678_ _20831_/Q _12672_/X _09628_/X _12674_/X vssd1 vssd1 vccd1 vccd1 _20831_/D
+ sky130_fd_sc_hd__a22o_1
X_15466_ _15609_/A _15466_/B _16616_/B vssd1 vssd1 vccd1 vccd1 _16297_/C sky130_fd_sc_hd__or3_4
XFILLER_187_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17205_ _18021_/A vssd1 vssd1 vccd1 vccd1 _17205_/X sky130_fd_sc_hd__buf_2
X_14417_ _21486_/Q vssd1 vssd1 vccd1 vccd1 _14417_/Y sky130_fd_sc_hd__inv_2
X_11629_ _21107_/Q _11628_/Y _11623_/B vssd1 vssd1 vccd1 vccd1 _21107_/D sky130_fd_sc_hd__o21a_1
XFILLER_8_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13220__B1 _13219_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17838__A _17838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18185_ _18184_/X _20267_/Q _18904_/S vssd1 vssd1 vccd1 vccd1 _18185_/X sky130_fd_sc_hd__mux2_1
XANTENNA__18433__S _18907_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15397_ _15397_/A _15655_/B _16311_/C vssd1 vssd1 vccd1 vccd1 _15405_/A sky130_fd_sc_hd__or3_4
XPHY_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17136_ _17136_/A vssd1 vssd1 vccd1 vccd1 _17175_/B sky130_fd_sc_hd__buf_2
X_14348_ _20212_/Q vssd1 vssd1 vccd1 vccd1 _14351_/A sky130_fd_sc_hd__inv_2
XFILLER_144_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17067_ _20255_/Q _20253_/Q vssd1 vssd1 vccd1 vccd1 _17067_/X sky130_fd_sc_hd__or2_1
X_14279_ _14279_/A _14288_/A vssd1 vssd1 vccd1 vccd1 _14283_/B sky130_fd_sc_hd__nor2_1
XANTENNA__14262__A _14262_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14720__B1 _14262_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16018_ _16465_/A vssd1 vssd1 vccd1 vccd1 _16297_/A sky130_fd_sc_hd__buf_1
XFILLER_143_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19813__CLK _19813_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18462__A1 _10584_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17969_ _18191_/X _17928_/X _18197_/X _17960_/X vssd1 vssd1 vccd1 vccd1 _17969_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_214_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_109_HCLK_A clkbuf_opt_3_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_226_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19708_ _19777_/CLK _19708_/D vssd1 vssd1 vccd1 vccd1 _19708_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_214_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20980_ _20980_/CLK _20980_/D repeater272/X vssd1 vssd1 vccd1 vccd1 _20980_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_65_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19937__RESET_B repeater251/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19639_ _20326_/CLK _19639_/D vssd1 vssd1 vccd1 vccd1 _19639_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13039__B1 _12872_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18608__S _18908_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_214_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21463_ _21481_/CLK _21463_/D repeater205/X vssd1 vssd1 vccd1 vccd1 _21463_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18343__S _18906_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20414_ _20957_/CLK _20414_/D repeater186/X vssd1 vssd1 vccd1 vccd1 _20414_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_119_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18150__A0 _17281_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21394_ _21401_/CLK _21394_/D repeater253/X vssd1 vssd1 vccd1 vccd1 _21394_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_175_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20345_ _20428_/CLK _20345_/D repeater269/X vssd1 vssd1 vccd1 vccd1 _20345_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_135_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20276_ _20286_/CLK _20276_/D repeater262/X vssd1 vssd1 vccd1 vccd1 _20276_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_191_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18453__A1 _10592_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21283__RESET_B repeater211/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11980_ _11978_/A _11972_/A _11978_/Y vssd1 vssd1 vccd1 vccd1 _21000_/D sky130_fd_sc_hd__a21oi_1
XFILLER_84_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10859__B _10859_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_244_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10931_ _10931_/A _10931_/B _10931_/C _10931_/D vssd1 vssd1 vccd1 vccd1 _10931_/X
+ sky130_fd_sc_hd__or4_1
XANTENNA__18518__S _18902_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13650_ _20368_/Q _13645_/X _13442_/X _13646_/X vssd1 vssd1 vccd1 vccd1 _20368_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_44_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10862_ _09931_/X _21268_/Q _10862_/S vssd1 vssd1 vccd1 vccd1 _21268_/D sky130_fd_sc_hd__mux2_1
XFILLER_232_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12601_ _12601_/A vssd1 vssd1 vccd1 vccd1 _12601_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_169_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13581_ _13595_/A vssd1 vssd1 vccd1 vccd1 _13581_/X sky130_fd_sc_hd__buf_1
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10793_ _10793_/A vssd1 vssd1 vccd1 vccd1 _10793_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13450__B1 _13449_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12532_ _12524_/X _12525_/Y _19987_/Q _20910_/Q _12518_/X vssd1 vssd1 vccd1 vccd1
+ _20910_/D sky130_fd_sc_hd__a32o_1
XFILLER_185_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15320_ _20242_/Q _15320_/B vssd1 vssd1 vccd1 vccd1 _15320_/Y sky130_fd_sc_hd__nor2_1
XFILLER_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15251_ _20496_/Q vssd1 vssd1 vccd1 vccd1 _15251_/Y sky130_fd_sc_hd__inv_2
X_12463_ _20933_/Q _12461_/Y _12480_/A _12423_/B vssd1 vssd1 vccd1 vccd1 _20933_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__18253__S _18896_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13202__B1 _12996_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11414_ _11418_/A vssd1 vssd1 vccd1 vccd1 _11414_/X sky130_fd_sc_hd__buf_1
X_14202_ _20276_/Q _14201_/Y _14087_/B _14191_/X vssd1 vssd1 vccd1 vccd1 _20276_/D
+ sky130_fd_sc_hd__o211a_1
X_15182_ _20065_/Q _15181_/Y _15166_/X _15080_/B vssd1 vssd1 vccd1 vccd1 _20065_/D
+ sky130_fd_sc_hd__o211a_1
X_12394_ _12469_/B vssd1 vssd1 vccd1 vccd1 _12490_/B sky130_fd_sc_hd__buf_1
XFILLER_165_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14133_ _20548_/Q vssd1 vssd1 vccd1 vccd1 _14133_/Y sky130_fd_sc_hd__inv_2
X_11345_ _21181_/Q _21180_/Q _11783_/C vssd1 vssd1 vccd1 vccd1 _11348_/C sky130_fd_sc_hd__or3_1
X_19990_ _21196_/CLK _19990_/D repeater217/X vssd1 vssd1 vccd1 vccd1 _19990_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_99_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18941_ _16701_/X _20900_/Q _18946_/S vssd1 vssd1 vccd1 vccd1 _18941_/X sky130_fd_sc_hd__mux2_1
X_14064_ _20264_/Q vssd1 vssd1 vccd1 vccd1 _14075_/A sky130_fd_sc_hd__inv_2
X_11276_ _20917_/Q vssd1 vssd1 vccd1 vccd1 _11304_/D sky130_fd_sc_hd__inv_2
XFILLER_125_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13015_ _20684_/Q _13012_/X _12928_/X _13013_/X vssd1 vssd1 vccd1 vccd1 _20684_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_79_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10227_ _10227_/A _10227_/B _10227_/C vssd1 vssd1 vccd1 vccd1 _21377_/D sky130_fd_sc_hd__nor3_1
X_18872_ _18871_/X _11024_/Y _18910_/S vssd1 vssd1 vccd1 vccd1 _18872_/X sky130_fd_sc_hd__mux2_1
XFILLER_121_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater204_A repeater205/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16455__B1 _11486_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17823_ _17823_/A vssd1 vssd1 vccd1 vccd1 _17954_/A sky130_fd_sc_hd__clkbuf_2
X_10158_ _10158_/A _10182_/A vssd1 vssd1 vccd1 vccd1 _10159_/B sky130_fd_sc_hd__or2_2
XANTENNA__13269__B1 _13265_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18001__B _18001_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13426__A input41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17754_ _19605_/Q _17773_/B vssd1 vssd1 vccd1 vccd1 _17754_/X sky130_fd_sc_hd__or2_1
XFILLER_236_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14966_ _14881_/B _14880_/A _14965_/X _14881_/A vssd1 vssd1 vccd1 vccd1 _14967_/C
+ sky130_fd_sc_hd__o31a_1
X_10089_ _20773_/Q vssd1 vssd1 vccd1 vccd1 _10089_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16705_ _16709_/A _18940_/X vssd1 vssd1 vccd1 vccd1 _19896_/D sky130_fd_sc_hd__and2_1
X_13917_ _20653_/Q vssd1 vssd1 vccd1 vccd1 _13917_/Y sky130_fd_sc_hd__inv_2
XFILLER_47_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17685_ _18707_/X _17775_/B vssd1 vssd1 vccd1 vccd1 _17685_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__18428__S _18680_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14897_ _20566_/Q vssd1 vssd1 vccd1 vccd1 _14897_/Y sky130_fd_sc_hd__inv_2
X_19424_ _19521_/CLK _19424_/D vssd1 vssd1 vccd1 vccd1 _19424_/Q sky130_fd_sc_hd__dfxtp_1
X_16636_ _16663_/A vssd1 vssd1 vccd1 vccd1 _16643_/A sky130_fd_sc_hd__buf_1
XFILLER_90_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13848_ _13848_/A vssd1 vssd1 vccd1 vccd1 _13974_/B sky130_fd_sc_hd__buf_1
XFILLER_222_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19355_ _21453_/CLK _19355_/D vssd1 vssd1 vccd1 vccd1 _19355_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16567_ _16744_/A _16738_/B _16556_/B _16566_/X vssd1 vssd1 vccd1 vccd1 _19996_/D
+ sky130_fd_sc_hd__o31ai_1
XFILLER_50_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_188_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13779_ _20599_/Q _14566_/A _13775_/Y _20195_/Q _13778_/X vssd1 vssd1 vccd1 vccd1
+ _13786_/C sky130_fd_sc_hd__o221a_1
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18306_ _18848_/A0 _10352_/Y _18884_/S vssd1 vssd1 vccd1 vccd1 _18306_/X sky130_fd_sc_hd__mux2_1
X_15518_ _15788_/A vssd1 vssd1 vccd1 vccd1 _15518_/X sky130_fd_sc_hd__buf_1
XFILLER_200_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19286_ _19282_/X _19283_/X _19284_/X _19285_/X _21018_/Q _21019_/Q vssd1 vssd1 vccd1
+ vccd1 _19286_/X sky130_fd_sc_hd__mux4_2
X_16498_ _16498_/A _16502_/A vssd1 vssd1 vccd1 vccd1 _16498_/Y sky130_fd_sc_hd__nor2_4
XFILLER_149_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18237_ _20861_/Q input10/X _18242_/S vssd1 vssd1 vccd1 vccd1 _18237_/X sky130_fd_sc_hd__mux2_1
X_15449_ _15459_/A vssd1 vssd1 vccd1 vccd1 _15449_/X sky130_fd_sc_hd__buf_1
XANTENNA__18163__S _18902_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18168_ _18167_/X _10422_/Y _18617_/S vssd1 vssd1 vccd1 vccd1 _18168_/X sky130_fd_sc_hd__mux2_1
XFILLER_190_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17119_ _19606_/Q vssd1 vssd1 vccd1 vccd1 _17119_/Y sky130_fd_sc_hd__inv_2
X_18099_ _20842_/Q vssd1 vssd1 vccd1 vccd1 _18099_/Y sky130_fd_sc_hd__inv_2
X_20130_ _21235_/CLK _20130_/D repeater249/X vssd1 vssd1 vccd1 vccd1 _20130_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_116_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09941_ _11488_/B vssd1 vssd1 vccd1 vccd1 _17133_/A sky130_fd_sc_hd__clkbuf_2
X_20061_ _20066_/CLK _20061_/D repeater281/X vssd1 vssd1 vccd1 vccd1 _20061_/Q sky130_fd_sc_hd__dfrtp_1
X_09872_ _09872_/A vssd1 vssd1 vccd1 vccd1 _09878_/B sky130_fd_sc_hd__buf_1
XFILLER_140_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09814__A _09827_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater220 repeater223/X vssd1 vssd1 vccd1 vccd1 repeater220/X sky130_fd_sc_hd__buf_8
Xrepeater231 repeater234/X vssd1 vssd1 vccd1 vccd1 repeater231/X sky130_fd_sc_hd__buf_8
Xrepeater242 repeater250/X vssd1 vssd1 vccd1 vccd1 repeater242/X sky130_fd_sc_hd__buf_8
Xrepeater253 repeater255/X vssd1 vssd1 vccd1 vccd1 repeater253/X sky130_fd_sc_hd__buf_4
Xrepeater264 repeater265/X vssd1 vssd1 vccd1 vccd1 repeater264/X sky130_fd_sc_hd__buf_8
XPHY_4407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_116_HCLK clkbuf_opt_3_HCLK/A vssd1 vssd1 vccd1 vccd1 _20937_/CLK sky130_fd_sc_hd__clkbuf_16
Xrepeater275 repeater277/X vssd1 vssd1 vccd1 vccd1 repeater275/X sky130_fd_sc_hd__clkbuf_8
XPHY_4418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20963_ _20981_/CLK _20963_/D repeater185/X vssd1 vssd1 vccd1 vccd1 _20963_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_4429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18338__S _18898_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_241_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_226_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20894_ _21141_/CLK _20894_/D repeater192/X vssd1 vssd1 vccd1 vccd1 _20894_/Q sky130_fd_sc_hd__dfstp_1
XPHY_3739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20676__RESET_B repeater208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_241_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21446_ _21449_/CLK _21446_/D repeater248/X vssd1 vssd1 vccd1 vccd1 _21446_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_119_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20836__CLK _20930_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21377_ _21379_/CLK _21377_/D repeater213/X vssd1 vssd1 vccd1 vccd1 _21377_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18801__S _18835_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11130_ _21222_/Q vssd1 vssd1 vccd1 vccd1 _15756_/A sky130_fd_sc_hd__buf_1
XFILLER_122_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20328_ _20331_/CLK _20328_/D repeater190/X vssd1 vssd1 vccd1 vccd1 _20328_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_162_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11061_ _11061_/A _11074_/A vssd1 vssd1 vccd1 vccd1 _11071_/A sky130_fd_sc_hd__or2_1
XFILLER_122_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20259_ _20661_/CLK _20259_/D repeater262/X vssd1 vssd1 vccd1 vccd1 _20259_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_150_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10012_ _17032_/A _10000_/X _20018_/Q _20019_/Q vssd1 vssd1 vccd1 vccd1 _10013_/B
+ sky130_fd_sc_hd__a31oi_1
XANTENNA__16437__B1 _11486_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19859__RESET_B repeater226/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14820_ _20111_/Q _20112_/Q _14823_/S vssd1 vssd1 vccd1 vccd1 _20112_/D sky130_fd_sc_hd__mux2_1
XFILLER_218_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input15_A HADDR[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14751_ _14751_/A _14751_/B vssd1 vssd1 vccd1 vccd1 _14757_/A sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_155_HCLK_A clkbuf_opt_1_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11963_ _20598_/Q vssd1 vssd1 vccd1 vccd1 _11973_/A sky130_fd_sc_hd__buf_1
XANTENNA__13671__B1 _13555_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13702_ _20338_/Q _13699_/X _13509_/X _13700_/X vssd1 vssd1 vccd1 vccd1 _20338_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_244_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17470_ _17462_/Y _17286_/X _17463_/Y _17147_/X _17469_/X vssd1 vssd1 vccd1 vccd1
+ _17470_/X sky130_fd_sc_hd__o221a_2
X_10914_ _20170_/Q vssd1 vssd1 vccd1 vccd1 _10917_/A sky130_fd_sc_hd__inv_2
XFILLER_189_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11894_ _11881_/A _11889_/X _11881_/A _11889_/X vssd1 vssd1 vccd1 vccd1 _21020_/D
+ sky130_fd_sc_hd__o2bb2a_1
X_14682_ _14682_/A vssd1 vssd1 vccd1 vccd1 _14682_/Y sky130_fd_sc_hd__inv_2
XFILLER_204_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16421_ _16427_/A vssd1 vssd1 vccd1 vccd1 _16428_/A sky130_fd_sc_hd__inv_2
X_13633_ _13633_/A vssd1 vssd1 vccd1 vccd1 _13652_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_32_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10845_ _10853_/A vssd1 vssd1 vccd1 vccd1 _10849_/A sky130_fd_sc_hd__inv_2
XFILLER_204_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13423__B1 _13422_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19140_ _19656_/Q _19648_/Q _19632_/Q _19816_/Q _19285_/S0 _21017_/Q vssd1 vssd1
+ vccd1 vccd1 _19140_/X sky130_fd_sc_hd__mux4_2
X_16352_ _16352_/A vssd1 vssd1 vccd1 vccd1 _16352_/X sky130_fd_sc_hd__buf_1
X_10776_ _10776_/A _10801_/A vssd1 vssd1 vccd1 vccd1 _10777_/B sky130_fd_sc_hd__or2_2
XANTENNA__18362__A0 _17281_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13564_ _20418_/Q _13559_/X _13477_/X _13561_/X vssd1 vssd1 vccd1 vccd1 _20418_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_158_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15303_ _20042_/Q _15302_/X _20041_/Q _18962_/S vssd1 vssd1 vccd1 vccd1 _20042_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_185_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12515_ _12515_/A _12520_/A vssd1 vssd1 vccd1 vccd1 _12528_/A sky130_fd_sc_hd__or2_2
X_19071_ _16732_/X _21139_/Q _19908_/D vssd1 vssd1 vccd1 vccd1 _19071_/X sky130_fd_sc_hd__mux2_1
XANTENNA__19079__S _19908_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13495_ _20448_/Q _13492_/X _13418_/X _13494_/X vssd1 vssd1 vccd1 vccd1 _20448_/D
+ sky130_fd_sc_hd__a22o_1
X_16283_ _20329_/Q vssd1 vssd1 vccd1 vccd1 _16283_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_repeater154_A _18617_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18022_ _18311_/X _18021_/X _18287_/X _17960_/X vssd1 vssd1 vccd1 vccd1 _18022_/X
+ sky130_fd_sc_hd__o22a_2
X_15234_ _20466_/Q vssd1 vssd1 vccd1 vccd1 _15234_/Y sky130_fd_sc_hd__inv_2
X_12446_ _12431_/A _12431_/B _12445_/X _12443_/Y vssd1 vssd1 vccd1 vccd1 _20942_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_8_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09618__B _13046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12377_ _12377_/A vssd1 vssd1 vccd1 vccd1 _12377_/Y sky130_fd_sc_hd__inv_2
X_15165_ _15165_/A vssd1 vssd1 vccd1 vccd1 _15165_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18711__S _18879_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11328_ _21184_/Q vssd1 vssd1 vccd1 vccd1 _11390_/A sky130_fd_sc_hd__buf_1
XANTENNA_output83_A _17892_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14116_ _20537_/Q vssd1 vssd1 vccd1 vccd1 _14116_/Y sky130_fd_sc_hd__inv_2
XFILLER_180_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15096_ _20451_/Q vssd1 vssd1 vccd1 vccd1 _15096_/Y sky130_fd_sc_hd__inv_2
X_19973_ _20408_/CLK _19973_/D repeater184/X vssd1 vssd1 vccd1 vccd1 _19973_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_140_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18924_ _18923_/X _14313_/Y _18929_/S vssd1 vssd1 vccd1 vccd1 _18924_/X sky130_fd_sc_hd__mux2_1
X_11259_ _11543_/A vssd1 vssd1 vccd1 vccd1 _12506_/A sky130_fd_sc_hd__buf_1
X_14047_ _20281_/Q vssd1 vssd1 vccd1 vccd1 _14091_/A sky130_fd_sc_hd__inv_2
XFILLER_140_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_139_HCLK clkbuf_4_3_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _21401_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__19090__A1 _21056_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18855_ _18854_/X _12147_/Y _18909_/S vssd1 vssd1 vccd1 vccd1 _18855_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17806_ _17806_/A _17807_/B vssd1 vssd1 vccd1 vccd1 _17806_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__15100__B1 _20447_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18786_ _17079_/Y _12061_/Y _18908_/S vssd1 vssd1 vccd1 vccd1 _18786_/X sky130_fd_sc_hd__mux2_1
X_15998_ _19534_/Q _15993_/X _15951_/X _15994_/X vssd1 vssd1 vccd1 vccd1 _19534_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_243_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17737_ _17548_/X _17719_/X _17560_/X _17728_/X _17736_/X vssd1 vssd1 vccd1 vccd1
+ _17737_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_47_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14949_ _14901_/X _14949_/B _14949_/C _14949_/D vssd1 vssd1 vccd1 vccd1 _14950_/A
+ sky130_fd_sc_hd__and4b_1
XANTENNA__12995__A _13012_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16467__A _16473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18158__S _18617_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17668_ _19700_/Q vssd1 vssd1 vccd1 vccd1 _17668_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_14_HCLK_A clkbuf_opt_2_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19407_ _19813_/CLK _19407_/D vssd1 vssd1 vccd1 vccd1 _19407_/Q sky130_fd_sc_hd__dfxtp_1
X_16619_ _16619_/A _16619_/B vssd1 vssd1 vccd1 vccd1 _16619_/Y sky130_fd_sc_hd__nor2_1
XFILLER_196_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_77_HCLK_A clkbuf_4_13_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17599_ _19723_/Q vssd1 vssd1 vccd1 vccd1 _17599_/Y sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_2_HCLK_A clkbuf_opt_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19338_ _20172_/CLK _19338_/D vssd1 vssd1 vccd1 vccd1 _19338_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19269_ _17122_/Y _17123_/Y _17124_/Y _17125_/Y _20130_/Q _20131_/Q vssd1 vssd1 vccd1
+ vccd1 _19269_/X sky130_fd_sc_hd__mux4_1
X_21300_ _21302_/CLK _21300_/D repeater209/X vssd1 vssd1 vccd1 vccd1 _21300_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_136_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21231_ _21239_/CLK _21231_/D repeater249/X vssd1 vssd1 vccd1 vccd1 _21231_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18621__S _18897_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21162_ _21162_/CLK _21162_/D repeater226/X vssd1 vssd1 vccd1 vccd1 _21162_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_160_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20113_ _21419_/CLK _20113_/D repeater234/X vssd1 vssd1 vccd1 vccd1 _20113_/Q sky130_fd_sc_hd__dfrtp_1
X_09924_ _21434_/Q _21435_/Q _09924_/S vssd1 vssd1 vccd1 vccd1 _21435_/D sky130_fd_sc_hd__mux2_1
X_21093_ _21164_/CLK _21093_/D repeater226/X vssd1 vssd1 vccd1 vccd1 _21093_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_59_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20044_ _20075_/CLK _20044_/D repeater276/X vssd1 vssd1 vccd1 vccd1 _20044_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__19952__RESET_B repeater270/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09855_ _09851_/X _09852_/Y _09853_/X _09857_/A _21445_/Q vssd1 vssd1 vccd1 vccd1
+ _09855_/X sky130_fd_sc_hd__a41o_1
XANTENNA_input7_A HADDR[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13066__A _13072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09786_ _14530_/C vssd1 vssd1 vccd1 vccd1 _18976_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__20857__RESET_B repeater243/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13653__B1 _13446_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20946_ _20946_/CLK _20946_/D repeater275/X vssd1 vssd1 vccd1 vccd1 _20946_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_4259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20877_ _21459_/CLK _20877_/D repeater244/X vssd1 vssd1 vccd1 vccd1 _20877_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_41_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10630_ _20767_/Q vssd1 vssd1 vccd1 vccd1 _10630_/Y sky130_fd_sc_hd__inv_2
XPHY_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19838__D _19838_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10561_ _21328_/Q vssd1 vssd1 vccd1 vccd1 _10657_/A sky130_fd_sc_hd__inv_2
XFILLER_22_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12300_ _12476_/A _20508_/Q _20945_/Q _12296_/Y _12299_/X vssd1 vssd1 vccd1 vccd1
+ _12301_/D sky130_fd_sc_hd__o221a_1
XFILLER_167_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13280_ input56/X vssd1 vssd1 vccd1 vccd1 _13280_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_212_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10492_ _20688_/Q vssd1 vssd1 vccd1 vccd1 _18005_/A sky130_fd_sc_hd__inv_2
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12231_ _12419_/A _20510_/Q _12424_/A _20515_/Q _12230_/X vssd1 vssd1 vccd1 vccd1
+ _12232_/D sky130_fd_sc_hd__o221a_1
XFILLER_170_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21429_ _21429_/CLK _21429_/D repeater229/X vssd1 vssd1 vccd1 vccd1 _21429_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_108_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18531__S _18850_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12392__B1 _12359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12162_ _20969_/Q _20351_/Q _12322_/A _12161_/Y vssd1 vssd1 vccd1 vccd1 _12162_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_2_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11113_ _11113_/A vssd1 vssd1 vccd1 vccd1 _11113_/X sky130_fd_sc_hd__buf_1
XANTENNA__15456__A _15663_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16970_ _16970_/A vssd1 vssd1 vccd1 vccd1 _16970_/Y sky130_fd_sc_hd__inv_2
X_12093_ _12315_/A vssd1 vssd1 vccd1 vccd1 _12093_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_49_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11044_ _16885_/B vssd1 vssd1 vccd1 vccd1 _11045_/B sky130_fd_sc_hd__inv_2
X_15921_ _15927_/A vssd1 vssd1 vccd1 vccd1 _15928_/A sky130_fd_sc_hd__inv_2
XANTENNA__19072__A1 _21138_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_237_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18640_ _17079_/Y _15277_/Y _18908_/S vssd1 vssd1 vccd1 vccd1 _18640_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15852_ _19605_/Q _15849_/X _15725_/X _15851_/X vssd1 vssd1 vccd1 vccd1 _19605_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_77_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20598__RESET_B repeater235/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_225_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14803_ _14803_/A _14803_/B vssd1 vssd1 vccd1 vccd1 _14804_/A sky130_fd_sc_hd__nand2_1
XFILLER_76_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18571_ _18848_/A0 _17866_/Y _18666_/S vssd1 vssd1 vccd1 vccd1 _18571_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13644__B1 _13586_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15783_ _19636_/Q _15779_/X _15730_/X _15781_/X vssd1 vssd1 vccd1 vccd1 _19636_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_output121_A _18114_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12995_ _13012_/A vssd1 vssd1 vccd1 vccd1 _12995_/X sky130_fd_sc_hd__buf_1
X_17522_ _19442_/Q vssd1 vssd1 vccd1 vccd1 _17522_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13704__A _15421_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14734_ _20143_/Q _14731_/X _13704_/X _14733_/X vssd1 vssd1 vccd1 vccd1 _20143_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_233_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11946_ _11946_/A vssd1 vssd1 vccd1 vccd1 _21009_/D sky130_fd_sc_hd__inv_2
XFILLER_55_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17453_ _21075_/Q vssd1 vssd1 vccd1 vccd1 _17453_/Y sky130_fd_sc_hd__inv_2
X_14665_ _20174_/Q _14663_/A _20174_/Q _14663_/A vssd1 vssd1 vccd1 vccd1 _14665_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_221_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20180__RESET_B repeater200/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18706__S _18930_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11877_ _11877_/A vssd1 vssd1 vccd1 vccd1 _11889_/B sky130_fd_sc_hd__inv_2
XFILLER_220_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16404_ _19333_/Q _16399_/X _16342_/X _16400_/X vssd1 vssd1 vccd1 vccd1 _19333_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_60_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13616_ _20390_/Q _13613_/X _13553_/X _13614_/X vssd1 vssd1 vccd1 vccd1 _20390_/D
+ sky130_fd_sc_hd__a22o_1
X_17384_ _16633_/Y _17286_/X _17375_/Y _17376_/X _17383_/X vssd1 vssd1 vccd1 vccd1
+ _17384_/X sky130_fd_sc_hd__o221a_2
X_10828_ _10762_/A _10762_/B _10827_/X _10825_/Y vssd1 vssd1 vccd1 vccd1 _21285_/D
+ sky130_fd_sc_hd__a211oi_2
X_14596_ _14596_/A vssd1 vssd1 vccd1 vccd1 _14596_/Y sky130_fd_sc_hd__inv_2
XFILLER_186_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19123_ _16484_/Y _16483_/Y _19123_/S vssd1 vssd1 vccd1 vccd1 _19123_/X sky130_fd_sc_hd__mux2_2
X_16335_ _16335_/A vssd1 vssd1 vccd1 vccd1 _16335_/X sky130_fd_sc_hd__buf_1
X_13547_ input58/X vssd1 vssd1 vccd1 vccd1 _13547_/X sky130_fd_sc_hd__clkbuf_4
X_10759_ _10759_/A _10833_/A vssd1 vssd1 vccd1 vccd1 _10760_/B sky130_fd_sc_hd__or2_1
XFILLER_40_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14535__A _20132_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19054_ _16767_/X _20815_/Q _19058_/S vssd1 vssd1 vccd1 vccd1 _19922_/D sky130_fd_sc_hd__mux2_1
X_16266_ _19404_/Q _16262_/X _16113_/X _16264_/X vssd1 vssd1 vccd1 vccd1 _19404_/D
+ sky130_fd_sc_hd__a22o_1
X_13478_ _20454_/Q _13472_/X _13477_/X _13473_/X vssd1 vssd1 vccd1 vccd1 _20454_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__21386__RESET_B repeater252/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18005_ _18005_/A _18006_/B vssd1 vssd1 vccd1 vccd1 _18005_/Y sky130_fd_sc_hd__nor2_1
X_15217_ _20494_/Q vssd1 vssd1 vccd1 vccd1 _18078_/A sky130_fd_sc_hd__inv_2
X_12429_ _12429_/A _12429_/B vssd1 vssd1 vccd1 vccd1 _12447_/A sky130_fd_sc_hd__or2_1
X_16197_ _16206_/A vssd1 vssd1 vccd1 vccd1 _16208_/A sky130_fd_sc_hd__inv_2
XANTENNA__18441__S _18910_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15148_ _20454_/Q vssd1 vssd1 vccd1 vccd1 _15148_/Y sky130_fd_sc_hd__inv_2
XFILLER_114_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19956_ _21234_/CLK _19956_/D repeater188/X vssd1 vssd1 vccd1 vccd1 _19956_/Q sky130_fd_sc_hd__dfrtp_1
X_15079_ _15079_/A _15181_/A vssd1 vssd1 vccd1 vccd1 _15080_/B sky130_fd_sc_hd__or2_1
XANTENNA__19554__CLK _19706_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18907_ _18906_/X _14914_/Y _18907_/S vssd1 vssd1 vccd1 vccd1 _18907_/X sky130_fd_sc_hd__mux2_2
X_19887_ _20915_/CLK _19887_/D repeater217/X vssd1 vssd1 vccd1 vccd1 _19889_/D sky130_fd_sc_hd__dfstp_1
XFILLER_206_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09640_ input44/X vssd1 vssd1 vccd1 vccd1 _12849_/A sky130_fd_sc_hd__buf_4
X_18838_ _18837_/X _16753_/A _18880_/S vssd1 vssd1 vccd1 vccd1 _18838_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18769_ _18845_/A0 _17451_/Y _18879_/S vssd1 vssd1 vccd1 vccd1 _18769_/X sky130_fd_sc_hd__mux2_1
XFILLER_222_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13635__B1 _13418_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20268__RESET_B repeater263/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20800_ _21405_/CLK _20800_/D repeater255/X vssd1 vssd1 vccd1 vccd1 _20800_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_236_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13614__A _13626_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18023__C1 _18022_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18574__A0 _18848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20731_ _21375_/CLK _20731_/D repeater257/X vssd1 vssd1 vccd1 vccd1 _20731_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__15388__B1 _15343_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18616__S _18891_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18326__A0 _18325_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20662_ _20665_/CLK _20662_/D repeater261/X vssd1 vssd1 vccd1 vccd1 _20662_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10973__A _20888_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20593_ _20665_/CLK _20593_/D repeater259/X vssd1 vssd1 vccd1 vccd1 _20593_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_191_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18351__S _18667_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21214_ _21223_/CLK _21214_/D repeater241/X vssd1 vssd1 vccd1 vccd1 _21214_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_191_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21145_ _21147_/CLK _21145_/D repeater215/X vssd1 vssd1 vccd1 vccd1 _21145_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_116_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09907_ _21255_/Q vssd1 vssd1 vccd1 vccd1 _09907_/Y sky130_fd_sc_hd__inv_2
X_21076_ _21087_/CLK _21076_/D repeater228/X vssd1 vssd1 vccd1 vccd1 _21076_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_76_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_247_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20027_ _21486_/CLK _20027_/D repeater209/X vssd1 vssd1 vccd1 vccd1 _20027_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_247_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09838_ _15881_/A vssd1 vssd1 vccd1 vccd1 _09838_/X sky130_fd_sc_hd__buf_1
XFILLER_74_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09769_ _09769_/A _09769_/B _09769_/C _09769_/D vssd1 vssd1 vccd1 vccd1 _14309_/A
+ sky130_fd_sc_hd__and4_4
XFILLER_74_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11800_ _11800_/A vssd1 vssd1 vccd1 vccd1 _12968_/A sky130_fd_sc_hd__buf_2
XPHY_4034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18565__A0 _17079_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12780_ _20791_/Q _12777_/X _09633_/X _12778_/X vssd1 vssd1 vccd1 vccd1 _20791_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11731_ _21062_/Q _11727_/X _11684_/X _11729_/X vssd1 vssd1 vccd1 vccd1 _21062_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20929_ _20929_/CLK _20929_/D repeater266/X vssd1 vssd1 vccd1 vccd1 _20929_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_203_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18526__S _18906_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16835__A _16835_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13929__A1 _13928_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14450_ _14401_/X _14450_/B _14450_/C _14450_/D vssd1 vssd1 vccd1 vccd1 _14464_/B
+ sky130_fd_sc_hd__and4b_1
XPHY_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11662_ _11504_/X _11652_/X _19112_/S _11659_/Y _21093_/Q vssd1 vssd1 vccd1 vccd1
+ _21093_/D sky130_fd_sc_hd__a32o_1
XANTENNA_clkbuf_leaf_60_HCLK_A clkbuf_4_14_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18317__A0 _18848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13401_ _20491_/Q _13398_/X _13280_/X _13399_/X vssd1 vssd1 vccd1 vccd1 _20491_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10613_ _21326_/Q _10609_/Y _21320_/Q _10610_/Y _10612_/X vssd1 vssd1 vccd1 vccd1
+ _10622_/B sky130_fd_sc_hd__o221a_1
XPHY_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14381_ _20238_/Q _14467_/A vssd1 vssd1 vccd1 vccd1 _14382_/B sky130_fd_sc_hd__nand2_1
XPHY_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11593_ _11589_/Y _11592_/Y _11017_/A _11587_/X vssd1 vssd1 vccd1 vccd1 _21123_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_167_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16120_ _20327_/Q vssd1 vssd1 vccd1 vccd1 _16120_/X sky130_fd_sc_hd__clkbuf_2
X_10544_ _21315_/Q vssd1 vssd1 vccd1 vccd1 _10703_/A sky130_fd_sc_hd__inv_2
X_13332_ _13357_/A vssd1 vssd1 vccd1 vccd1 _13359_/A sky130_fd_sc_hd__inv_2
XPHY_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16051_ _16057_/A vssd1 vssd1 vccd1 vccd1 _16051_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13263_ _13299_/A vssd1 vssd1 vccd1 vccd1 _13293_/A sky130_fd_sc_hd__buf_1
XANTENNA__15551__B1 _15550_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10475_ _20681_/Q vssd1 vssd1 vccd1 vccd1 _10475_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18261__S _18910_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15002_ _15002_/A _15002_/B vssd1 vssd1 vccd1 vccd1 _15012_/A sky130_fd_sc_hd__or2_1
X_12214_ _20944_/Q vssd1 vssd1 vccd1 vccd1 _12432_/C sky130_fd_sc_hd__inv_2
XANTENNA__17828__C1 _17827_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13194_ _13227_/A vssd1 vssd1 vccd1 vccd1 _13217_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_151_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12145_ _12103_/X _12145_/B _12145_/C _12145_/D vssd1 vssd1 vccd1 vccd1 _12145_/X
+ sky130_fd_sc_hd__and4b_1
X_19810_ _19812_/CLK _19810_/D vssd1 vssd1 vccd1 vccd1 _19810_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17843__A2 _17839_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20554__CLK _20592_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12076_ _20386_/Q vssd1 vssd1 vccd1 vccd1 _18000_/A sky130_fd_sc_hd__inv_2
X_16953_ _19967_/Q vssd1 vssd1 vccd1 vccd1 _16958_/A sky130_fd_sc_hd__buf_1
X_19741_ _19811_/CLK _19741_/D vssd1 vssd1 vccd1 vccd1 _19741_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20708__RESET_B repeater210/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19092__S _19870_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15904_ _15911_/A vssd1 vssd1 vccd1 vccd1 _15904_/X sky130_fd_sc_hd__buf_1
X_11027_ _19952_/Q _16886_/A _19953_/Q vssd1 vssd1 vccd1 vccd1 _16896_/A sky130_fd_sc_hd__or3_1
XFILLER_237_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19672_ _19821_/CLK _19672_/D vssd1 vssd1 vccd1 vccd1 _19672_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__19140__S1 _21017_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16884_ _16894_/A _19950_/Q vssd1 vssd1 vccd1 vccd1 _16884_/Y sky130_fd_sc_hd__nor2_1
XFILLER_37_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18623_ _18848_/A0 _18070_/Y _18666_/S vssd1 vssd1 vccd1 vccd1 _18623_/X sky130_fd_sc_hd__mux2_1
XFILLER_92_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15835_ _15841_/A vssd1 vssd1 vccd1 vccd1 _15842_/A sky130_fd_sc_hd__inv_2
XANTENNA__13617__B1 _13555_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18554_ _18553_/X _12169_/Y _18909_/S vssd1 vssd1 vccd1 vccd1 _18554_/X sky130_fd_sc_hd__mux2_1
X_15766_ _15766_/A vssd1 vssd1 vccd1 vccd1 _15766_/X sky130_fd_sc_hd__buf_1
X_12978_ _13600_/A vssd1 vssd1 vccd1 vccd1 _12978_/X sky130_fd_sc_hd__buf_1
XFILLER_206_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_233_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17505_ _21023_/Q _17425_/X _17502_/X _17503_/X _17504_/Y vssd1 vssd1 vccd1 vccd1
+ _17505_/X sky130_fd_sc_hd__o221a_1
X_14717_ _14723_/A vssd1 vssd1 vccd1 vccd1 _14717_/X sky130_fd_sc_hd__buf_1
XANTENNA__12840__A1 _20758_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18485_ _18484_/X _15141_/Y _18784_/S vssd1 vssd1 vccd1 vccd1 _18485_/X sky130_fd_sc_hd__mux2_2
X_11929_ _11929_/A vssd1 vssd1 vccd1 vccd1 _11930_/A sky130_fd_sc_hd__inv_2
XFILLER_233_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15697_ _15788_/A vssd1 vssd1 vccd1 vccd1 _15697_/X sky130_fd_sc_hd__buf_1
XANTENNA__18436__S _18885_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17436_ _19489_/Q vssd1 vssd1 vccd1 vccd1 _17436_/Y sky130_fd_sc_hd__inv_2
X_14648_ _14648_/A vssd1 vssd1 vccd1 vccd1 _14648_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_221_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17367_ _19335_/Q vssd1 vssd1 vccd1 vccd1 _17368_/A sky130_fd_sc_hd__inv_2
X_14579_ _14579_/A _14579_/B vssd1 vssd1 vccd1 vccd1 _14627_/A sky130_fd_sc_hd__or2_1
XANTENNA__15790__B1 _15788_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19106_ _16664_/Y _21072_/Q _19870_/D vssd1 vssd1 vccd1 vccd1 _19106_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16318_ _19378_/Q _16312_/X _16006_/X _16314_/X vssd1 vssd1 vccd1 vccd1 _19378_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_158_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17298_ _17285_/Y _17286_/X _17288_/X _17297_/X vssd1 vssd1 vccd1 vccd1 _17298_/X
+ sky130_fd_sc_hd__o211a_2
X_19037_ _16841_/Y _20832_/Q _19046_/S vssd1 vssd1 vccd1 vccd1 _19939_/D sky130_fd_sc_hd__mux2_1
X_16249_ _16255_/A vssd1 vssd1 vccd1 vccd1 _16256_/A sky130_fd_sc_hd__inv_2
XANTENNA__18171__S _18886_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput102 _18097_/Y vssd1 vssd1 vccd1 vccd1 HRDATA[30] sky130_fd_sc_hd__clkbuf_2
XFILLER_133_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput113 _17091_/X vssd1 vssd1 vccd1 vccd1 IRQ[10] sky130_fd_sc_hd__clkbuf_2
XFILLER_127_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput124 _17086_/X vssd1 vssd1 vccd1 vccd1 IRQ[6] sky130_fd_sc_hd__clkbuf_2
Xoutput135 _17043_/Y vssd1 vssd1 vccd1 vccd1 SSn_S3 sky130_fd_sc_hd__clkbuf_2
XFILLER_142_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15096__A _20451_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19939_ _20930_/CLK _19939_/D repeater269/X vssd1 vssd1 vccd1 vccd1 _19939_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_229_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09623_ _09677_/A vssd1 vssd1 vccd1 vccd1 _09660_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_44_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18547__A0 _18848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_197_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18346__S _18787_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20714_ _21366_/CLK _20714_/D repeater254/X vssd1 vssd1 vccd1 vccd1 _20714_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_12_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19198__S1 _20131_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20645_ _20657_/CLK _20645_/D repeater198/X vssd1 vssd1 vccd1 vccd1 _20645_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21237__RESET_B repeater249/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20576_ _20946_/CLK _20576_/D repeater275/X vssd1 vssd1 vccd1 vccd1 _20576_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_176_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15533__B1 _15454_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10260_ _10260_/A _10260_/B vssd1 vssd1 vccd1 vccd1 _10418_/A sky130_fd_sc_hd__or2_1
X_10191_ _21393_/Q _10190_/Y _10183_/X _10155_/B vssd1 vssd1 vccd1 vccd1 _21393_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_160_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20872__RESET_B repeater247/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21128_ _21134_/CLK _21128_/D repeater192/X vssd1 vssd1 vccd1 vccd1 _21128_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_78_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20801__RESET_B repeater252/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21059_ _21147_/CLK _21059_/D repeater230/X vssd1 vssd1 vccd1 vccd1 _21059_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_87_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13950_ _20646_/Q _13972_/C _13948_/Y _20303_/Q _13949_/X vssd1 vssd1 vccd1 vccd1
+ _13950_/X sky130_fd_sc_hd__a221o_1
XANTENNA__18786__A0 _17079_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20119__RESET_B repeater247/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10125__A2 _20774_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12901_ _12924_/A vssd1 vssd1 vccd1 vccd1 _12901_/X sky130_fd_sc_hd__buf_1
X_13881_ _13971_/C _13881_/B vssd1 vssd1 vccd1 vccd1 _14002_/A sky130_fd_sc_hd__or2_1
XFILLER_100_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15620_ _19713_/Q _15618_/X _15480_/X _15619_/X vssd1 vssd1 vccd1 vccd1 _19713_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13254__A _13600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12832_ _20764_/Q _12829_/X _12666_/X _12830_/X vssd1 vssd1 vccd1 vccd1 _20764_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18538__A0 _18537_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14272__B1 _13714_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_215_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_opt_5_HCLK_A clkbuf_opt_7_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15551_ _19747_/Q _15543_/X _15550_/X _15546_/X vssd1 vssd1 vccd1 vccd1 _19747_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12763_ _20802_/Q _12757_/X _12658_/X _12760_/X vssd1 vssd1 vccd1 vccd1 _20802_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_243_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18256__S _18896_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_230_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14502_ _14502_/A _14502_/B vssd1 vssd1 vccd1 vccd1 _14507_/A sky130_fd_sc_hd__or2_1
XPHY_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11714_ _11720_/A vssd1 vssd1 vccd1 vccd1 _11721_/A sky130_fd_sc_hd__inv_2
XPHY_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18270_ _17811_/Y _20746_/Q _18879_/S vssd1 vssd1 vccd1 vccd1 _18270_/X sky130_fd_sc_hd__mux2_1
XFILLER_159_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15482_ _19777_/Q _15479_/X _15480_/X _15481_/X vssd1 vssd1 vccd1 vccd1 _19777_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12694_ _12708_/A vssd1 vssd1 vccd1 vccd1 _12694_/X sky130_fd_sc_hd__buf_1
XPHY_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17221_ _18904_/X _17211_/X _18892_/X _17214_/X _17220_/X vssd1 vssd1 vccd1 vccd1
+ _17235_/C sky130_fd_sc_hd__o221a_2
X_14433_ _14430_/Y _20226_/Q _14431_/Y _20221_/Q _14432_/X vssd1 vssd1 vccd1 vccd1
+ _14434_/D sky130_fd_sc_hd__o221a_1
XANTENNA__19189__S1 _20122_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11645_ _18979_/X _11640_/X _21101_/Q _11642_/X vssd1 vssd1 vccd1 vccd1 _21101_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17152_ _21044_/Q vssd1 vssd1 vccd1 vccd1 _17152_/Y sky130_fd_sc_hd__inv_2
XPHY_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14364_ _14460_/D _14364_/B vssd1 vssd1 vccd1 vccd1 _14493_/A sky130_fd_sc_hd__or2_1
Xinput15 HADDR[22] vssd1 vssd1 vccd1 vccd1 input15/X sky130_fd_sc_hd__clkbuf_1
X_11576_ _16546_/A _19993_/Q vssd1 vssd1 vccd1 vccd1 _11577_/A sky130_fd_sc_hd__nand2_1
Xinput26 HADDR[3] vssd1 vssd1 vccd1 vccd1 input26/X sky130_fd_sc_hd__buf_1
XPHY_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput37 HTRANS[1] vssd1 vssd1 vccd1 vccd1 input37/X sky130_fd_sc_hd__clkbuf_2
XPHY_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16103_ _19481_/Q _16101_/X _15876_/X _16102_/X vssd1 vssd1 vccd1 vccd1 _19481_/D
+ sky130_fd_sc_hd__a22o_1
Xinput48 HWDATA[19] vssd1 vssd1 vccd1 vccd1 input48/X sky130_fd_sc_hd__clkbuf_4
XFILLER_7_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput59 HWDATA[29] vssd1 vssd1 vccd1 vccd1 input59/X sky130_fd_sc_hd__buf_4
X_13315_ _13321_/A vssd1 vssd1 vccd1 vccd1 _13315_/X sky130_fd_sc_hd__buf_1
X_17083_ _17083_/A vssd1 vssd1 vccd1 vccd1 _17814_/A sky130_fd_sc_hd__inv_2
X_10527_ _20735_/Q vssd1 vssd1 vccd1 vccd1 _10527_/Y sky130_fd_sc_hd__inv_2
X_14295_ _14292_/X _14294_/Y _14292_/X _14294_/Y vssd1 vssd1 vccd1 vccd1 _14302_/C
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_155_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16034_ _16034_/A _16229_/B _16229_/C vssd1 vssd1 vccd1 vccd1 _16042_/A sky130_fd_sc_hd__or3_4
X_10458_ _10783_/A _20696_/Q _21307_/Q _10454_/Y _10457_/X vssd1 vssd1 vccd1 vccd1
+ _10471_/B sky130_fd_sc_hd__o221a_1
X_13246_ _20570_/Q _13239_/X _13245_/X _13241_/X vssd1 vssd1 vccd1 vccd1 _20570_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18004__B _18006_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13429__A input40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10389_ _21363_/Q _10388_/Y _10373_/X _10279_/B vssd1 vssd1 vccd1 vccd1 _21363_/D
+ sky130_fd_sc_hd__o211a_1
X_13177_ _20598_/Q _13717_/B vssd1 vssd1 vccd1 vccd1 _13177_/Y sky130_fd_sc_hd__nor2_1
XFILLER_123_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12128_ _20390_/Q vssd1 vssd1 vccd1 vccd1 _12128_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17985_ _18366_/X _17947_/X _18339_/X _17948_/X vssd1 vssd1 vccd1 vccd1 _17989_/A
+ sky130_fd_sc_hd__o22ai_2
XFILLER_123_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20542__RESET_B repeater264/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12059_ _20971_/Q _12054_/Y _20950_/Q _12055_/Y _12058_/X vssd1 vssd1 vccd1 vccd1
+ _12060_/D sky130_fd_sc_hd__o221a_1
X_16936_ _19963_/Q vssd1 vssd1 vccd1 vccd1 _16936_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19724_ _20432_/CLK _19724_/D vssd1 vssd1 vccd1 vccd1 _19724_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18777__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18020__A _18020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16867_ _19946_/Q vssd1 vssd1 vccd1 vccd1 _16867_/Y sky130_fd_sc_hd__inv_2
X_19655_ _21021_/CLK _19655_/D vssd1 vssd1 vccd1 vccd1 _19655_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18606_ _18605_/X _13738_/X _18748_/S vssd1 vssd1 vccd1 vccd1 _18606_/X sky130_fd_sc_hd__mux2_2
X_15818_ _15824_/A vssd1 vssd1 vccd1 vccd1 _15825_/A sky130_fd_sc_hd__inv_2
X_19586_ _21218_/CLK _19586_/D vssd1 vssd1 vccd1 vccd1 _19586_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14263__B1 _14262_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16798_ _19930_/Q _16794_/A _16797_/Y _16794_/Y vssd1 vssd1 vccd1 vccd1 _16799_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_240_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18537_ _17937_/Y _20349_/Q _18787_/S vssd1 vssd1 vccd1 vccd1 _18537_/X sky130_fd_sc_hd__mux2_1
XFILLER_80_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15749_ _19650_/Q _15743_/X _15694_/X _15745_/X vssd1 vssd1 vccd1 vccd1 _19650_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18166__S _18896_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_240_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18468_ _18467_/X _14402_/Y _18897_/S vssd1 vssd1 vccd1 vccd1 _18468_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17419_ _19713_/Q vssd1 vssd1 vccd1 vccd1 _17419_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21330__RESET_B repeater204/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18399_ _18845_/A0 _10304_/Y _18884_/S vssd1 vssd1 vccd1 vccd1 _18399_/X sky130_fd_sc_hd__mux2_1
X_20430_ _21001_/CLK _20430_/D repeater190/X vssd1 vssd1 vccd1 vccd1 _20430_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_158_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20361_ _20951_/CLK _20361_/D repeater272/X vssd1 vssd1 vccd1 vccd1 _20361_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_174_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20292_ _20661_/CLK _20292_/D repeater263/X vssd1 vssd1 vccd1 vccd1 _20292_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_103_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20283__RESET_B repeater262/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20212__RESET_B repeater203/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_229_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09606_ _13110_/A vssd1 vssd1 vccd1 vccd1 _13108_/A sky130_fd_sc_hd__buf_1
XFILLER_113_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15203__C1 _15160_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18804__S _18880_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11430_ _19916_/Q vssd1 vssd1 vccd1 vccd1 _11430_/Y sky130_fd_sc_hd__inv_2
XPHY_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20628_ _20697_/CLK _20628_/D repeater196/X vssd1 vssd1 vccd1 vccd1 _20628_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21000__RESET_B repeater190/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11361_ _21178_/Q vssd1 vssd1 vccd1 vccd1 _11363_/B sky130_fd_sc_hd__inv_2
XANTENNA__11240__B1 _19910_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15729__A input66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20559_ _20592_/CLK _20559_/D repeater260/X vssd1 vssd1 vccd1 vccd1 _20559_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_22_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10312_ _20733_/Q vssd1 vssd1 vccd1 vccd1 _10312_/Y sky130_fd_sc_hd__inv_2
X_13100_ _20637_/Q _13098_/X _12875_/X _13099_/X vssd1 vssd1 vccd1 vccd1 _20637_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_3_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11292_ _12502_/A _12500_/A _11545_/A _12504_/A vssd1 vssd1 vccd1 vccd1 _11322_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_152_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14080_ _14080_/A _14212_/A vssd1 vssd1 vccd1 vccd1 _14081_/B sky130_fd_sc_hd__or2_2
Xclkbuf_leaf_30_HCLK clkbuf_opt_4_HCLK/A vssd1 vssd1 vccd1 vccd1 _21423_/CLK sky130_fd_sc_hd__clkbuf_16
X_13031_ _20675_/Q _13026_/X _13030_/X _13027_/X vssd1 vssd1 vccd1 vccd1 _20675_/D
+ sky130_fd_sc_hd__a22o_1
X_10243_ _21360_/Q vssd1 vssd1 vccd1 vccd1 _10275_/A sky130_fd_sc_hd__inv_2
XFILLER_161_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input45_A HWDATA[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10174_ _21402_/Q _10169_/C _10170_/X _10172_/A vssd1 vssd1 vccd1 vccd1 _21402_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_121_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17770_ _19445_/Q vssd1 vssd1 vccd1 vccd1 _17770_/Y sky130_fd_sc_hd__inv_2
X_14982_ _20097_/Q _14981_/Y _14973_/X _14876_/B vssd1 vssd1 vccd1 vccd1 _20097_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_78_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16721_ _20983_/Q vssd1 vssd1 vccd1 vccd1 _16721_/Y sky130_fd_sc_hd__inv_2
X_13933_ _20656_/Q _13848_/A _20654_/Q _13971_/B vssd1 vssd1 vccd1 vccd1 _13933_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_219_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19440_ _21234_/CLK _19440_/D vssd1 vssd1 vccd1 vccd1 _19440_/Q sky130_fd_sc_hd__dfxtp_1
X_16652_ _16652_/A _18954_/X vssd1 vssd1 vccd1 vccd1 _19860_/D sky130_fd_sc_hd__and2_1
XFILLER_47_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13864_ _20292_/Q vssd1 vssd1 vccd1 vccd1 _14031_/C sky130_fd_sc_hd__inv_2
XFILLER_234_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19765__CLK _19765_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15603_ _15603_/A vssd1 vssd1 vccd1 vccd1 _15603_/X sky130_fd_sc_hd__buf_1
XFILLER_16_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19371_ _19789_/CLK _19371_/D vssd1 vssd1 vccd1 vccd1 _19371_/Q sky130_fd_sc_hd__dfxtp_1
X_12815_ _12815_/A _13108_/B vssd1 vssd1 vccd1 vccd1 _12816_/S sky130_fd_sc_hd__or2_1
X_16583_ _16583_/A _16583_/B vssd1 vssd1 vccd1 vccd1 _16744_/B sky130_fd_sc_hd__or2_1
XFILLER_222_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13795_ _20199_/Q vssd1 vssd1 vccd1 vccd1 _14588_/A sky130_fd_sc_hd__inv_2
XFILLER_27_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_repeater184_A repeater185/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_188_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18322_ _17281_/X _18017_/Y _18835_/S vssd1 vssd1 vccd1 vccd1 _18322_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13712__A _15429_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15534_ _19755_/Q _15529_/X _15456_/X _15531_/X vssd1 vssd1 vccd1 vccd1 _19755_/D
+ sky130_fd_sc_hd__a22o_1
X_12746_ _20807_/Q _12746_/B _12751_/B vssd1 vssd1 vccd1 vccd1 _12746_/X sky130_fd_sc_hd__or3_2
XFILLER_188_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14527__B _17169_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18253_ _18845_/A0 _10507_/Y _18896_/S vssd1 vssd1 vccd1 vccd1 _18253_/X sky130_fd_sc_hd__mux2_1
XFILLER_187_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15465_ _15638_/C vssd1 vssd1 vccd1 vccd1 _16616_/B sky130_fd_sc_hd__buf_1
XFILLER_230_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12677_ _20832_/Q _12672_/X _09626_/X _12674_/X vssd1 vssd1 vccd1 vccd1 _20832_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18714__S _18879_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17204_ _17204_/A vssd1 vssd1 vccd1 vccd1 _18021_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_187_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14416_ _20032_/Q vssd1 vssd1 vccd1 vccd1 _14416_/Y sky130_fd_sc_hd__inv_2
XPHY_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11628_ _11628_/A vssd1 vssd1 vccd1 vccd1 _11628_/Y sky130_fd_sc_hd__inv_2
X_18184_ _17809_/Y _20642_/Q _18903_/S vssd1 vssd1 vccd1 vccd1 _18184_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17838__B _17838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15396_ _15505_/A _15396_/B _16594_/B vssd1 vssd1 vccd1 vccd1 _16311_/C sky130_fd_sc_hd__or3_4
XFILLER_184_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17135_ _17286_/A vssd1 vssd1 vccd1 vccd1 _17136_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_14347_ _20213_/Q vssd1 vssd1 vccd1 vccd1 _14498_/A sky130_fd_sc_hd__inv_2
XFILLER_155_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11559_ _16332_/A vssd1 vssd1 vccd1 vccd1 _13163_/A sky130_fd_sc_hd__buf_4
XFILLER_183_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18015__A _20456_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20794__RESET_B repeater252/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17066_ _17072_/B _17066_/B vssd1 vssd1 vccd1 vccd1 _19909_/D sky130_fd_sc_hd__nor2_1
XFILLER_155_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14278_ _20121_/Q vssd1 vssd1 vccd1 vccd1 _14288_/A sky130_fd_sc_hd__inv_2
XFILLER_143_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20723__RESET_B repeater264/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16017_ _19526_/Q _16008_/X _16016_/X _16010_/X vssd1 vssd1 vccd1 vccd1 _19526_/D
+ sky130_fd_sc_hd__a22o_1
X_13229_ _20580_/Q _13226_/X _13140_/X _13228_/X vssd1 vssd1 vccd1 vccd1 _20580_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17854__A _17854_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19295__CLK _19813_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17968_ _20416_/Q vssd1 vssd1 vccd1 vccd1 _17968_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_214_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19707_ _19789_/CLK _19707_/D vssd1 vssd1 vccd1 vccd1 _19707_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_226_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16919_ _19958_/Q _16913_/A _16917_/Y _16913_/Y vssd1 vssd1 vccd1 vccd1 _16920_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_65_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17899_ _17974_/A vssd1 vssd1 vccd1 vccd1 _17938_/B sky130_fd_sc_hd__buf_4
XFILLER_53_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19638_ _20326_/CLK _19638_/D vssd1 vssd1 vccd1 vccd1 _19638_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_214_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19569_ _19812_/CLK _19569_/D vssd1 vssd1 vccd1 vccd1 _19569_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_213_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_222_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19270__S0 _20130_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12262__A2 _20504_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19906__RESET_B repeater202/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18624__S _18667_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11142__A _21005_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21462_ _21462_/CLK _21462_/D repeater245/X vssd1 vssd1 vccd1 vccd1 _21462_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_182_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_53_HCLK clkbuf_4_9_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _21147_/CLK sky130_fd_sc_hd__clkbuf_16
X_20413_ _20413_/CLK _20413_/D repeater185/X vssd1 vssd1 vccd1 vccd1 _20413_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_135_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11222__B1 _10886_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21393_ _21401_/CLK _21393_/D repeater253/X vssd1 vssd1 vccd1 vccd1 _21393_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_134_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20344_ _21372_/CLK _20344_/D repeater269/X vssd1 vssd1 vccd1 vccd1 _20344_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_134_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20275_ _20286_/CLK _20275_/D repeater265/X vssd1 vssd1 vccd1 vccd1 _20275_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_103_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12701__A _12707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10930_ _21211_/Q _21038_/Q _10928_/Y _11815_/A vssd1 vssd1 vccd1 vccd1 _10931_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_83_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20765__CLK _21342_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10861_ _10908_/A _10908_/B _17370_/A vssd1 vssd1 vccd1 vccd1 _10862_/S sky130_fd_sc_hd__or3_1
XFILLER_232_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12600_ _12600_/A vssd1 vssd1 vccd1 vccd1 _12600_/X sky130_fd_sc_hd__clkbuf_4
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12789__B1 _09649_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13580_ _13594_/A vssd1 vssd1 vccd1 vccd1 _13580_/X sky130_fd_sc_hd__buf_1
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_242_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10792_ _10781_/A _10781_/B _10824_/A _10790_/Y vssd1 vssd1 vccd1 vccd1 _21305_/D
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__19261__S0 _20132_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_212_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12531_ _11286_/C _12520_/X _11545_/A _12521_/X vssd1 vssd1 vccd1 vccd1 _20911_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18534__S _18904_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15250_ _15250_/A _15250_/B _15250_/C _15250_/D vssd1 vssd1 vccd1 vccd1 _15250_/X
+ sky130_fd_sc_hd__and4_1
X_12462_ _12462_/A vssd1 vssd1 vccd1 vccd1 _12480_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_200_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14201_ _14201_/A vssd1 vssd1 vccd1 vccd1 _14201_/Y sky130_fd_sc_hd__inv_2
X_11413_ _11421_/A _11413_/B vssd1 vssd1 vccd1 vccd1 _11413_/X sky130_fd_sc_hd__or2_2
XFILLER_153_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15181_ _15181_/A vssd1 vssd1 vccd1 vccd1 _15181_/Y sky130_fd_sc_hd__inv_2
X_12393_ _20396_/Q vssd1 vssd1 vccd1 vccd1 _12469_/B sky130_fd_sc_hd__inv_2
XFILLER_137_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_115_HCLK_A clkbuf_opt_3_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14132_ _20530_/Q _14070_/A _14129_/Y _20278_/Q _14131_/X vssd1 vssd1 vccd1 vccd1
+ _14138_/C sky130_fd_sc_hd__o221a_1
XFILLER_137_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11344_ _21183_/Q _21182_/Q vssd1 vssd1 vccd1 vccd1 _11783_/C sky130_fd_sc_hd__or2_2
XFILLER_153_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18940_ _16704_/X _21136_/Q _18946_/S vssd1 vssd1 vccd1 vccd1 _18940_/X sky130_fd_sc_hd__mux2_1
X_14063_ _20265_/Q vssd1 vssd1 vccd1 vccd1 _14076_/A sky130_fd_sc_hd__inv_2
X_11275_ _20913_/Q vssd1 vssd1 vccd1 vccd1 _11541_/B sky130_fd_sc_hd__inv_2
XFILLER_79_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20134__RESET_B repeater248/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13014_ _20685_/Q _13012_/X _12925_/X _13013_/X vssd1 vssd1 vccd1 vccd1 _20685_/D
+ sky130_fd_sc_hd__a22o_1
X_10226_ _10221_/A _10221_/B _10221_/C vssd1 vssd1 vccd1 vccd1 _10227_/B sky130_fd_sc_hd__o21a_1
X_18871_ _17193_/Y _16894_/A _18899_/S vssd1 vssd1 vccd1 vccd1 _18871_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13707__A _15424_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17822_ _18403_/X _17951_/A _18405_/X _17952_/A vssd1 vssd1 vccd1 vccd1 _17827_/A
+ sky130_fd_sc_hd__a22oi_1
X_10157_ _10157_/A _10157_/B vssd1 vssd1 vccd1 vccd1 _10182_/A sky130_fd_sc_hd__or2_1
XFILLER_67_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14965_ _14965_/A _14965_/B _14965_/C _14964_/X vssd1 vssd1 vccd1 vccd1 _14965_/X
+ sky130_fd_sc_hd__or4b_4
X_17753_ _19405_/Q vssd1 vssd1 vccd1 vccd1 _17753_/Y sky130_fd_sc_hd__inv_2
X_10088_ _10052_/C _20784_/Q _21387_/Q _10085_/Y _10087_/X vssd1 vssd1 vccd1 vccd1
+ _10098_/B sky130_fd_sc_hd__o221a_1
XFILLER_248_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18709__S _18835_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17404__B1 _18813_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16704_ _19896_/Q _14236_/B _14237_/B vssd1 vssd1 vccd1 vccd1 _16704_/X sky130_fd_sc_hd__a21bo_1
X_13916_ _20658_/Q _20315_/Q _13915_/Y _13891_/A vssd1 vssd1 vccd1 vccd1 _13922_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_48_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17684_ _17684_/A vssd1 vssd1 vccd1 vccd1 _17775_/B sky130_fd_sc_hd__buf_1
X_14896_ _20575_/Q vssd1 vssd1 vccd1 vccd1 _14896_/Y sky130_fd_sc_hd__inv_2
X_16635_ _19852_/Q _19853_/Q _15288_/B vssd1 vssd1 vccd1 vccd1 _16635_/X sky130_fd_sc_hd__a21bo_1
XFILLER_74_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19423_ _19521_/CLK _19423_/D vssd1 vssd1 vccd1 vccd1 _19423_/Q sky130_fd_sc_hd__dfxtp_1
X_13847_ _20313_/Q vssd1 vssd1 vccd1 vccd1 _13848_/A sky130_fd_sc_hd__inv_2
XFILLER_204_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13442__A _15421_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16566_ _16566_/A _16609_/A _16566_/C vssd1 vssd1 vccd1 vccd1 _16566_/X sky130_fd_sc_hd__or3_4
X_19354_ _21453_/CLK _19354_/D vssd1 vssd1 vccd1 vccd1 _19354_/Q sky130_fd_sc_hd__dfxtp_1
X_13778_ _20627_/Q _14593_/A _13777_/Y _20204_/Q vssd1 vssd1 vccd1 vccd1 _13778_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__19252__S0 _19275_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_76_HCLK clkbuf_4_13_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20693_/CLK sky130_fd_sc_hd__clkbuf_16
X_18305_ _18304_/X _14922_/Y _18907_/S vssd1 vssd1 vccd1 vccd1 _18305_/X sky130_fd_sc_hd__mux2_1
X_15517_ input63/X vssd1 vssd1 vccd1 vccd1 _15788_/A sky130_fd_sc_hd__buf_1
XFILLER_176_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12729_ _11179_/X _20808_/Q _12729_/S vssd1 vssd1 vccd1 vccd1 _20808_/D sky130_fd_sc_hd__mux2_1
X_19285_ _19661_/Q _19653_/Q _19637_/Q _19821_/Q _19285_/S0 _21017_/Q vssd1 vssd1
+ vccd1 vccd1 _19285_/X sky130_fd_sc_hd__mux4_2
X_16497_ _20002_/Q vssd1 vssd1 vccd1 vccd1 _16498_/A sky130_fd_sc_hd__inv_2
XANTENNA__18444__S _18910_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_230_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20975__RESET_B repeater278/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18236_ _20860_/Q input9/X _18236_/S vssd1 vssd1 vccd1 vccd1 _18236_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15448_ _15448_/A _15624_/B _15999_/C vssd1 vssd1 vccd1 vccd1 _15459_/A sky130_fd_sc_hd__or3_4
XANTENNA__15194__A1 _15099_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20904__RESET_B repeater217/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18167_ _18166_/X _10601_/Y _18891_/S vssd1 vssd1 vccd1 vccd1 _18167_/X sky130_fd_sc_hd__mux2_1
X_15379_ _15389_/A vssd1 vssd1 vccd1 vccd1 _15390_/A sky130_fd_sc_hd__inv_2
XFILLER_184_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17118_ _19622_/Q vssd1 vssd1 vccd1 vccd1 _17118_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12952__B1 _12950_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18098_ _20464_/Q vssd1 vssd1 vccd1 vccd1 _18098_/Y sky130_fd_sc_hd__inv_2
X_17049_ _20039_/Q _20037_/Q vssd1 vssd1 vccd1 vccd1 _17049_/X sky130_fd_sc_hd__or2_1
XFILLER_104_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09940_ _20871_/Q vssd1 vssd1 vccd1 vccd1 _11488_/B sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_37_HCLK_A _20004_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12704__B1 _12548_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20060_ _20066_/CLK _20060_/D repeater281/X vssd1 vssd1 vccd1 vccd1 _20060_/Q sky130_fd_sc_hd__dfrtp_4
X_09871_ _09871_/A vssd1 vssd1 vccd1 vccd1 _14307_/B sky130_fd_sc_hd__inv_2
XFILLER_140_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater210 repeater211/X vssd1 vssd1 vccd1 vccd1 repeater210/X sky130_fd_sc_hd__clkbuf_8
XFILLER_39_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater221 repeater223/X vssd1 vssd1 vccd1 vccd1 repeater221/X sky130_fd_sc_hd__buf_8
XFILLER_57_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrepeater232 repeater234/X vssd1 vssd1 vccd1 vccd1 repeater232/X sky130_fd_sc_hd__buf_4
Xrepeater243 repeater244/X vssd1 vssd1 vccd1 vccd1 repeater243/X sky130_fd_sc_hd__buf_8
Xrepeater254 repeater255/X vssd1 vssd1 vccd1 vccd1 repeater254/X sky130_fd_sc_hd__buf_8
XANTENNA__18619__S _18904_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater265 repeater267/X vssd1 vssd1 vccd1 vccd1 repeater265/X sky130_fd_sc_hd__clkbuf_8
Xrepeater276 repeater277/X vssd1 vssd1 vccd1 vccd1 repeater276/X sky130_fd_sc_hd__clkbuf_8
XPHY_4408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20962_ _20981_/CLK _20962_/D repeater186/X vssd1 vssd1 vccd1 vccd1 _20962_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_3707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15957__B1 _15887_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_214_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20893_ _21141_/CLK _20893_/D repeater192/X vssd1 vssd1 vccd1 vccd1 _20893_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__19243__S0 _19275_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16663__A _16663_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18354__S _18850_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13196__B1 _12984_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21445_ _21445_/CLK _21445_/D repeater244/X vssd1 vssd1 vccd1 vccd1 _21445_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_119_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21376_ _21406_/CLK _21376_/D repeater213/X vssd1 vssd1 vccd1 vccd1 _21376_/Q sky130_fd_sc_hd__dfrtp_1
X_20327_ _20327_/CLK _20327_/D repeater235/X vssd1 vssd1 vccd1 vccd1 _20327_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_190_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11060_ _11060_/A _11080_/A vssd1 vssd1 vccd1 vccd1 _11074_/A sky130_fd_sc_hd__or2_1
XFILLER_134_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20258_ _20915_/CLK _20258_/D repeater217/X vssd1 vssd1 vccd1 vccd1 _20258_/Q sky130_fd_sc_hd__dfstp_1
X_10011_ _21415_/Q _17032_/A _10008_/Y _10009_/Y _10010_/Y vssd1 vssd1 vccd1 vccd1
+ _10011_/X sky130_fd_sc_hd__o221a_1
XFILLER_95_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20189_ _21485_/CLK _20189_/D repeater200/X vssd1 vssd1 vccd1 vccd1 _20189_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_192_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17941__B _17943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18529__S _18748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14750_ _19123_/X vssd1 vssd1 vccd1 vccd1 _14753_/A sky130_fd_sc_hd__inv_2
Xclkbuf_1_1_1_HCLK clkbuf_1_1_1_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_11962_ _13182_/A vssd1 vssd1 vccd1 vccd1 _16515_/A sky130_fd_sc_hd__buf_1
XFILLER_233_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13701_ _20339_/Q _13699_/X _13506_/X _13700_/X vssd1 vssd1 vccd1 vccd1 _20339_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_45_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_99_HCLK clkbuf_4_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20665_/CLK sky130_fd_sc_hd__clkbuf_16
X_10913_ _20171_/Q vssd1 vssd1 vccd1 vccd1 _10918_/A sky130_fd_sc_hd__inv_2
XFILLER_72_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14681_ _10917_/A _14680_/X _14676_/Y vssd1 vssd1 vccd1 vccd1 _20170_/D sky130_fd_sc_hd__a21oi_1
X_11893_ _21021_/Q _11883_/X _11877_/A _11892_/X vssd1 vssd1 vccd1 vccd1 _21021_/D
+ sky130_fd_sc_hd__a31o_1
XANTENNA__10886__A _12548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16420_ _16427_/A vssd1 vssd1 vccd1 vccd1 _16420_/X sky130_fd_sc_hd__buf_1
XANTENNA__13262__A _17080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13632_ _13651_/A vssd1 vssd1 vccd1 vccd1 _13632_/X sky130_fd_sc_hd__buf_1
X_10844_ _10842_/A _09851_/X _14307_/C _10843_/X _09869_/B vssd1 vssd1 vccd1 vccd1
+ _10853_/A sky130_fd_sc_hd__a2111o_2
XANTENNA__19234__S0 _19275_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09627__B1 _09626_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16351_ _19362_/Q _16345_/X _16285_/X _16347_/X vssd1 vssd1 vccd1 vccd1 _19362_/D
+ sky130_fd_sc_hd__a22o_1
X_13563_ _20419_/Q _13559_/X _13475_/X _13561_/X vssd1 vssd1 vccd1 vccd1 _20419_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_13_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10775_ _10775_/A _10775_/B vssd1 vssd1 vccd1 vccd1 _10801_/A sky130_fd_sc_hd__or2_1
XANTENNA__18264__S _18904_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_212_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15302_ _15302_/A vssd1 vssd1 vccd1 vccd1 _15302_/X sky130_fd_sc_hd__buf_1
XFILLER_185_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12514_ _12523_/A vssd1 vssd1 vccd1 vccd1 _12520_/A sky130_fd_sc_hd__inv_2
X_19070_ _16733_/X _21140_/Q _19908_/D vssd1 vssd1 vccd1 vccd1 _19070_/X sky130_fd_sc_hd__mux2_1
XFILLER_158_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16282_ _19396_/Q _16276_/X _16281_/X _16279_/X vssd1 vssd1 vccd1 vccd1 _19396_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_200_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13494_ _13515_/A vssd1 vssd1 vccd1 vccd1 _13494_/X sky130_fd_sc_hd__buf_1
XFILLER_200_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18021_ _18021_/A vssd1 vssd1 vccd1 vccd1 _18021_/X sky130_fd_sc_hd__buf_1
Xclkbuf_leaf_5_HCLK clkbuf_opt_2_HCLK/A vssd1 vssd1 vccd1 vccd1 _19776_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_8_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15233_ _20486_/Q vssd1 vssd1 vccd1 vccd1 _15233_/Y sky130_fd_sc_hd__inv_2
X_12445_ _12445_/A vssd1 vssd1 vccd1 vccd1 _12445_/X sky130_fd_sc_hd__buf_2
XFILLER_60_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_repeater147_A _19058_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11510__A _20251_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15164_ _15088_/A _15088_/B _15089_/Y _15201_/B vssd1 vssd1 vccd1 vccd1 _20074_/D
+ sky130_fd_sc_hd__a211oi_2
X_12376_ _12376_/A _12376_/B _12376_/C vssd1 vssd1 vccd1 vccd1 _20960_/D sky130_fd_sc_hd__nor3_2
XFILLER_126_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19095__S _19870_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14115_ _14112_/Y _20286_/Q _20544_/Q _14083_/A _14114_/X vssd1 vssd1 vccd1 vccd1
+ _14120_/C sky130_fd_sc_hd__o221a_1
XFILLER_114_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11327_ _16683_/A vssd1 vssd1 vccd1 vccd1 _11327_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_153_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15095_ _20464_/Q _15090_/Y _15091_/Y _15092_/X _15094_/X vssd1 vssd1 vccd1 vccd1
+ _15110_/A sky130_fd_sc_hd__a221o_1
X_19972_ _20422_/CLK _19972_/D repeater184/X vssd1 vssd1 vccd1 vccd1 _19972_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_141_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18923_ _18922_/X _09745_/Y _18928_/S vssd1 vssd1 vccd1 vccd1 _18923_/X sky130_fd_sc_hd__mux2_1
XANTENNA__20930__CLK _20930_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14046_ _20282_/Q vssd1 vssd1 vccd1 vccd1 _14092_/A sky130_fd_sc_hd__inv_2
XFILLER_140_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11258_ _11300_/A vssd1 vssd1 vccd1 vccd1 _11543_/A sky130_fd_sc_hd__buf_1
XFILLER_79_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13437__A _13447_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10209_ _10207_/A _10207_/B _10177_/A _10207_/Y vssd1 vssd1 vccd1 vccd1 _21386_/D
+ sky130_fd_sc_hd__a211oi_2
X_18854_ _17079_/Y _12074_/Y _18908_/S vssd1 vssd1 vccd1 vccd1 _18854_/X sky130_fd_sc_hd__mux2_1
X_11189_ _15847_/A _11549_/A vssd1 vssd1 vccd1 vccd1 _16487_/A sky130_fd_sc_hd__or2_2
XFILLER_39_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15100__A1 _15097_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17805_ _17548_/X _17788_/X _17560_/X _17797_/X _17804_/X vssd1 vssd1 vccd1 vccd1
+ _17805_/Y sky130_fd_sc_hd__o221ai_4
XANTENNA__15100__B2 _15099_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21174__RESET_B repeater216/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15997_ _19535_/Q _15993_/X _15949_/X _15994_/X vssd1 vssd1 vccd1 vccd1 _19535_/D
+ sky130_fd_sc_hd__a22o_1
X_18785_ _18784_/X _14938_/Y _18907_/S vssd1 vssd1 vccd1 vccd1 _18785_/X sky130_fd_sc_hd__mux2_2
XANTENNA__16748__A _16758_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18439__S _18667_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14948_ _14936_/X _14948_/B _14948_/C _14948_/D vssd1 vssd1 vccd1 vccd1 _14949_/D
+ sky130_fd_sc_hd__and4b_1
XFILLER_94_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17736_ _12606_/A _17729_/X _17731_/X _17734_/X _17735_/X vssd1 vssd1 vccd1 vccd1
+ _17736_/X sky130_fd_sc_hd__o2111a_1
XFILLER_236_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_236_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15939__B1 _15891_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14879_ _14965_/A _14972_/A vssd1 vssd1 vccd1 vccd1 _14880_/B sky130_fd_sc_hd__or2_2
X_17667_ _19644_/Q vssd1 vssd1 vccd1 vccd1 _17667_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19406_ _19813_/CLK _19406_/D vssd1 vssd1 vccd1 vccd1 _19406_/Q sky130_fd_sc_hd__dfxtp_1
X_16618_ _16618_/A vssd1 vssd1 vccd1 vccd1 _16618_/Y sky130_fd_sc_hd__inv_2
XFILLER_211_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13414__A1 _20482_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19225__S0 _19275_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17598_ _19507_/Q vssd1 vssd1 vccd1 vccd1 _17598_/Y sky130_fd_sc_hd__inv_2
X_16549_ _19991_/Q vssd1 vssd1 vccd1 vccd1 _16553_/A sky130_fd_sc_hd__inv_2
X_19337_ _20142_/CLK _19337_/D vssd1 vssd1 vccd1 vccd1 _19337_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18174__S _18874_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19268_ _17118_/Y _17119_/Y _17120_/Y _17121_/Y _20130_/Q _20131_/Q vssd1 vssd1 vccd1
+ vccd1 _19268_/X sky130_fd_sc_hd__mux4_2
XFILLER_191_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18219_ _20843_/Q input1/X _18242_/S vssd1 vssd1 vccd1 vccd1 _18219_/X sky130_fd_sc_hd__mux2_1
X_19199_ _17765_/Y _17766_/Y _17767_/Y _17768_/Y _20130_/Q _20131_/Q vssd1 vssd1 vccd1
+ vccd1 _19199_/X sky130_fd_sc_hd__mux4_1
XFILLER_117_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18902__S _18902_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21230_ _21239_/CLK _21230_/D repeater249/X vssd1 vssd1 vccd1 vccd1 _21230_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_191_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21161_ _21162_/CLK _21161_/D repeater226/X vssd1 vssd1 vccd1 vccd1 _21161_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_131_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_161_HCLK_A clkbuf_opt_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20112_ _21433_/CLK _20112_/D repeater234/X vssd1 vssd1 vccd1 vccd1 _20112_/Q sky130_fd_sc_hd__dfrtp_1
X_09923_ _21435_/Q _21436_/Q _09924_/S vssd1 vssd1 vccd1 vccd1 _21436_/D sky130_fd_sc_hd__mux2_1
X_21092_ _21193_/CLK _21092_/D repeater226/X vssd1 vssd1 vccd1 vccd1 _21092_/Q sky130_fd_sc_hd__dfrtp_2
X_20043_ _20075_/CLK _20043_/D repeater276/X vssd1 vssd1 vccd1 vccd1 _20043_/Q sky130_fd_sc_hd__dfrtp_2
X_09854_ _21443_/Q vssd1 vssd1 vccd1 vccd1 _09857_/A sky130_fd_sc_hd__buf_1
XFILLER_59_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09785_ _14309_/A vssd1 vssd1 vccd1 vccd1 _14530_/C sky130_fd_sc_hd__inv_2
XFILLER_46_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18349__S _18885_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13102__B1 _12881_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19921__RESET_B repeater211/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20945_ _20946_/CLK _20945_/D repeater275/X vssd1 vssd1 vccd1 vccd1 _20945_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19216__S0 _21005_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20876_ _21459_/CLK _20876_/D repeater244/X vssd1 vssd1 vccd1 vccd1 _20876_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_81_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20826__RESET_B repeater251/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_241_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10560_ _10660_/A _10659_/A _10652_/A _10651_/A vssd1 vssd1 vccd1 vccd1 _10566_/C
+ sky130_fd_sc_hd__or4_4
XFILLER_128_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18812__S _18897_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10491_ _21281_/Q vssd1 vssd1 vccd1 vccd1 _10758_/A sky130_fd_sc_hd__inv_2
XFILLER_182_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12230_ _12429_/A _20520_/Q _20939_/Q _12229_/Y vssd1 vssd1 vccd1 vccd1 _12230_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_136_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21428_ _21429_/CLK _21428_/D repeater229/X vssd1 vssd1 vccd1 vccd1 _21428_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_30_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17936__B _17936_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12161_ _20351_/Q vssd1 vssd1 vccd1 vccd1 _12161_/Y sky130_fd_sc_hd__inv_2
X_21359_ _21367_/CLK _21359_/D repeater254/X vssd1 vssd1 vccd1 vccd1 _21359_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_2_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11112_ _11112_/A vssd1 vssd1 vccd1 vccd1 _11112_/X sky130_fd_sc_hd__buf_1
XFILLER_123_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12092_ _20962_/Q vssd1 vssd1 vccd1 vccd1 _12315_/A sky130_fd_sc_hd__inv_2
XANTENNA__13341__B1 _13277_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_20_HCLK_A clkbuf_4_3_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11043_ _19981_/Q _19980_/Q _17008_/A vssd1 vssd1 vccd1 vccd1 _16885_/B sky130_fd_sc_hd__or3_4
X_15920_ _15927_/A vssd1 vssd1 vccd1 vccd1 _15920_/X sky130_fd_sc_hd__buf_1
XFILLER_104_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_83_HCLK_A clkbuf_4_13_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_237_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15851_ _15857_/A vssd1 vssd1 vccd1 vccd1 _15851_/X sky130_fd_sc_hd__buf_1
XANTENNA__18259__S _18908_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14802_ _14791_/Y _14797_/A _20119_/Q _14796_/A vssd1 vssd1 vccd1 vccd1 _14803_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_218_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18570_ _18569_/X _10764_/A _18617_/S vssd1 vssd1 vccd1 vccd1 _18570_/X sky130_fd_sc_hd__mux2_2
X_15782_ _19637_/Q _15779_/X _15725_/X _15781_/X vssd1 vssd1 vccd1 vccd1 _19637_/D
+ sky130_fd_sc_hd__a22o_1
X_12994_ _20694_/Q _12983_/X _12993_/X _12987_/X vssd1 vssd1 vccd1 vccd1 _20694_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17521_ _19329_/Q vssd1 vssd1 vccd1 vccd1 _17521_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14733_ _14733_/A vssd1 vssd1 vccd1 vccd1 _14733_/X sky130_fd_sc_hd__buf_1
X_11945_ _11943_/X _11940_/B _11944_/Y _11917_/X _11936_/Y vssd1 vssd1 vccd1 vccd1
+ _11946_/A sky130_fd_sc_hd__o32a_1
XANTENNA_output114_A _17092_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_217_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17452_ _20400_/Q vssd1 vssd1 vccd1 vccd1 _17452_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19207__S0 _20130_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14664_ _14655_/Y _19124_/S _14660_/A _14663_/Y vssd1 vssd1 vccd1 vccd1 _14664_/X
+ sky130_fd_sc_hd__o211a_1
X_11876_ _21245_/Q _16592_/A vssd1 vssd1 vccd1 vccd1 _11877_/A sky130_fd_sc_hd__or2_2
XFILLER_220_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16403_ _19334_/Q _16399_/X _16340_/X _16400_/X vssd1 vssd1 vccd1 vccd1 _19334_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_221_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13615_ _20391_/Q _13613_/X _13550_/X _13614_/X vssd1 vssd1 vccd1 vccd1 _20391_/D
+ sky130_fd_sc_hd__a22o_1
X_10827_ _10827_/A vssd1 vssd1 vccd1 vccd1 _10827_/X sky130_fd_sc_hd__buf_2
X_17383_ _17377_/Y _17301_/A _11665_/Y _17378_/X _17382_/X vssd1 vssd1 vccd1 vccd1
+ _17383_/X sky130_fd_sc_hd__o221a_1
X_14595_ _14595_/A _14595_/B vssd1 vssd1 vccd1 vccd1 _14596_/A sky130_fd_sc_hd__or2_1
XFILLER_201_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19122_ _16484_/Y _14526_/Y _19124_/S vssd1 vssd1 vccd1 vccd1 _19122_/X sky130_fd_sc_hd__mux2_2
X_16334_ _16334_/A vssd1 vssd1 vccd1 vccd1 _16334_/X sky130_fd_sc_hd__buf_1
X_13546_ _20426_/Q _13537_/X _13545_/X _13541_/X vssd1 vssd1 vccd1 vccd1 _20426_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_186_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10758_ _10758_/A _10758_/B vssd1 vssd1 vccd1 vccd1 _10833_/A sky130_fd_sc_hd__or2_1
XFILLER_9_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19053_ _16771_/X _20816_/Q _19058_/S vssd1 vssd1 vccd1 vccd1 _19923_/D sky130_fd_sc_hd__mux2_1
XANTENNA__18007__B _18007_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16265_ _19405_/Q _16262_/X _16109_/X _16264_/X vssd1 vssd1 vccd1 vccd1 _19405_/D
+ sky130_fd_sc_hd__a22o_1
X_13477_ input51/X vssd1 vssd1 vccd1 vccd1 _13477_/X sky130_fd_sc_hd__clkbuf_2
X_10689_ _10657_/A _10657_/B _10685_/X _10687_/Y vssd1 vssd1 vccd1 vccd1 _21328_/D
+ sky130_fd_sc_hd__a211oi_4
XANTENNA__18722__S _18902_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16361__A3 _19889_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18004_ _18004_/A _18006_/B vssd1 vssd1 vccd1 vccd1 _18004_/Y sky130_fd_sc_hd__nor2_1
X_15216_ _20044_/Q _14970_/X _15214_/A _15160_/X vssd1 vssd1 vccd1 vccd1 _20044_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12907__B1 _12658_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12428_ _12428_/A _12451_/A vssd1 vssd1 vccd1 vccd1 _12429_/B sky130_fd_sc_hd__or2_2
XFILLER_173_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16196_ _21453_/Q vssd1 vssd1 vccd1 vccd1 _16196_/X sky130_fd_sc_hd__buf_1
Xclkbuf_leaf_106_HCLK clkbuf_4_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20944_/CLK sky130_fd_sc_hd__clkbuf_16
X_15147_ _20437_/Q _15128_/X _15145_/Y _20047_/Q _15146_/X vssd1 vssd1 vccd1 vccd1
+ _15157_/A sky130_fd_sc_hd__o221a_1
XFILLER_153_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12359_ _12359_/A vssd1 vssd1 vccd1 vccd1 _12359_/X sky130_fd_sc_hd__buf_1
XFILLER_99_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09645__A _12853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19955_ _21234_/CLK _19955_/D repeater188/X vssd1 vssd1 vccd1 vccd1 _19955_/Q sky130_fd_sc_hd__dfrtp_1
X_15078_ _15112_/A _15078_/B vssd1 vssd1 vccd1 vccd1 _15181_/A sky130_fd_sc_hd__or2_1
XANTENNA__21355__RESET_B repeater252/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18906_ _18905_/X _15136_/Y _18906_/S vssd1 vssd1 vccd1 vccd1 _18906_/X sky130_fd_sc_hd__mux2_2
XFILLER_68_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14029_ _20295_/Q _14033_/A _14026_/A _13965_/X vssd1 vssd1 vccd1 vccd1 _20295_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__17862__A _17862_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19886_ _20256_/CLK _19886_/D repeater217/X vssd1 vssd1 vccd1 vccd1 _19888_/D sky130_fd_sc_hd__dfstp_1
XFILLER_206_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18837_ _18845_/A0 _17283_/Y _18879_/S vssd1 vssd1 vccd1 vccd1 _18837_/X sky130_fd_sc_hd__mux2_1
XFILLER_121_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18169__S _18884_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18768_ _18767_/X _16895_/Y _18875_/S vssd1 vssd1 vccd1 vccd1 _18768_/X sky130_fd_sc_hd__mux2_2
XFILLER_48_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_222_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17719_ _17711_/Y _17301_/X _17714_/X _17718_/X vssd1 vssd1 vccd1 vccd1 _17719_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_82_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18699_ _18698_/X _12150_/Y _18909_/S vssd1 vssd1 vccd1 vccd1 _18699_/X sky130_fd_sc_hd__mux2_1
XFILLER_222_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20730_ _21375_/CLK _20730_/D repeater257/X vssd1 vssd1 vccd1 vccd1 _20730_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_223_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20661_ _20661_/CLK _20661_/D repeater261/X vssd1 vssd1 vccd1 vccd1 _20661_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_189_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20237__RESET_B repeater204/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20592_ _20592_/CLK _20592_/D repeater259/X vssd1 vssd1 vccd1 vccd1 _20592_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__10973__B _20887_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10621__B2 _10619_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18632__S _18669_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13571__B1 _13489_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21213_ _21255_/CLK _21213_/D repeater241/X vssd1 vssd1 vccd1 vccd1 _21213_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_144_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21144_ _21147_/CLK _21144_/D repeater215/X vssd1 vssd1 vccd1 vccd1 _21144_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_120_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13323__B1 _13166_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09906_ _20006_/Q vssd1 vssd1 vccd1 vccd1 _17020_/A sky130_fd_sc_hd__buf_1
X_21075_ _21087_/CLK _21075_/D repeater228/X vssd1 vssd1 vccd1 vccd1 _21075_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_99_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20026_ _21486_/CLK _20026_/D repeater209/X vssd1 vssd1 vccd1 vccd1 _20026_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_76_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18262__A0 _18848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09837_ _21446_/Q vssd1 vssd1 vccd1 vccd1 _16163_/A sky130_fd_sc_hd__buf_1
XFILLER_19_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09768_ _09768_/A _09768_/B _09768_/C _09768_/D vssd1 vssd1 vccd1 vccd1 _09769_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_100_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09699_ _21464_/Q _09690_/X _09698_/X _09694_/X vssd1 vssd1 vccd1 vccd1 _21464_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18807__S _18841_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_215_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11730_ _21063_/Q _11727_/X _11680_/X _11729_/X vssd1 vssd1 vccd1 vccd1 _21063_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20928_ _20930_/CLK _20928_/D repeater266/X vssd1 vssd1 vccd1 vccd1 _20928_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11661_ _11502_/X _11652_/X _19112_/S _11659_/Y _21094_/Q vssd1 vssd1 vccd1 vccd1
+ _21094_/D sky130_fd_sc_hd__a32o_1
XPHY_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20859_ _21445_/CLK _20859_/D repeater243/X vssd1 vssd1 vccd1 vccd1 _20859_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13400_ _20492_/Q _13398_/X _13277_/X _13399_/X vssd1 vssd1 vccd1 vccd1 _20492_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10612_ _10569_/A _20760_/Q _21311_/Q _10611_/Y vssd1 vssd1 vccd1 vccd1 _10612_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14380_ _20237_/Q _20236_/Q _14380_/C vssd1 vssd1 vccd1 vccd1 _14467_/A sky130_fd_sc_hd__and3_1
XFILLER_167_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_129_HCLK clkbuf_4_4_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _21242_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11592_ _21122_/Q _11592_/B vssd1 vssd1 vccd1 vccd1 _11592_/Y sky130_fd_sc_hd__nand2_1
XPHY_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13331_ _13351_/A vssd1 vssd1 vccd1 vccd1 _13331_/X sky130_fd_sc_hd__buf_1
XFILLER_183_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10543_ _10543_/A vssd1 vssd1 vccd1 vccd1 _10704_/A sky130_fd_sc_hd__clkbuf_2
Xclkbuf_2_1_0_HCLK clkbuf_2_1_0_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_3_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XPHY_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18542__S _18907_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16050_ _16056_/A vssd1 vssd1 vccd1 vccd1 _16057_/A sky130_fd_sc_hd__inv_2
XANTENNA_input75_A scl_i_S4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13262_ _17080_/A _13262_/B vssd1 vssd1 vccd1 vccd1 _13299_/A sky130_fd_sc_hd__or2_2
XFILLER_155_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10474_ _21292_/Q vssd1 vssd1 vccd1 vccd1 _10768_/A sky130_fd_sc_hd__inv_2
X_15001_ _15001_/A _15015_/A vssd1 vssd1 vccd1 vccd1 _15002_/B sky130_fd_sc_hd__or2_2
XANTENNA__21131__CLK _21134_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13562__B1 _13560_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12213_ _12395_/A _20526_/Q _20921_/Q _12209_/Y _12212_/Y vssd1 vssd1 vccd1 vccd1
+ _12232_/A sky130_fd_sc_hd__o221a_1
XANTENNA__17828__B1 _17838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13193_ _13225_/A vssd1 vssd1 vccd1 vccd1 _13227_/A sky130_fd_sc_hd__inv_2
XANTENNA__10376__B1 _10375_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12144_ _12144_/A _12144_/B _12144_/C _12144_/D vssd1 vssd1 vccd1 vccd1 _12145_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_2_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15303__B2 _18962_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12117__B2 _17895_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13314__B1 _13313_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19740_ _19765_/CLK _19740_/D vssd1 vssd1 vccd1 vccd1 _19740_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12075_ _20955_/Q vssd1 vssd1 vccd1 vccd1 _12309_/A sky130_fd_sc_hd__inv_2
X_16952_ _16950_/Y _16951_/Y _16939_/X vssd1 vssd1 vccd1 vccd1 _16952_/X sky130_fd_sc_hd__o21a_1
XFILLER_49_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21281__CLK _21342_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18253__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15903_ _16093_/A _16150_/B _16377_/C vssd1 vssd1 vccd1 vccd1 _15911_/A sky130_fd_sc_hd__or3_4
X_11026_ _19951_/Q _19950_/Q vssd1 vssd1 vccd1 vccd1 _16886_/A sky130_fd_sc_hd__or2_1
X_19671_ _19821_/CLK _19671_/D vssd1 vssd1 vccd1 vccd1 _19671_/Q sky130_fd_sc_hd__dfxtp_1
X_16883_ _16971_/A vssd1 vssd1 vccd1 vccd1 _16894_/A sky130_fd_sc_hd__buf_2
XFILLER_237_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18622_ _18621_/X _10781_/A _18898_/S vssd1 vssd1 vccd1 vccd1 _18622_/X sky130_fd_sc_hd__mux2_1
XFILLER_66_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15834_ _15841_/A vssd1 vssd1 vccd1 vccd1 _15834_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_64_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20748__RESET_B repeater207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18553_ _17079_/Y _12127_/Y _18908_/S vssd1 vssd1 vccd1 vccd1 _18553_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12977_ _12891_/X _20699_/Q _12977_/S vssd1 vssd1 vccd1 vccd1 _20699_/D sky130_fd_sc_hd__mux2_1
X_15765_ _19643_/Q _15757_/X _15764_/X _15760_/X vssd1 vssd1 vccd1 vccd1 _19643_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_205_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18717__S _18879_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17504_ _19589_/Q _19588_/Q _19587_/Q _19586_/Q vssd1 vssd1 vccd1 vccd1 _17504_/Y
+ sky130_fd_sc_hd__nor4_2
X_14716_ _20152_/Q _14711_/X _13586_/X _14712_/X vssd1 vssd1 vccd1 vccd1 _20152_/D
+ sky130_fd_sc_hd__a22o_1
X_11928_ _21008_/Q vssd1 vssd1 vccd1 vccd1 _11928_/Y sky130_fd_sc_hd__inv_2
XFILLER_233_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18484_ _17079_/Y _15269_/Y _18908_/S vssd1 vssd1 vccd1 vccd1 _18484_/X sky130_fd_sc_hd__mux2_1
X_15696_ _15696_/A vssd1 vssd1 vccd1 vccd1 _15696_/X sky130_fd_sc_hd__buf_1
XFILLER_72_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14647_ _14570_/A _14570_/B _14639_/X _14645_/Y vssd1 vssd1 vccd1 vccd1 _20180_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_32_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17435_ _19577_/Q vssd1 vssd1 vccd1 vccd1 _17435_/Y sky130_fd_sc_hd__inv_2
X_11859_ _11859_/A vssd1 vssd1 vccd1 vccd1 _11860_/B sky130_fd_sc_hd__inv_2
XFILLER_177_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18018__A _18018_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20330__RESET_B repeater190/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14578_ _14578_/A _14630_/A vssd1 vssd1 vccd1 vccd1 _14579_/B sky130_fd_sc_hd__or2_1
XFILLER_32_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17366_ _20141_/Q vssd1 vssd1 vccd1 vccd1 _17366_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19105_ _16665_/X _21073_/Q _19870_/D vssd1 vssd1 vccd1 vccd1 _19105_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10603__B2 _10602_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16317_ _19379_/Q _16312_/X _16237_/X _16314_/X vssd1 vssd1 vccd1 vccd1 _19379_/D
+ sky130_fd_sc_hd__a22o_1
X_13529_ _13181_/C _13528_/X _13524_/Y vssd1 vssd1 vccd1 vccd1 _20431_/D sky130_fd_sc_hd__a21oi_1
X_17297_ _17289_/Y _17290_/X _17291_/Y _17292_/X _17296_/X vssd1 vssd1 vccd1 vccd1
+ _17297_/X sky130_fd_sc_hd__o221a_1
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18452__S _18884_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19036_ _16846_/X _20833_/Q _19046_/S vssd1 vssd1 vccd1 vccd1 _19940_/D sky130_fd_sc_hd__mux2_1
X_16248_ _16255_/A vssd1 vssd1 vccd1 vccd1 _16248_/X sky130_fd_sc_hd__buf_1
XFILLER_133_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput103 _18105_/Y vssd1 vssd1 vccd1 vccd1 HRDATA[31] sky130_fd_sc_hd__clkbuf_2
XFILLER_114_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput114 _17092_/X vssd1 vssd1 vccd1 vccd1 IRQ[11] sky130_fd_sc_hd__clkbuf_2
X_16179_ _16179_/A _16405_/B _16194_/C vssd1 vssd1 vccd1 vccd1 _16187_/A sky130_fd_sc_hd__or3_4
XFILLER_127_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput125 _17088_/X vssd1 vssd1 vccd1 vccd1 IRQ[7] sky130_fd_sc_hd__clkbuf_2
Xoutput136 _20982_/Q vssd1 vssd1 vccd1 vccd1 pwm_S6 sky130_fd_sc_hd__clkbuf_2
XANTENNA__18492__A0 _18491_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13305__B1 _13146_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19938_ _20159_/CLK _19938_/D repeater269/X vssd1 vssd1 vccd1 vccd1 _19938_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_102_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19869_ _21183_/CLK _19869_/D repeater216/X vssd1 vssd1 vccd1 vccd1 _19869_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_96_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09622_ _09672_/A vssd1 vssd1 vccd1 vccd1 _09677_/A sky130_fd_sc_hd__inv_2
XANTENNA__13625__A _13625_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18627__S _18841_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20418__RESET_B repeater187/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__21004__CLK _21009_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_212_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20713_ _20724_/CLK _20713_/D repeater254/X vssd1 vssd1 vccd1 vccd1 _20713_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_196_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20071__RESET_B repeater276/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20644_ _20657_/CLK _20644_/D repeater198/X vssd1 vssd1 vccd1 vccd1 _20644_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_149_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20000__RESET_B repeater225/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18362__S _18787_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20575_ _20947_/CLK _20575_/D repeater266/X vssd1 vssd1 vccd1 vccd1 _20575_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_165_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__21277__RESET_B repeater205/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13544__B1 _13543_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10190_ _10190_/A vssd1 vssd1 vccd1 vccd1 _10190_/Y sky130_fd_sc_hd__inv_2
XFILLER_160_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21127_ _21134_/CLK _21127_/D repeater192/X vssd1 vssd1 vccd1 vccd1 _21127_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_160_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21058_ _21147_/CLK _21058_/D repeater212/X vssd1 vssd1 vccd1 vccd1 _21058_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_59_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12900_ _12934_/A vssd1 vssd1 vccd1 vccd1 _12924_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__13535__A _13657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20009_ _21438_/CLK _20009_/D repeater240/X vssd1 vssd1 vccd1 vccd1 _20009_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_247_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13880_ _13971_/D _14006_/A vssd1 vssd1 vccd1 vccd1 _13881_/B sky130_fd_sc_hd__or2_1
XFILLER_234_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17994__C1 _17993_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12831_ _20765_/Q _12829_/X _12663_/X _12830_/X vssd1 vssd1 vccd1 vccd1 _20765_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_36_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18537__S _18787_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15550_ _15663_/A vssd1 vssd1 vccd1 vccd1 _15550_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_215_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12762_ _20803_/Q _12757_/X _12656_/X _12760_/X vssd1 vssd1 vccd1 vccd1 _20803_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_199_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14501_ _14501_/A _14510_/A vssd1 vssd1 vccd1 vccd1 _14502_/B sky130_fd_sc_hd__or2_1
XFILLER_202_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11713_ _11720_/A vssd1 vssd1 vccd1 vccd1 _11713_/X sky130_fd_sc_hd__buf_1
XPHY_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15481_ _15481_/A vssd1 vssd1 vccd1 vccd1 _15481_/X sky130_fd_sc_hd__buf_1
X_12693_ _12707_/A vssd1 vssd1 vccd1 vccd1 _12693_/X sky130_fd_sc_hd__buf_1
XFILLER_230_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13270__A input61/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14432_ _21485_/Q _14333_/A _21484_/Q _14460_/A vssd1 vssd1 vccd1 vccd1 _14432_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17220_ _18930_/X _17854_/A _18910_/X _17219_/X vssd1 vssd1 vccd1 vccd1 _17220_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11644_ _18978_/X _11640_/X _21102_/Q _11642_/X vssd1 vssd1 vccd1 vccd1 _21102_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17151_ _17378_/A vssd1 vssd1 vccd1 vccd1 _17151_/X sky130_fd_sc_hd__buf_1
XPHY_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14363_ _14517_/A _14463_/A vssd1 vssd1 vccd1 vccd1 _14364_/B sky130_fd_sc_hd__or2_2
XPHY_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11575_ _19881_/Q vssd1 vssd1 vccd1 vccd1 _16546_/A sky130_fd_sc_hd__buf_1
Xinput16 HADDR[23] vssd1 vssd1 vccd1 vccd1 input16/X sky130_fd_sc_hd__buf_1
XANTENNA__18272__S _18908_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput27 HADDR[4] vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_hd__buf_1
XPHY_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16102_ _16102_/A vssd1 vssd1 vccd1 vccd1 _16102_/X sky130_fd_sc_hd__buf_1
XPHY_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput38 HWDATA[0] vssd1 vssd1 vccd1 vccd1 input38/X sky130_fd_sc_hd__buf_6
X_13314_ _20538_/Q _13307_/X _13313_/X _13308_/X vssd1 vssd1 vccd1 vccd1 _20538_/D
+ sky130_fd_sc_hd__a22o_1
X_10526_ _21343_/Q _10824_/A _10421_/Y vssd1 vssd1 vccd1 vccd1 _21343_/D sky130_fd_sc_hd__o21a_1
Xinput49 HWDATA[1] vssd1 vssd1 vccd1 vccd1 input49/X sky130_fd_sc_hd__buf_2
X_17082_ _17808_/A vssd1 vssd1 vccd1 vccd1 _18902_/S sky130_fd_sc_hd__clkinv_16
X_14294_ _14293_/X _14280_/X _14783_/B vssd1 vssd1 vccd1 vccd1 _14294_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16033_ _19518_/Q _16028_/X _15776_/X _16029_/X vssd1 vssd1 vccd1 vccd1 _19518_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_115_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13245_ _14264_/A vssd1 vssd1 vccd1 vccd1 _13245_/X sky130_fd_sc_hd__buf_2
X_10457_ _10779_/A _20692_/Q _21288_/Q _10456_/Y vssd1 vssd1 vccd1 vccd1 _10457_/X
+ sky130_fd_sc_hd__o22a_1
X_13176_ _13717_/B vssd1 vssd1 vccd1 vccd1 _16525_/B sky130_fd_sc_hd__buf_1
X_10388_ _10388_/A vssd1 vssd1 vccd1 vccd1 _10388_/Y sky130_fd_sc_hd__inv_2
XFILLER_123_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12127_ _20375_/Q vssd1 vssd1 vccd1 vccd1 _12127_/Y sky130_fd_sc_hd__inv_2
XFILLER_97_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17984_ _20417_/Q _18007_/B vssd1 vssd1 vccd1 vccd1 _17984_/Y sky130_fd_sc_hd__nand2_1
XFILLER_78_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19723_ _20327_/CLK _19723_/D vssd1 vssd1 vccd1 vccd1 _19723_/Q sky130_fd_sc_hd__dfxtp_1
X_12058_ _12311_/A _20371_/Q _20957_/Q _12057_/Y vssd1 vssd1 vccd1 vccd1 _12058_/X
+ sky130_fd_sc_hd__o22a_1
X_16935_ _16956_/A _16935_/B vssd1 vssd1 vccd1 vccd1 _16935_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__13445__A input63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11009_ _11909_/B vssd1 vssd1 vccd1 vccd1 _15374_/B sky130_fd_sc_hd__buf_1
X_19654_ _19821_/CLK _19654_/D vssd1 vssd1 vccd1 vccd1 _19654_/Q sky130_fd_sc_hd__dfxtp_1
X_16866_ _16865_/Y _16862_/A _19945_/Q _16862_/Y _16779_/A vssd1 vssd1 vccd1 vccd1
+ _16866_/X sky130_fd_sc_hd__o221a_1
XANTENNA__16788__B1 _16779_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18605_ _18604_/X _14403_/Y _18669_/S vssd1 vssd1 vccd1 vccd1 _18605_/X sky130_fd_sc_hd__mux2_1
X_15817_ _15824_/A vssd1 vssd1 vccd1 vccd1 _15817_/X sky130_fd_sc_hd__clkbuf_2
X_19585_ _21021_/CLK _19585_/D vssd1 vssd1 vccd1 vccd1 _19585_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18529__A1 _20193_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16797_ _19930_/Q vssd1 vssd1 vccd1 vccd1 _16797_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18447__S _18885_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20511__RESET_B repeater267/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18536_ _18535_/X _16815_/A _18667_/S vssd1 vssd1 vccd1 vccd1 _18536_/X sky130_fd_sc_hd__mux2_1
XFILLER_179_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15748_ _19651_/Q _15743_/X _15733_/X _15745_/X vssd1 vssd1 vccd1 vccd1 _19651_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18467_ _18845_/A0 _13764_/Y _18896_/S vssd1 vssd1 vccd1 vccd1 _18467_/X sky130_fd_sc_hd__mux2_1
XANTENNA__14276__A _20124_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15679_ _19683_/Q _15674_/X _15663_/X _15676_/X vssd1 vssd1 vccd1 vccd1 _19683_/D
+ sky130_fd_sc_hd__a22o_1
X_17418_ _19721_/Q vssd1 vssd1 vccd1 vccd1 _17418_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18398_ _18397_/X _10761_/A _18880_/S vssd1 vssd1 vccd1 vccd1 _18398_/X sky130_fd_sc_hd__mux2_1
XFILLER_193_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12577__A1 _20887_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17349_ _19600_/Q _17369_/B vssd1 vssd1 vccd1 vccd1 _17349_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__18182__S _18669_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20360_ _20951_/CLK _20360_/D repeater272/X vssd1 vssd1 vccd1 vccd1 _20360_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__21370__RESET_B repeater255/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19019_ _16916_/X _20404_/Q _19019_/S vssd1 vssd1 vccd1 vccd1 _19957_/D sky130_fd_sc_hd__mux2_1
X_20291_ _20293_/CLK _20291_/D repeater263/X vssd1 vssd1 vccd1 vccd1 _20291_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_228_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18910__S _18910_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09605_ _17204_/A _13048_/A vssd1 vssd1 vccd1 vccd1 _13110_/A sky130_fd_sc_hd__or2_2
XFILLER_28_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18357__S _18850_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18940__A1 _21136_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21458__RESET_B repeater245/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20627_ _20697_/CLK _20627_/D repeater193/X vssd1 vssd1 vccd1 vccd1 _20627_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11360_ _11409_/A _11411_/A vssd1 vssd1 vccd1 vccd1 _11782_/B sky130_fd_sc_hd__nor2_1
XFILLER_20_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20558_ _20592_/CLK _20558_/D repeater260/X vssd1 vssd1 vccd1 vccd1 _20558_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_137_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18105__B _18105_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13517__B1 _13449_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10311_ _21346_/Q _10308_/Y _10262_/A _20705_/Q _10310_/X vssd1 vssd1 vccd1 vccd1
+ _10311_/X sky130_fd_sc_hd__a221o_1
XFILLER_125_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11291_ _16568_/A _18970_/X vssd1 vssd1 vccd1 vccd1 _12504_/A sky130_fd_sc_hd__or2b_1
XANTENNA__21040__RESET_B repeater247/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18820__S _18908_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20489_ _20495_/CLK _20489_/D repeater274/X vssd1 vssd1 vccd1 vccd1 _20489_/Q sky130_fd_sc_hd__dfrtp_4
X_13030_ _13311_/A vssd1 vssd1 vccd1 vccd1 _13030_/X sky130_fd_sc_hd__clkbuf_4
X_10242_ _21361_/Q vssd1 vssd1 vccd1 vccd1 _10276_/A sky130_fd_sc_hd__inv_2
XANTENNA__17944__B _17944_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10173_ _21403_/Q _10172_/Y _10034_/B _10172_/A _10166_/X vssd1 vssd1 vccd1 vccd1
+ _21403_/D sky130_fd_sc_hd__o221a_1
XFILLER_239_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18208__A0 _17079_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input38_A HWDATA[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14981_ _14981_/A vssd1 vssd1 vccd1 vccd1 _14981_/Y sky130_fd_sc_hd__inv_2
XANTENNA__10889__A _12550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16720_ _16720_/A _18933_/X vssd1 vssd1 vccd1 vccd1 _19903_/D sky130_fd_sc_hd__and2_1
XANTENNA__17960__A _18045_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13265__A input62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13932_ _20654_/Q vssd1 vssd1 vccd1 vccd1 _13932_/Y sky130_fd_sc_hd__inv_2
XFILLER_170_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16651_ _19860_/Q _15294_/B _15295_/B vssd1 vssd1 vccd1 vccd1 _16651_/X sky130_fd_sc_hd__a21bo_1
XFILLER_74_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13863_ _20293_/Q vssd1 vssd1 vccd1 vccd1 _13865_/B sky130_fd_sc_hd__inv_2
XANTENNA__18267__S _18904_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12814_ _12809_/X _16779_/A _12814_/S vssd1 vssd1 vccd1 vccd1 _20771_/D sky130_fd_sc_hd__mux2_1
X_15602_ _19722_/Q _15596_/X _15477_/X _15598_/X vssd1 vssd1 vccd1 vccd1 _19722_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_138_HCLK_A clkbuf_4_12_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19370_ _19706_/CLK _19370_/D vssd1 vssd1 vccd1 vccd1 _19370_/Q sky130_fd_sc_hd__dfxtp_1
X_16582_ _16551_/Y _16737_/A _19992_/Q vssd1 vssd1 vccd1 vccd1 _16583_/B sky130_fd_sc_hd__a21oi_1
X_13794_ _20179_/Q vssd1 vssd1 vccd1 vccd1 _14569_/A sky130_fd_sc_hd__inv_2
XFILLER_15_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18321_ _18320_/X _12268_/Y _18910_/S vssd1 vssd1 vccd1 vccd1 _18321_/X sky130_fd_sc_hd__mux2_1
X_15533_ _19756_/Q _15529_/X _15454_/X _15531_/X vssd1 vssd1 vccd1 vccd1 _19756_/D
+ sky130_fd_sc_hd__a22o_1
X_12745_ _14686_/A _12740_/B _12738_/B _12751_/B vssd1 vssd1 vccd1 vccd1 _12745_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_31_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_repeater177_A _18666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18252_ _18037_/Y _16986_/Y _18680_/S vssd1 vssd1 vccd1 vccd1 _18252_/X sky130_fd_sc_hd__mux2_2
X_15464_ _19782_/Q _15459_/X _15431_/X _15460_/X vssd1 vssd1 vccd1 vccd1 _19782_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12676_ _20833_/Q _12672_/X _09621_/X _12674_/X vssd1 vssd1 vccd1 vccd1 _20833_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14415_ _21478_/Q vssd1 vssd1 vccd1 vccd1 _14415_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19098__S _19870_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17203_ _18048_/A vssd1 vssd1 vccd1 vccd1 _17203_/X sky130_fd_sc_hd__buf_2
XPHY_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11627_ _11638_/A _11632_/A _21106_/Q vssd1 vssd1 vccd1 vccd1 _11628_/A sky130_fd_sc_hd__or3b_1
XPHY_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18183_ _18182_/X _20184_/Q _18748_/S vssd1 vssd1 vccd1 vccd1 _18183_/X sky130_fd_sc_hd__mux2_2
X_15395_ _21014_/Q vssd1 vssd1 vccd1 vccd1 _15655_/B sky130_fd_sc_hd__buf_1
XPHY_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14346_ _20632_/Q vssd1 vssd1 vccd1 vccd1 _14517_/A sky130_fd_sc_hd__inv_2
X_17134_ _21072_/Q vssd1 vssd1 vccd1 vccd1 _17134_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18695__A0 _17079_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11558_ input64/X vssd1 vssd1 vccd1 vccd1 _16332_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_155_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13508__B1 _13506_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17065_ _12006_/A _19288_/Q _12008_/A vssd1 vssd1 vccd1 vccd1 _17066_/B sky130_fd_sc_hd__o21a_1
XFILLER_195_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10509_ _10774_/A _20687_/Q _10505_/X _20675_/Q _10508_/X vssd1 vssd1 vccd1 vccd1
+ _10522_/B sky130_fd_sc_hd__o221a_1
XFILLER_143_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14277_ _20122_/Q vssd1 vssd1 vccd1 vccd1 _14279_/A sky130_fd_sc_hd__inv_2
XFILLER_155_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12344__A _12359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18730__S _18910_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11489_ _13383_/A _17140_/B _11489_/C vssd1 vssd1 vccd1 vccd1 _15847_/B sky130_fd_sc_hd__or3_4
X_16016_ _16016_/A vssd1 vssd1 vccd1 vccd1 _16016_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_170_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13228_ _13249_/A vssd1 vssd1 vccd1 vccd1 _13228_/X sky130_fd_sc_hd__buf_1
X_13159_ _13167_/A vssd1 vssd1 vccd1 vccd1 _13159_/X sky130_fd_sc_hd__buf_1
XFILLER_3_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20763__RESET_B repeater211/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17967_ _20830_/Q vssd1 vssd1 vccd1 vccd1 _17967_/Y sky130_fd_sc_hd__inv_2
X_19706_ _19706_/CLK _19706_/D vssd1 vssd1 vccd1 vccd1 _19706_/Q sky130_fd_sc_hd__dfxtp_1
X_16918_ _16971_/A vssd1 vssd1 vccd1 vccd1 _16956_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_214_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17898_ _17898_/A _17898_/B vssd1 vssd1 vccd1 vccd1 _17898_/Y sky130_fd_sc_hd__nor2_1
XFILLER_238_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19637_ _20142_/CLK _19637_/D vssd1 vssd1 vccd1 vccd1 _19637_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_226_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16849_ _19941_/Q _16844_/Y _16847_/Y _16844_/A _16848_/X vssd1 vssd1 vccd1 vccd1
+ _16849_/X sky130_fd_sc_hd__o221a_1
XANTENNA__18177__S _18897_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_214_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19568_ _19706_/CLK _19568_/D vssd1 vssd1 vccd1 vccd1 _19568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18519_ _18518_/X _13923_/Y _18849_/S vssd1 vssd1 vccd1 vccd1 _18519_/X sky130_fd_sc_hd__mux2_1
XFILLER_222_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19499_ _20327_/CLK _19499_/D vssd1 vssd1 vccd1 vccd1 _19499_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_230_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19270__S1 _20131_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18905__S _18908_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21461_ _21461_/CLK _21461_/D repeater245/X vssd1 vssd1 vccd1 vccd1 _21461_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18686__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20412_ _20413_/CLK _20412_/D repeater184/X vssd1 vssd1 vccd1 vccd1 _20412_/Q sky130_fd_sc_hd__dfrtp_1
X_21392_ _21401_/CLK _21392_/D repeater253/X vssd1 vssd1 vccd1 vccd1 _21392_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_190_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20343_ _20949_/CLK _20343_/D repeater269/X vssd1 vssd1 vccd1 vccd1 _20343_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__18640__S _18908_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18438__A0 _18848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20274_ _20724_/CLK _20274_/D repeater263/X vssd1 vssd1 vccd1 vccd1 _20274_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_248_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21342__CLK _21342_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20433__RESET_B repeater278/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_229_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13813__A _20602_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10860_ _11654_/A _17195_/A vssd1 vssd1 vccd1 vccd1 _10908_/B sky130_fd_sc_hd__or2_2
XFILLER_231_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10791_ _21306_/Q _10790_/Y _10787_/X _10783_/B vssd1 vssd1 vccd1 vccd1 _21306_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19261__S1 _20133_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18815__S _18849_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12530_ _11270_/B _12527_/X _11272_/B _12528_/X vssd1 vssd1 vccd1 vccd1 _20912_/D
+ sky130_fd_sc_hd__o22ai_1
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_235_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12461_ _12461_/A vssd1 vssd1 vccd1 vccd1 _12461_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21221__RESET_B repeater235/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14200_ _14087_/A _14087_/B _14198_/Y _14193_/X vssd1 vssd1 vccd1 vccd1 _20277_/D
+ sky130_fd_sc_hd__a211oi_2
X_11412_ _16595_/B _11412_/B _11412_/C _11412_/D vssd1 vssd1 vccd1 vccd1 _11413_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_184_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15180_ _15129_/X _15080_/B _15176_/Y _15179_/X vssd1 vssd1 vccd1 vccd1 _20066_/D
+ sky130_fd_sc_hd__a211oi_2
X_12392_ _20950_/Q _12445_/A _12359_/A _12389_/A vssd1 vssd1 vccd1 vccd1 _20950_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_165_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14131_ _20558_/Q _14097_/A _14130_/Y _20287_/Q vssd1 vssd1 vccd1 vccd1 _14131_/X
+ sky130_fd_sc_hd__o22a_1
X_11343_ _21176_/Q vssd1 vssd1 vccd1 vccd1 _11347_/B sky130_fd_sc_hd__inv_2
XFILLER_152_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12164__A _20347_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18550__S _18884_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18429__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14062_ _20266_/Q vssd1 vssd1 vccd1 vccd1 _14077_/A sky130_fd_sc_hd__inv_2
X_11274_ _11299_/C _11294_/A _11283_/C _12505_/B vssd1 vssd1 vccd1 vccd1 _11541_/C
+ sky130_fd_sc_hd__or4_4
XFILLER_4_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20037__SET_B repeater216/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13013_ _13013_/A vssd1 vssd1 vccd1 vccd1 _13013_/X sky130_fd_sc_hd__buf_1
XFILLER_79_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10225_ _10041_/B _10224_/A _21378_/Q _10227_/A _10166_/X vssd1 vssd1 vccd1 vccd1
+ _21378_/D sky130_fd_sc_hd__o221a_1
X_18870_ _18869_/X _19266_/X _18930_/S vssd1 vssd1 vccd1 vccd1 _18870_/X sky130_fd_sc_hd__mux2_1
X_17821_ _17821_/A vssd1 vssd1 vccd1 vccd1 _17952_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_121_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10156_ _10156_/A _10187_/A vssd1 vssd1 vccd1 vccd1 _10157_/B sky130_fd_sc_hd__or2_2
XANTENNA_output144_A _21042_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20174__RESET_B repeater249/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17752_ _19299_/Q vssd1 vssd1 vccd1 vccd1 _17752_/Y sky130_fd_sc_hd__inv_2
XFILLER_248_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14964_ _20497_/Q _14964_/B vssd1 vssd1 vccd1 vccd1 _14964_/X sky130_fd_sc_hd__or2_1
X_10087_ _21407_/Q _10086_/Y _10079_/Y _20804_/Q vssd1 vssd1 vccd1 vccd1 _10087_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_236_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20103__RESET_B repeater259/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16703_ _16709_/A _18941_/X vssd1 vssd1 vccd1 vccd1 _19895_/D sky130_fd_sc_hd__and2_1
XFILLER_47_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17404__B2 _17326_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13915_ _20658_/Q vssd1 vssd1 vccd1 vccd1 _13915_/Y sky130_fd_sc_hd__inv_2
XFILLER_208_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17683_ _18708_/X _17703_/B vssd1 vssd1 vccd1 vccd1 _17683_/X sky130_fd_sc_hd__and2_1
X_14895_ _20581_/Q vssd1 vssd1 vccd1 vccd1 _14895_/Y sky130_fd_sc_hd__inv_2
X_19422_ _19521_/CLK _19422_/D vssd1 vssd1 vccd1 vccd1 _19422_/Q sky130_fd_sc_hd__dfxtp_1
X_16634_ _16634_/A _18962_/X vssd1 vssd1 vccd1 vccd1 _19852_/D sky130_fd_sc_hd__nor2_1
X_13846_ _20314_/Q vssd1 vssd1 vccd1 vccd1 _13974_/C sky130_fd_sc_hd__inv_2
XFILLER_16_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19353_ _19626_/CLK _19353_/D vssd1 vssd1 vccd1 vccd1 _19353_/Q sky130_fd_sc_hd__dfxtp_1
X_16565_ _16744_/A _16738_/B _16539_/X _16564_/X vssd1 vssd1 vccd1 vccd1 _19995_/D
+ sky130_fd_sc_hd__o31ai_1
XFILLER_204_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13777_ _20627_/Q vssd1 vssd1 vccd1 vccd1 _13777_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21309__RESET_B repeater211/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18725__S _18908_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19252__S1 _21004_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10989_ _21017_/Q vssd1 vssd1 vccd1 vccd1 _10991_/A sky130_fd_sc_hd__inv_2
XANTENNA__11243__A _19910_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18304_ _18303_/X _18015_/Y _18906_/S vssd1 vssd1 vccd1 vccd1 _18304_/X sky130_fd_sc_hd__mux2_1
XFILLER_204_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15516_ _15516_/A vssd1 vssd1 vccd1 vccd1 _15516_/X sky130_fd_sc_hd__buf_1
X_12728_ _13535_/B _13108_/B vssd1 vssd1 vccd1 vccd1 _12729_/S sky130_fd_sc_hd__or2_1
X_19284_ _19693_/Q _19381_/Q _19677_/Q _19669_/Q _19285_/S0 _21017_/Q vssd1 vssd1
+ vccd1 vccd1 _19284_/X sky130_fd_sc_hd__mux4_2
X_16496_ _19875_/Q vssd1 vssd1 vccd1 vccd1 _16496_/Y sky130_fd_sc_hd__inv_2
XFILLER_188_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18235_ _20859_/Q input8/X _18236_/S vssd1 vssd1 vccd1 vccd1 _18235_/X sky130_fd_sc_hd__mux2_1
XFILLER_230_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15447_ _20127_/Q vssd1 vssd1 vccd1 vccd1 _15624_/B sky130_fd_sc_hd__buf_1
XPHY_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12659_ _20840_/Q _12650_/X _12658_/X _12654_/X vssd1 vssd1 vccd1 vccd1 _20840_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18668__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09648__A input42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18166_ _18845_/A0 _10518_/Y _18896_/S vssd1 vssd1 vccd1 vccd1 _18166_/X sky130_fd_sc_hd__mux2_1
X_15378_ _15657_/A vssd1 vssd1 vccd1 vccd1 _15378_/X sky130_fd_sc_hd__buf_1
XFILLER_172_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17117_ _19341_/Q vssd1 vssd1 vccd1 vccd1 _17117_/Y sky130_fd_sc_hd__inv_2
X_14329_ _20234_/Q vssd1 vssd1 vccd1 vccd1 _14465_/A sky130_fd_sc_hd__inv_2
XFILLER_171_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18460__S _18898_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18097_ _17925_/A _18097_/B _18097_/C vssd1 vssd1 vccd1 vccd1 _18097_/Y sky130_fd_sc_hd__nand3b_4
XFILLER_128_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17048_ _17054_/B _17048_/B vssd1 vssd1 vccd1 vccd1 _19871_/D sky130_fd_sc_hd__nor2_1
XFILLER_131_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09870_ _09870_/A _09872_/A vssd1 vssd1 vccd1 vccd1 _09870_/X sky130_fd_sc_hd__or2_1
Xrepeater200 repeater206/X vssd1 vssd1 vccd1 vccd1 repeater200/X sky130_fd_sc_hd__buf_8
X_18999_ _17002_/X _20424_/Q _19026_/S vssd1 vssd1 vccd1 vccd1 _19977_/D sky130_fd_sc_hd__mux2_1
XFILLER_57_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater211 repeater212/X vssd1 vssd1 vccd1 vccd1 repeater211/X sky130_fd_sc_hd__clkbuf_8
XFILLER_97_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater222 repeater224/X vssd1 vssd1 vccd1 vccd1 repeater222/X sky130_fd_sc_hd__buf_8
Xrepeater233 repeater234/X vssd1 vssd1 vccd1 vccd1 repeater233/X sky130_fd_sc_hd__buf_6
XFILLER_245_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater244 repeater245/X vssd1 vssd1 vccd1 vccd1 repeater244/X sky130_fd_sc_hd__buf_6
XFILLER_39_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater255 repeater256/X vssd1 vssd1 vccd1 vccd1 repeater255/X sky130_fd_sc_hd__buf_8
XFILLER_54_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater266 repeater267/X vssd1 vssd1 vccd1 vccd1 repeater266/X sky130_fd_sc_hd__buf_8
X_20961_ _20971_/CLK _20961_/D repeater187/X vssd1 vssd1 vccd1 vccd1 _20961_/Q sky130_fd_sc_hd__dfrtp_2
Xrepeater277 repeater278/X vssd1 vssd1 vccd1 vccd1 repeater277/X sky130_fd_sc_hd__clkbuf_8
XPHY_4409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11691__A1 _21083_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20892_ _21338_/CLK _20892_/D repeater221/X vssd1 vssd1 vccd1 vccd1 _20892_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_3719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_20_HCLK clkbuf_4_3_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _21438_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_clkbuf_leaf_121_HCLK_A clkbuf_opt_3_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_241_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18635__S _18891_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19243__S1 _21004_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_222_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18659__A0 _17281_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14393__B1 _21477_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21444_ _21444_/CLK _21444_/D repeater243/X vssd1 vssd1 vccd1 vccd1 _21444_/Q sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_162_HCLK clkbuf_opt_0_HCLK/A vssd1 vssd1 vccd1 vccd1 _21462_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_5_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21375_ _21375_/CLK _21375_/D repeater257/X vssd1 vssd1 vccd1 vccd1 _21375_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18370__S _18841_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20685__RESET_B repeater208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20326_ _20326_/CLK _20326_/D repeater250/X vssd1 vssd1 vccd1 vccd1 _20326_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__19755__CLK _19765_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20257_ _20908_/CLK _20257_/D repeater217/X vssd1 vssd1 vccd1 vccd1 _20257_/Q sky130_fd_sc_hd__dfstp_1
X_10010_ _21415_/Q _17032_/A vssd1 vssd1 vccd1 vccd1 _10010_/Y sky130_fd_sc_hd__nand2_1
X_20188_ _21485_/CLK _20188_/D repeater200/X vssd1 vssd1 vccd1 vccd1 _20188_/Q sky130_fd_sc_hd__dfrtp_1
X_09999_ _20016_/Q vssd1 vssd1 vccd1 vccd1 _09999_/X sky130_fd_sc_hd__buf_1
XFILLER_77_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11961_ _13185_/B vssd1 vssd1 vccd1 vccd1 _11961_/Y sky130_fd_sc_hd__inv_2
XFILLER_217_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14563__A1_N _20133_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13700_ _13708_/A vssd1 vssd1 vccd1 vccd1 _13700_/X sky130_fd_sc_hd__buf_1
XFILLER_72_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13543__A input61/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10912_ _12750_/A _20701_/Q vssd1 vssd1 vccd1 vccd1 _12742_/A sky130_fd_sc_hd__or2_2
XFILLER_217_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14680_ _14680_/A _14682_/A vssd1 vssd1 vccd1 vccd1 _14680_/X sky130_fd_sc_hd__or2_1
XFILLER_45_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11892_ _11881_/A _11881_/B _11881_/Y _11889_/X vssd1 vssd1 vccd1 vccd1 _11892_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__21473__RESET_B repeater204/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13631_ _13631_/A vssd1 vssd1 vccd1 vccd1 _13651_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_44_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10843_ _20034_/Q _10843_/B _10843_/C vssd1 vssd1 vccd1 vccd1 _10843_/X sky130_fd_sc_hd__and3_1
XANTENNA__13262__B _13262_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18545__S _18775_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19234__S1 _21004_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21402__RESET_B repeater255/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13562_ _20420_/Q _13559_/X _13560_/X _13561_/X vssd1 vssd1 vccd1 vccd1 _20420_/D
+ sky130_fd_sc_hd__a22o_1
X_16350_ _19363_/Q _16345_/X _16283_/X _16347_/X vssd1 vssd1 vccd1 vccd1 _19363_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19868__RESET_B repeater202/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10774_ _10774_/A _10804_/A vssd1 vssd1 vccd1 vccd1 _10775_/B sky130_fd_sc_hd__or2_2
X_15301_ _15305_/A vssd1 vssd1 vccd1 vccd1 _18962_/S sky130_fd_sc_hd__clkbuf_8
X_12513_ _11316_/X _12511_/Y _12512_/Y vssd1 vssd1 vccd1 vccd1 _12523_/A sky130_fd_sc_hd__o21ai_2
XFILLER_212_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_43_HCLK_A _20004_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16281_ _20330_/Q vssd1 vssd1 vccd1 vccd1 _16281_/X sky130_fd_sc_hd__clkbuf_2
X_13493_ _13493_/A vssd1 vssd1 vccd1 vccd1 _13515_/A sky130_fd_sc_hd__clkbuf_2
X_18020_ _18020_/A vssd1 vssd1 vccd1 vccd1 _18020_/X sky130_fd_sc_hd__buf_1
X_15232_ _15232_/A _15232_/B _15232_/C _15232_/D vssd1 vssd1 vccd1 vccd1 _15232_/X
+ sky130_fd_sc_hd__and4_1
X_12444_ _12432_/A _12443_/A _20943_/Q _12443_/Y _12411_/X vssd1 vssd1 vccd1 vccd1
+ _20943_/D sky130_fd_sc_hd__o221a_1
XANTENNA__11198__B1 _10900_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15163_ _15193_/A vssd1 vssd1 vccd1 vccd1 _15201_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_3_0_0_HCLK_A clkbuf_3_1_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12375_ _12139_/X _12377_/A _12081_/X vssd1 vssd1 vccd1 vccd1 _12376_/C sky130_fd_sc_hd__o21a_1
XFILLER_125_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17322__B1 _18853_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14114_ _20559_/Q _14098_/A _18031_/A _20283_/Q vssd1 vssd1 vccd1 vccd1 _14114_/X
+ sky130_fd_sc_hd__o22a_1
X_11326_ _11371_/A vssd1 vssd1 vccd1 vccd1 _16683_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__17873__A1 _18570_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15094_ _20441_/Q _15093_/X _20450_/Q _15075_/A vssd1 vssd1 vccd1 vccd1 _15094_/X
+ sky130_fd_sc_hd__a22o_1
X_19971_ _20422_/CLK _19971_/D repeater184/X vssd1 vssd1 vccd1 vccd1 _19971_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_181_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14687__A1 _10985_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18922_ _18921_/X _18112_/A _18927_/S vssd1 vssd1 vccd1 vccd1 _18922_/X sky130_fd_sc_hd__mux2_1
X_14045_ _20283_/Q vssd1 vssd1 vccd1 vccd1 _14093_/A sky130_fd_sc_hd__inv_2
XANTENNA__13718__A _13727_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11257_ _20917_/Q vssd1 vssd1 vccd1 vccd1 _11300_/A sky130_fd_sc_hd__buf_1
XFILLER_125_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12698__B1 _12697_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19170__S0 _19280_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10208_ _21387_/Q _10207_/Y _10166_/A _10149_/B vssd1 vssd1 vccd1 vccd1 _21387_/D
+ sky130_fd_sc_hd__o211a_1
X_18853_ _18852_/X _14897_/Y _18907_/S vssd1 vssd1 vccd1 vccd1 _18853_/X sky130_fd_sc_hd__mux2_2
X_11188_ _11199_/A _17133_/B _11200_/A vssd1 vssd1 vccd1 vccd1 _11549_/A sky130_fd_sc_hd__or3_4
XFILLER_39_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15636__B1 _15590_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17804_ _12606_/A _17798_/X _17800_/X _17802_/X _17803_/X vssd1 vssd1 vccd1 vccd1
+ _17804_/X sky130_fd_sc_hd__o2111a_1
XFILLER_39_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10139_ _10260_/B vssd1 vssd1 vccd1 vccd1 _10183_/A sky130_fd_sc_hd__buf_1
X_18784_ _18783_/X _15145_/Y _18784_/S vssd1 vssd1 vccd1 vccd1 _18784_/X sky130_fd_sc_hd__mux2_2
XFILLER_227_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15996_ _19536_/Q _15993_/X _15947_/X _15994_/X vssd1 vssd1 vccd1 vccd1 _19536_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_94_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09931__A _16342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_43_HCLK _20004_/CLK vssd1 vssd1 vccd1 vccd1 _21055_/CLK sky130_fd_sc_hd__clkbuf_16
X_17735_ _18682_/X _17856_/A _18691_/X _17480_/X vssd1 vssd1 vccd1 vccd1 _17735_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_48_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14947_ _20592_/Q _14881_/B _14896_/Y _20086_/Q _14946_/X vssd1 vssd1 vccd1 vccd1
+ _14948_/D sky130_fd_sc_hd__o221a_1
XFILLER_75_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17666_ _19500_/Q vssd1 vssd1 vccd1 vccd1 _17666_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12870__B1 _12548_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14878_ _14965_/B _14878_/B vssd1 vssd1 vccd1 vccd1 _14972_/A sky130_fd_sc_hd__or2_1
X_19405_ _21011_/CLK _19405_/D vssd1 vssd1 vccd1 vccd1 _19405_/Q sky130_fd_sc_hd__dfxtp_1
X_16617_ _16617_/A _16617_/B vssd1 vssd1 vccd1 vccd1 _16617_/X sky130_fd_sc_hd__or2_1
XFILLER_90_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13829_ _13824_/Y _20182_/Q _13825_/Y _20192_/Q _13828_/X vssd1 vssd1 vccd1 vccd1
+ _13836_/C sky130_fd_sc_hd__o221a_1
XFILLER_90_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19225__S1 _21004_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18455__S _18885_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17597_ _19387_/Q vssd1 vssd1 vccd1 vccd1 _17597_/Y sky130_fd_sc_hd__inv_2
XFILLER_211_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19336_ _20241_/CLK _19336_/D vssd1 vssd1 vccd1 vccd1 _19336_/Q sky130_fd_sc_hd__dfxtp_1
X_16548_ _16548_/A vssd1 vssd1 vccd1 vccd1 _16566_/A sky130_fd_sc_hd__inv_2
XFILLER_188_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19267_ _17114_/Y _17115_/Y _17116_/Y _17117_/Y _20130_/Q _20131_/Q vssd1 vssd1 vccd1
+ vccd1 _19267_/X sky130_fd_sc_hd__mux4_1
X_16479_ _16479_/A vssd1 vssd1 vccd1 vccd1 _18930_/S sky130_fd_sc_hd__clkinv_8
X_18218_ _12566_/X _18218_/A1 _19986_/D vssd1 vssd1 vccd1 vccd1 _19985_/D sky130_fd_sc_hd__mux2_2
XFILLER_176_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19198_ _17761_/Y _17762_/Y _17763_/Y _17764_/Y _20130_/Q _20131_/Q vssd1 vssd1 vccd1
+ vccd1 _19198_/X sky130_fd_sc_hd__mux4_2
XFILLER_191_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18149_ _18148_/X _20281_/Q _18904_/S vssd1 vssd1 vccd1 vccd1 _18149_/X sky130_fd_sc_hd__mux2_1
XANTENNA__18190__S _18669_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14127__B1 _20541_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21160_ _21162_/CLK _21160_/D repeater227/X vssd1 vssd1 vccd1 vccd1 _21160_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_132_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20096__RESET_B repeater259/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20111_ _21433_/CLK _20111_/D repeater234/X vssd1 vssd1 vccd1 vccd1 _20111_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_104_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09922_ _21436_/Q _21437_/Q _09924_/S vssd1 vssd1 vccd1 vccd1 _21437_/D sky130_fd_sc_hd__mux2_1
XFILLER_236_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21091_ _21424_/CLK _21091_/D repeater230/X vssd1 vssd1 vccd1 vccd1 _21091_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12689__B1 _09641_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20042_ _20042_/CLK _20042_/D repeater219/X vssd1 vssd1 vccd1 vccd1 _20042_/Q sky130_fd_sc_hd__dfstp_1
X_09853_ _21444_/Q vssd1 vssd1 vccd1 vccd1 _09853_/X sky130_fd_sc_hd__buf_1
XFILLER_59_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09784_ _21459_/Q vssd1 vssd1 vccd1 vccd1 _16619_/A sky130_fd_sc_hd__buf_1
XFILLER_100_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20944_ _20944_/CLK _20944_/D repeater275/X vssd1 vssd1 vccd1 vccd1 _20944_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_4239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18365__S _18617_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20875_ _21459_/CLK _20875_/D repeater244/X vssd1 vssd1 vccd1 vccd1 _20875_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19216__S1 _21006_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_241_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19961__RESET_B repeater185/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_241_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12707__A _12707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20866__RESET_B repeater247/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10490_ _20676_/Q vssd1 vssd1 vccd1 vccd1 _10490_/Y sky130_fd_sc_hd__inv_2
XFILLER_194_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21427_ _21429_/CLK _21427_/D repeater229/X vssd1 vssd1 vccd1 vccd1 _21427_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_163_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12160_ _20354_/Q vssd1 vssd1 vccd1 vccd1 _12160_/Y sky130_fd_sc_hd__inv_2
XFILLER_123_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21358_ _21367_/CLK _21358_/D repeater254/X vssd1 vssd1 vccd1 vccd1 _21358_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_146_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11111_ _11111_/A vssd1 vssd1 vccd1 vccd1 _21228_/D sky130_fd_sc_hd__inv_2
XFILLER_107_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13538__A input62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20309_ _20316_/CLK _20309_/D repeater197/X vssd1 vssd1 vccd1 vccd1 _20309_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_146_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12091_ _20966_/Q _20380_/Q _12089_/X _12090_/Y vssd1 vssd1 vccd1 vccd1 _12103_/A
+ sky130_fd_sc_hd__o22a_1
X_21289_ _21357_/CLK _21289_/D repeater209/X vssd1 vssd1 vccd1 vccd1 _21289_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_150_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19152__S0 _19285_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11042_ _19979_/Q _19978_/Q _17004_/A vssd1 vssd1 vccd1 vccd1 _17008_/A sky130_fd_sc_hd__or3_4
Xclkbuf_leaf_66_HCLK clkbuf_4_11_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20915_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__19870__D _19870_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15850_ _15856_/A vssd1 vssd1 vccd1 vccd1 _15857_/A sky130_fd_sc_hd__inv_2
XFILLER_237_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15094__A1 _20441_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14801_ _14795_/Y _19125_/S _14800_/Y vssd1 vssd1 vccd1 vccd1 _14803_/A sky130_fd_sc_hd__o21ai_1
XANTENNA_input20_A HADDR[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15781_ _15789_/A vssd1 vssd1 vccd1 vccd1 _15781_/X sky130_fd_sc_hd__buf_1
XFILLER_18_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12993_ input58/X vssd1 vssd1 vccd1 vccd1 _12993_/X sky130_fd_sc_hd__buf_2
XFILLER_57_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17520_ _19353_/Q vssd1 vssd1 vccd1 vccd1 _17520_/Y sky130_fd_sc_hd__inv_2
XFILLER_245_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10458__A2 _20696_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14732_ _14732_/A vssd1 vssd1 vccd1 vccd1 _14733_/A sky130_fd_sc_hd__inv_2
XANTENNA__12852__B1 _12849_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11944_ _11944_/A _11944_/B vssd1 vssd1 vccd1 vccd1 _11944_/Y sky130_fd_sc_hd__nor2_1
XFILLER_233_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17451_ _20814_/Q vssd1 vssd1 vccd1 vccd1 _17451_/Y sky130_fd_sc_hd__inv_2
XFILLER_233_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14663_ _14663_/A _14663_/B vssd1 vssd1 vccd1 vccd1 _14663_/Y sky130_fd_sc_hd__nand2_1
X_11875_ _16594_/A _11875_/B vssd1 vssd1 vccd1 vccd1 _16592_/A sky130_fd_sc_hd__or2_1
XANTENNA__19207__S1 _20131_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output107_A _17737_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_233_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16402_ _19335_/Q _16399_/X _16338_/X _16400_/X vssd1 vssd1 vccd1 vccd1 _19335_/D
+ sky130_fd_sc_hd__a22o_1
X_10826_ _10505_/X _10825_/A _21286_/Q _10825_/Y _10787_/X vssd1 vssd1 vccd1 vccd1
+ _21286_/D sky130_fd_sc_hd__o221a_1
X_13614_ _13626_/A vssd1 vssd1 vccd1 vccd1 _13614_/X sky130_fd_sc_hd__buf_1
X_17382_ _17379_/Y _17292_/A _17380_/Y _17381_/X vssd1 vssd1 vccd1 vccd1 _17382_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12604__B1 _18222_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14594_ _14594_/A _14602_/A vssd1 vssd1 vccd1 vccd1 _14595_/B sky130_fd_sc_hd__or2_2
XFILLER_13_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19121_ _19124_/S _16483_/Y _19123_/S vssd1 vssd1 vccd1 vccd1 _19121_/X sky130_fd_sc_hd__mux2_1
X_16333_ _19370_/Q _16326_/X _16332_/X _16328_/X vssd1 vssd1 vccd1 vccd1 _19370_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_201_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10757_ _10757_/A _10836_/A vssd1 vssd1 vccd1 vccd1 _10758_/B sky130_fd_sc_hd__or2_2
X_13545_ input59/X vssd1 vssd1 vccd1 vccd1 _13545_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_40_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19052_ _16775_/X _20817_/Q _19058_/S vssd1 vssd1 vccd1 vccd1 _19924_/D sky130_fd_sc_hd__mux2_1
X_13476_ _20455_/Q _13472_/X _13475_/X _13473_/X vssd1 vssd1 vccd1 vccd1 _20455_/D
+ sky130_fd_sc_hd__a22o_1
X_16264_ _16270_/A vssd1 vssd1 vccd1 vccd1 _16264_/X sky130_fd_sc_hd__buf_1
X_10688_ _21329_/Q _10687_/Y _10680_/X _10659_/B vssd1 vssd1 vccd1 vccd1 _21329_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_187_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20536__RESET_B repeater267/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12907__A1 _20732_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18003_ _18003_/A _18006_/B vssd1 vssd1 vccd1 vccd1 _18003_/Y sky130_fd_sc_hd__nor2_1
X_15215_ _20045_/Q _15214_/Y _15061_/B _15177_/X vssd1 vssd1 vccd1 vccd1 _20045_/D
+ sky130_fd_sc_hd__o211a_1
X_12427_ _12427_/A _12427_/B vssd1 vssd1 vccd1 vccd1 _12451_/A sky130_fd_sc_hd__or2_1
X_16195_ _16206_/A vssd1 vssd1 vccd1 vccd1 _16195_/X sky130_fd_sc_hd__buf_1
XANTENNA__17846__A1 _18593_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15146_ _20445_/Q _15070_/A _20453_/Q _15112_/X vssd1 vssd1 vccd1 vccd1 _15146_/X
+ sky130_fd_sc_hd__o22a_1
X_12358_ _12358_/A vssd1 vssd1 vccd1 vccd1 _12358_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17846__B2 _17203_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11309_ _20908_/Q vssd1 vssd1 vccd1 vccd1 _11310_/B sky130_fd_sc_hd__inv_2
X_15077_ _15077_/A _15184_/A vssd1 vssd1 vccd1 vccd1 _15078_/B sky130_fd_sc_hd__or2_2
X_19954_ _20809_/CLK _19954_/D repeater188/X vssd1 vssd1 vccd1 vccd1 _19954_/Q sky130_fd_sc_hd__dfrtp_1
X_12289_ _20527_/Q vssd1 vssd1 vccd1 vccd1 _12289_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19143__S0 _19285_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18905_ _17174_/Y _15218_/Y _18908_/S vssd1 vssd1 vccd1 vccd1 _18905_/X sky130_fd_sc_hd__mux2_1
X_14028_ _14028_/A vssd1 vssd1 vccd1 vccd1 _14033_/A sky130_fd_sc_hd__inv_2
X_19885_ _21338_/CLK _19885_/D repeater221/X vssd1 vssd1 vccd1 vccd1 _19885_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_141_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18836_ _18835_/X _16889_/A _18875_/S vssd1 vssd1 vccd1 vccd1 _18836_/X sky130_fd_sc_hd__mux2_2
XANTENNA__15663__A _15663_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18767_ _17281_/X _17452_/Y _18835_/S vssd1 vssd1 vccd1 vccd1 _18767_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13096__B1 _12957_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15979_ _15979_/A vssd1 vssd1 vccd1 vccd1 _15979_/X sky130_fd_sc_hd__buf_1
XANTENNA__21324__RESET_B repeater204/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17718_ _17715_/Y _11678_/A _16628_/A _17553_/X _17717_/X vssd1 vssd1 vccd1 vccd1
+ _17718_/X sky130_fd_sc_hd__o221a_1
XFILLER_222_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12843__B1 _09630_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18698_ _17079_/Y _12107_/Y _18908_/S vssd1 vssd1 vccd1 vccd1 _18698_/X sky130_fd_sc_hd__mux2_1
X_17649_ _17648_/Y _17639_/X _17062_/Y _17162_/B vssd1 vssd1 vccd1 vccd1 _17649_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_90_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18185__S _18904_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20660_ _20661_/CLK _20660_/D repeater261/X vssd1 vssd1 vccd1 vccd1 _20660_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_195_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19319_ _19961_/CLK _19319_/D vssd1 vssd1 vccd1 vccd1 _19319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20591_ _20592_/CLK _20591_/D repeater260/X vssd1 vssd1 vccd1 vccd1 _20591_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_31_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10621__A2 _10618_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21212_ _21401_/CLK _21212_/D repeater241/X vssd1 vssd1 vccd1 vccd1 _21212_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_117_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_89_HCLK clkbuf_4_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _21367_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_172_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21143_ _21191_/CLK _21143_/D repeater192/X vssd1 vssd1 vccd1 vccd1 _21143_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_116_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19134__S0 _19285_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09905_ _09902_/Y _17021_/A _21254_/Q _09904_/A vssd1 vssd1 vccd1 vccd1 _09905_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_120_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21074_ _21424_/CLK _21074_/D repeater229/X vssd1 vssd1 vccd1 vccd1 _21074_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_58_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20025_ _21486_/CLK _20025_/D repeater209/X vssd1 vssd1 vccd1 vccd1 _20025_/Q sky130_fd_sc_hd__dfrtp_2
X_09836_ _15881_/A _09827_/X _09835_/X _09829_/X vssd1 vssd1 vccd1 vccd1 _21447_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_219_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09767_ _21232_/Q _09762_/Y _11113_/A _20144_/Q _09766_/X vssd1 vssd1 vccd1 vccd1
+ _09768_/D sky130_fd_sc_hd__o221a_1
XFILLER_86_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12834__B1 _12670_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09698_ _10898_/A vssd1 vssd1 vccd1 vccd1 _09698_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_215_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19943__CLK _20930_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20927_ _20929_/CLK _20927_/D repeater267/X vssd1 vssd1 vccd1 vccd1 _20927_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_4069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_230_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11660_ _11486_/X _11652_/X _19112_/S _21095_/Q _11659_/Y vssd1 vssd1 vccd1 vccd1
+ _21095_/D sky130_fd_sc_hd__a32o_1
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20858_ _21445_/CLK _20858_/D repeater243/X vssd1 vssd1 vccd1 vccd1 _20858_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20920__CLK _20930_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10611_ _20739_/Q vssd1 vssd1 vccd1 vccd1 _10611_/Y sky130_fd_sc_hd__inv_2
XPHY_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11591_ _11591_/A _11591_/B vssd1 vssd1 vccd1 vccd1 _11592_/B sky130_fd_sc_hd__and2_1
XPHY_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20789_ _21374_/CLK _20789_/D repeater253/X vssd1 vssd1 vccd1 vccd1 _20789_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13330_ _13357_/A vssd1 vssd1 vccd1 vccd1 _13351_/A sky130_fd_sc_hd__buf_1
XPHY_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10542_ _21316_/Q vssd1 vssd1 vccd1 vccd1 _10543_/A sky130_fd_sc_hd__inv_2
XPHY_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10612__A2 _20760_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13261_ _13261_/A vssd1 vssd1 vccd1 vccd1 _17080_/A sky130_fd_sc_hd__buf_2
XFILLER_183_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10473_ _20683_/Q vssd1 vssd1 vccd1 vccd1 _17942_/A sky130_fd_sc_hd__inv_2
XANTENNA__13011__B1 _12922_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12212_ _12470_/A _20502_/Q _12424_/A _20515_/Q vssd1 vssd1 vccd1 vccd1 _12212_/Y
+ sky130_fd_sc_hd__a22oi_1
X_15000_ _15000_/A _15017_/A vssd1 vssd1 vccd1 vccd1 _15015_/A sky130_fd_sc_hd__or2_1
XFILLER_136_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17828__B2 _17819_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13192_ _13215_/A vssd1 vssd1 vccd1 vccd1 _13192_/X sky130_fd_sc_hd__buf_1
XANTENNA_input68_A HWDATA[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12143_ _20952_/Q _12137_/Y _12139_/X _20373_/Q _12142_/X vssd1 vssd1 vccd1 vccd1
+ _12144_/D sky130_fd_sc_hd__o221a_1
XANTENNA__17963__A _18048_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13314__A1 _20538_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16951_ _16951_/A _16951_/B vssd1 vssd1 vccd1 vccd1 _16951_/Y sky130_fd_sc_hd__nor2_1
X_12074_ _20365_/Q vssd1 vssd1 vccd1 vccd1 _12074_/Y sky130_fd_sc_hd__inv_2
XFILLER_150_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11025_ _19975_/Q _19974_/Q vssd1 vssd1 vccd1 vccd1 _11041_/C sky130_fd_sc_hd__or2_1
X_15902_ _16484_/B _15902_/B vssd1 vssd1 vccd1 vccd1 _16377_/C sky130_fd_sc_hd__or2_2
X_19670_ _19821_/CLK _19670_/D vssd1 vssd1 vccd1 vccd1 _19670_/Q sky130_fd_sc_hd__dfxtp_1
X_16882_ _16984_/A vssd1 vssd1 vccd1 vccd1 _16971_/A sky130_fd_sc_hd__inv_2
X_18621_ _18620_/X _10631_/Y _18897_/S vssd1 vssd1 vccd1 vccd1 _18621_/X sky130_fd_sc_hd__mux2_1
XFILLER_77_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15833_ _16093_/A _15833_/B _16194_/C vssd1 vssd1 vccd1 vccd1 _15841_/A sky130_fd_sc_hd__or3_4
XANTENNA__11516__A _16340_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18552_ _18551_/X _10270_/A _18841_/S vssd1 vssd1 vccd1 vccd1 _18552_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12825__B1 _12651_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15764_ _15764_/A vssd1 vssd1 vccd1 vccd1 _15764_/X sky130_fd_sc_hd__buf_1
X_12976_ _17087_/A _12981_/A vssd1 vssd1 vccd1 vccd1 _12977_/S sky130_fd_sc_hd__or2_1
XFILLER_61_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17503_ _21023_/Q _17425_/A _17348_/X _17501_/Y vssd1 vssd1 vccd1 vccd1 _17503_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_17_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14715_ _20153_/Q _14711_/X _13584_/X _14712_/X vssd1 vssd1 vccd1 vccd1 _20153_/D
+ sky130_fd_sc_hd__a22o_1
X_11927_ _11916_/Y _11917_/X _11165_/X _11926_/X vssd1 vssd1 vccd1 vccd1 _21011_/D
+ sky130_fd_sc_hd__o22ai_1
X_18483_ _18482_/X _14081_/A _18904_/S vssd1 vssd1 vccd1 vccd1 _18483_/X sky130_fd_sc_hd__mux2_1
X_15695_ _19674_/Q _15688_/X _15694_/X _15690_/X vssd1 vssd1 vccd1 vccd1 _19674_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17434_ _19593_/Q vssd1 vssd1 vccd1 vccd1 _17434_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17203__A _18048_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14646_ _20181_/Q _14645_/Y _14642_/X _14572_/B vssd1 vssd1 vccd1 vccd1 _20181_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_60_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11858_ _11858_/A vssd1 vssd1 vccd1 vccd1 _21029_/D sky130_fd_sc_hd__inv_2
XFILLER_32_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20717__RESET_B repeater254/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10809_ _10827_/A vssd1 vssd1 vccd1 vccd1 _10809_/X sky130_fd_sc_hd__buf_2
X_17365_ _19464_/Q vssd1 vssd1 vccd1 vccd1 _17365_/Y sky130_fd_sc_hd__inv_2
X_11789_ _21041_/Q _11418_/X _11396_/X vssd1 vssd1 vccd1 vccd1 _21041_/D sky130_fd_sc_hd__o21a_1
X_14577_ _14577_/A _14577_/B vssd1 vssd1 vccd1 vccd1 _14630_/A sky130_fd_sc_hd__or2_1
XFILLER_159_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18733__S _18928_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13250__B1 _13166_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19104_ _16666_/X _21074_/Q _19870_/D vssd1 vssd1 vccd1 vccd1 _19104_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16316_ _19380_/Q _16312_/X _16235_/X _16314_/X vssd1 vssd1 vccd1 vccd1 _19380_/D
+ sky130_fd_sc_hd__a22o_1
X_13528_ _13528_/A _13530_/A _13528_/C vssd1 vssd1 vccd1 vccd1 _13528_/X sky130_fd_sc_hd__or3_1
X_17296_ _17293_/Y _17141_/A _17294_/Y _17295_/X vssd1 vssd1 vccd1 vccd1 _17296_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_174_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20370__RESET_B repeater187/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19035_ _16849_/X _20834_/Q _19046_/S vssd1 vssd1 vccd1 vccd1 _19941_/D sky130_fd_sc_hd__mux2_1
XANTENNA__13002__B1 _13001_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16247_ _16247_/A _16344_/B _16261_/C vssd1 vssd1 vccd1 vccd1 _16255_/A sky130_fd_sc_hd__or3_4
X_13459_ _13491_/A vssd1 vssd1 vccd1 vccd1 _13493_/A sky130_fd_sc_hd__inv_2
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput104 _17483_/Y vssd1 vssd1 vccd1 vccd1 HRDATA[3] sky130_fd_sc_hd__clkbuf_2
Xoutput115 _18117_/LO vssd1 vssd1 vccd1 vccd1 IRQ[12] sky130_fd_sc_hd__clkbuf_2
X_16178_ _19446_/Q _16173_/X _16163_/X _16174_/X vssd1 vssd1 vccd1 vccd1 _19446_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_154_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput126 _17089_/X vssd1 vssd1 vccd1 vccd1 IRQ[8] sky130_fd_sc_hd__clkbuf_2
Xoutput137 _20043_/Q vssd1 vssd1 vccd1 vccd1 pwm_S7 sky130_fd_sc_hd__clkbuf_2
XFILLER_141_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15129_ _15129_/A vssd1 vssd1 vccd1 vccd1 _15129_/X sky130_fd_sc_hd__buf_1
X_19937_ _20159_/CLK _19937_/D repeater251/X vssd1 vssd1 vccd1 vccd1 _19937_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_68_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19868_ _20256_/CLK input77/X repeater202/X vssd1 vssd1 vccd1 vccd1 _19869_/D sky130_fd_sc_hd__dfrtp_1
XFILLER_229_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12810__A _12815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09621_ input52/X vssd1 vssd1 vccd1 vccd1 _09621_/X sky130_fd_sc_hd__buf_4
XFILLER_28_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18819_ _18818_/X _14909_/Y _18907_/S vssd1 vssd1 vccd1 vccd1 _18819_/X sky130_fd_sc_hd__mux2_2
XANTENNA__13069__B1 _12918_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19799_ _19820_/CLK _19799_/D vssd1 vssd1 vccd1 vccd1 _19799_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_244_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18908__S _18908_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_237_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12816__A0 _12809_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16007__B1 _16006_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_4_3_0_HCLK_A clkbuf_4_3_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20712_ _21366_/CLK _20712_/D repeater254/X vssd1 vssd1 vccd1 vccd1 _20712_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_197_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20458__RESET_B repeater276/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20643_ _20657_/CLK _20643_/D repeater198/X vssd1 vssd1 vccd1 vccd1 _20643_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_177_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18643__S _18884_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20574_ _20946_/CLK _20574_/D repeater275/X vssd1 vssd1 vccd1 vccd1 _20574_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11555__B1 _10884_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17783__A _21087_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21126_ _21185_/CLK _21126_/D repeater223/X vssd1 vssd1 vccd1 vccd1 _21126_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_133_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21057_ _21147_/CLK _21057_/D repeater215/X vssd1 vssd1 vccd1 vccd1 _21057_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__12720__A _12898_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20008_ _21223_/CLK _20008_/D repeater238/X vssd1 vssd1 vccd1 vccd1 _20008_/Q sky130_fd_sc_hd__dfrtp_1
X_09819_ _15869_/A _09813_/X _09818_/X _09815_/X vssd1 vssd1 vccd1 vccd1 _21452_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18818__S _18906_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12830_ _12842_/A vssd1 vssd1 vccd1 vccd1 _12830_/X sky130_fd_sc_hd__buf_1
XANTENNA__12807__B1 _11741_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12761_ _20804_/Q _12757_/X _12651_/X _12760_/X vssd1 vssd1 vccd1 vccd1 _20804_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14500_ _14500_/A _14500_/B vssd1 vssd1 vccd1 vccd1 _14510_/A sky130_fd_sc_hd__or2_1
XFILLER_199_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13551__A _13567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20881__RESET_B repeater243/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11712_ _14256_/A _15312_/D vssd1 vssd1 vccd1 vccd1 _11720_/A sky130_fd_sc_hd__or2_2
XPHY_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15480_ _15769_/A vssd1 vssd1 vccd1 vccd1 _15480_/X sky130_fd_sc_hd__clkbuf_2
X_12692_ _20823_/Q _12686_/X _09652_/X _12688_/X vssd1 vssd1 vccd1 vccd1 _20823_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_199_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20199__RESET_B repeater193/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14431_ _21475_/Q vssd1 vssd1 vccd1 vccd1 _14431_/Y sky130_fd_sc_hd__inv_2
X_11643_ _18977_/X _11640_/X _21103_/Q _11642_/X vssd1 vssd1 vccd1 vccd1 _21103_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13232__B1 _13148_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18553__S _18908_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20128__RESET_B repeater245/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17150_ _17292_/A vssd1 vssd1 vccd1 vccd1 _17150_/X sky130_fd_sc_hd__buf_1
XPHY_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14362_ _14498_/A _14497_/C _14362_/C _14362_/D vssd1 vssd1 vccd1 vccd1 _14463_/A
+ sky130_fd_sc_hd__or4_4
X_11574_ _21127_/Q _11562_/X _11573_/X _11566_/X vssd1 vssd1 vccd1 vccd1 _21127_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput17 HADDR[24] vssd1 vssd1 vccd1 vccd1 input17/X sky130_fd_sc_hd__buf_1
XPHY_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10597__B2 _20762_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16101_ _16101_/A vssd1 vssd1 vccd1 vccd1 _16101_/X sky130_fd_sc_hd__buf_1
Xinput28 HADDR[5] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__buf_1
XPHY_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10525_ _10827_/A vssd1 vssd1 vccd1 vccd1 _10824_/A sky130_fd_sc_hd__clkbuf_2
Xinput39 HWDATA[10] vssd1 vssd1 vccd1 vccd1 input39/X sky130_fd_sc_hd__buf_2
XPHY_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13313_ _13313_/A vssd1 vssd1 vccd1 vccd1 _13313_/X sky130_fd_sc_hd__buf_2
X_14293_ _20123_/Q vssd1 vssd1 vccd1 vccd1 _14293_/X sky130_fd_sc_hd__buf_1
XFILLER_6_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17081_ _18079_/A vssd1 vssd1 vccd1 vccd1 _17808_/A sky130_fd_sc_hd__buf_4
X_13244_ _20571_/Q _13239_/X _13243_/X _13241_/X vssd1 vssd1 vccd1 vccd1 _20571_/D
+ sky130_fd_sc_hd__a22o_1
X_16032_ _19519_/Q _16028_/X _15774_/X _16029_/X vssd1 vssd1 vccd1 vccd1 _19519_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_109_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10456_ _20677_/Q vssd1 vssd1 vccd1 vccd1 _10456_/Y sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_4_14_0_HCLK_A clkbuf_3_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13175_ _13175_/A vssd1 vssd1 vccd1 vccd1 _16525_/A sky130_fd_sc_hd__buf_1
X_10387_ _10279_/A _10279_/B _10385_/Y _10383_/X vssd1 vssd1 vccd1 vccd1 _21364_/D
+ sky130_fd_sc_hd__a211oi_2
X_12126_ _20384_/Q vssd1 vssd1 vccd1 vccd1 _17975_/A sky130_fd_sc_hd__inv_2
XFILLER_124_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17983_ _20831_/Q _18007_/B vssd1 vssd1 vccd1 vccd1 _17983_/Y sky130_fd_sc_hd__nand2_1
XFILLER_238_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19722_ _20327_/CLK _19722_/D vssd1 vssd1 vccd1 vccd1 _19722_/Q sky130_fd_sc_hd__dfxtp_1
X_12057_ _20371_/Q vssd1 vssd1 vccd1 vccd1 _12057_/Y sky130_fd_sc_hd__inv_2
X_16934_ _19962_/Q _16930_/A _16933_/Y _16930_/Y vssd1 vssd1 vccd1 vccd1 _16935_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_78_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11008_ _15413_/A _11008_/B vssd1 vssd1 vccd1 vccd1 _11909_/B sky130_fd_sc_hd__or2_1
X_19653_ _19821_/CLK _19653_/D vssd1 vssd1 vccd1 vccd1 _19653_/Q sky130_fd_sc_hd__dfxtp_1
X_16865_ _19945_/Q vssd1 vssd1 vccd1 vccd1 _16865_/Y sky130_fd_sc_hd__inv_2
XFILLER_226_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18728__S _18908_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17985__B1 _18339_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18604_ _18845_/A0 _13819_/Y _18896_/S vssd1 vssd1 vccd1 vccd1 _18604_/X sky130_fd_sc_hd__mux2_1
XFILLER_219_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15816_ _15816_/A _16165_/B _16419_/C vssd1 vssd1 vccd1 vccd1 _15824_/A sky130_fd_sc_hd__or3_4
XANTENNA__20969__RESET_B repeater186/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15941__A _16332_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_225_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19584_ _21021_/CLK _19584_/D vssd1 vssd1 vccd1 vccd1 _19584_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16796_ _16794_/Y _16795_/Y _16779_/X vssd1 vssd1 vccd1 vccd1 _16796_/X sky130_fd_sc_hd__o21a_1
XFILLER_225_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18535_ _18848_/A0 _17921_/Y _18666_/S vssd1 vssd1 vccd1 vccd1 _18535_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15747_ _19652_/Q _15743_/X _15730_/X _15745_/X vssd1 vssd1 vccd1 vccd1 _19652_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13471__B1 _13284_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12959_ _20707_/Q _12948_/X _12872_/X _12951_/X vssd1 vssd1 vccd1 vccd1 _20707_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13461__A _13483_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18466_ _17830_/X _10928_/Y _18928_/S vssd1 vssd1 vccd1 vccd1 _18466_/X sky130_fd_sc_hd__mux2_1
XFILLER_179_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15678_ _19684_/Q _15674_/X _15661_/X _15676_/X vssd1 vssd1 vccd1 vccd1 _19684_/D
+ sky130_fd_sc_hd__a22o_1
X_17417_ _19505_/Q vssd1 vssd1 vccd1 vccd1 _17417_/Y sky130_fd_sc_hd__inv_2
X_14629_ _14579_/A _14579_/B _14621_/X _14627_/Y vssd1 vssd1 vccd1 vccd1 _20190_/D
+ sky130_fd_sc_hd__a211oi_2
X_18397_ _18396_/X _10583_/Y _18879_/S vssd1 vssd1 vccd1 vccd1 _18397_/X sky130_fd_sc_hd__mux2_1
XANTENNA__18463__S _18617_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09978__B1 _09685_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20346__CLK _20930_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14971__B1 _14970_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17348_ _17348_/A vssd1 vssd1 vccd1 vccd1 _17348_/X sky130_fd_sc_hd__buf_1
XFILLER_147_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17279_ _21432_/Q _17449_/A vssd1 vssd1 vccd1 vccd1 _17279_/X sky130_fd_sc_hd__and2_1
X_19018_ _16920_/Y _20405_/Q _19019_/S vssd1 vssd1 vccd1 vccd1 _19958_/D sky130_fd_sc_hd__mux2_1
XFILLER_228_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20290_ _20661_/CLK _20290_/D repeater261/X vssd1 vssd1 vccd1 vccd1 _20290_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_228_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11537__B1 _10896_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18217__A1 input70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_8_HCLK_A clkbuf_opt_2_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_119_HCLK clkbuf_opt_3_HCLK/A vssd1 vssd1 vccd1 vccd1 _20980_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_29_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18638__S _18849_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09604_ _14304_/A vssd1 vssd1 vccd1 vccd1 _13048_/A sky130_fd_sc_hd__buf_1
XFILLER_244_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_244_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13462__B1 _13265_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_240_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20292__RESET_B repeater263/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18373__S _18787_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20221__RESET_B repeater202/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20626_ _20626_/CLK _20626_/D repeater193/X vssd1 vssd1 vccd1 vccd1 _20626_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18153__A0 _18152_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10579__B2 _20755_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20557_ _20592_/CLK _20557_/D repeater267/X vssd1 vssd1 vccd1 vccd1 _20557_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12715__A _12715_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10310_ _21357_/Q _20716_/Q _10272_/A _10309_/Y vssd1 vssd1 vccd1 vccd1 _10310_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_4_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14714__B1 _12863_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11290_ _11290_/A _11290_/B _11290_/C _11299_/D vssd1 vssd1 vccd1 vccd1 _16568_/A
+ sky130_fd_sc_hd__nor4_2
XFILLER_165_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20488_ _20937_/CLK _20488_/D repeater277/X vssd1 vssd1 vccd1 vccd1 _20488_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_138_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10241_ _21362_/Q vssd1 vssd1 vccd1 vccd1 _10277_/A sky130_fd_sc_hd__inv_2
XFILLER_133_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17664__C1 _17661_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10172_ _10172_/A vssd1 vssd1 vccd1 vccd1 _10172_/Y sky130_fd_sc_hd__inv_2
XFILLER_160_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21109_ _21417_/CLK _21109_/D repeater234/X vssd1 vssd1 vccd1 vccd1 _21109_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_154_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14980_ _14963_/D _14876_/B _14977_/Y _14975_/X vssd1 vssd1 vccd1 vccd1 _20098_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_120_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13931_ _20660_/Q vssd1 vssd1 vccd1 vccd1 _13931_/Y sky130_fd_sc_hd__inv_2
XFILLER_208_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18548__S _18903_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16650_ _16652_/A _18955_/X vssd1 vssd1 vccd1 vccd1 _19859_/D sky130_fd_sc_hd__and2_1
XFILLER_19_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13862_ _20294_/Q vssd1 vssd1 vccd1 vccd1 _13865_/A sky130_fd_sc_hd__inv_2
XFILLER_234_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15601_ _19723_/Q _15596_/X _15475_/X _15598_/X vssd1 vssd1 vccd1 vccd1 _19723_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_74_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12813_ _12815_/A _13106_/B vssd1 vssd1 vccd1 vccd1 _12814_/S sky130_fd_sc_hd__or2_1
X_16581_ _16689_/B vssd1 vssd1 vccd1 vccd1 _16585_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_16_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13793_ _20604_/Q vssd1 vssd1 vccd1 vccd1 _13793_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13453__B1 _13452_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18320_ _18319_/X _12191_/Y _18909_/S vssd1 vssd1 vccd1 vccd1 _18320_/X sky130_fd_sc_hd__mux2_1
X_15532_ _19757_/Q _15529_/X _15450_/X _15531_/X vssd1 vssd1 vccd1 vccd1 _19757_/D
+ sky130_fd_sc_hd__a22o_1
X_12744_ _12968_/A _16526_/A _20807_/Q _12739_/Y _12743_/X vssd1 vssd1 vccd1 vccd1
+ _12751_/B sky130_fd_sc_hd__a41o_1
XANTENNA__18392__A0 _18391_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18251_ _18250_/X _20585_/Q _18907_/S vssd1 vssd1 vccd1 vccd1 _18251_/X sky130_fd_sc_hd__mux2_1
X_15463_ _19783_/Q _15459_/X _15429_/X _15460_/X vssd1 vssd1 vccd1 vccd1 _19783_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14527__D _17320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13205__B1 _13003_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12675_ _20834_/Q _12672_/X _12673_/X _12674_/X vssd1 vssd1 vccd1 vccd1 _20834_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18283__S _18644_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17202_ _17575_/A vssd1 vssd1 vccd1 vccd1 _18048_/A sky130_fd_sc_hd__buf_2
X_14414_ _21463_/Q vssd1 vssd1 vccd1 vccd1 _14414_/Y sky130_fd_sc_hd__inv_2
XPHY_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11626_ _21105_/Q vssd1 vssd1 vccd1 vccd1 _11632_/A sky130_fd_sc_hd__inv_2
X_18182_ _17810_/Y _21471_/Q _18669_/S vssd1 vssd1 vccd1 vccd1 _18182_/X sky130_fd_sc_hd__mux2_1
XPHY_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15394_ _19814_/Q _15389_/X _15355_/X _15390_/X vssd1 vssd1 vccd1 vccd1 _19814_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17133_ _17133_/A _17133_/B vssd1 vssd1 vccd1 vccd1 _18920_/S sky130_fd_sc_hd__nor2_4
X_14345_ _20221_/Q vssd1 vssd1 vccd1 vccd1 _14460_/D sky130_fd_sc_hd__inv_2
X_11557_ _21132_/Q _11552_/X _10889_/X _11554_/X vssd1 vssd1 vccd1 vccd1 _21132_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10508_ _21278_/Q _10506_/Y _21304_/Q _10507_/Y vssd1 vssd1 vccd1 vccd1 _10508_/X
+ sky130_fd_sc_hd__o22a_1
X_17064_ _17064_/A _17064_/B vssd1 vssd1 vccd1 vccd1 _19880_/D sky130_fd_sc_hd__and2_1
X_14276_ _20124_/Q vssd1 vssd1 vccd1 vccd1 _14276_/Y sky130_fd_sc_hd__inv_2
XANTENNA_output99_A _18076_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11488_ _20872_/Q _11488_/B vssd1 vssd1 vccd1 vccd1 _17140_/B sky130_fd_sc_hd__or2_1
XANTENNA__21168__RESET_B repeater220/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16015_ _19527_/Q _16008_/X _16014_/X _16010_/X vssd1 vssd1 vccd1 vccd1 _19527_/D
+ sky130_fd_sc_hd__a22o_1
X_10439_ _10780_/A _20693_/Q _21291_/Q _17900_/A _10438_/X vssd1 vssd1 vccd1 vccd1
+ _10446_/C sky130_fd_sc_hd__o221a_1
XANTENNA__15936__A _15943_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13227_ _13227_/A vssd1 vssd1 vccd1 vccd1 _13249_/A sky130_fd_sc_hd__buf_1
XANTENNA__18447__A1 _10635_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16458__B1 _16332_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09934__A _20890_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13158_ _13165_/A vssd1 vssd1 vccd1 vccd1 _13158_/X sky130_fd_sc_hd__buf_1
XFILLER_69_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18031__B _18032_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12109_ _12308_/A vssd1 vssd1 vccd1 vccd1 _12109_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__13456__A _13657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17966_ _17925_/X _17966_/B _17966_/C vssd1 vssd1 vccd1 vccd1 _17966_/Y sky130_fd_sc_hd__nand3b_4
X_13089_ _20644_/Q _13086_/X _12863_/X _13087_/X vssd1 vssd1 vccd1 vccd1 _20644_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16917_ _19958_/Q vssd1 vssd1 vccd1 vccd1 _16917_/Y sky130_fd_sc_hd__inv_2
X_19705_ _19828_/CLK _19705_/D vssd1 vssd1 vccd1 vccd1 _19705_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13692__B1 _12857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17897_ _17897_/A _17898_/B vssd1 vssd1 vccd1 vccd1 _17897_/Y sky130_fd_sc_hd__nor2_1
XFILLER_238_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18458__S _18896_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19636_ _20142_/CLK _19636_/D vssd1 vssd1 vccd1 vccd1 _19636_/Q sky130_fd_sc_hd__dfxtp_1
X_16848_ _16848_/A vssd1 vssd1 vccd1 vccd1 _16848_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_38_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_226_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20732__RESET_B repeater257/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19567_ _19812_/CLK _19567_/D vssd1 vssd1 vccd1 vccd1 _19567_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16779_ _16779_/A vssd1 vssd1 vccd1 vccd1 _16779_/X sky130_fd_sc_hd__buf_2
XFILLER_241_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18518_ _18848_/A0 _14133_/Y _18902_/S vssd1 vssd1 vccd1 vccd1 _18518_/X sky130_fd_sc_hd__mux2_1
XFILLER_230_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19498_ _20327_/CLK _19498_/D vssd1 vssd1 vccd1 vccd1 _19498_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18449_ _18845_/A0 _10342_/Y _18884_/S vssd1 vssd1 vccd1 vccd1 _18449_/X sky130_fd_sc_hd__mux2_1
XFILLER_221_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18193__S _18644_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21460_ _21461_/CLK _21460_/D repeater245/X vssd1 vssd1 vccd1 vccd1 _21460_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__14944__B1 _20594_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20411_ _20413_/CLK _20411_/D repeater185/X vssd1 vssd1 vccd1 vccd1 _20411_/Q sky130_fd_sc_hd__dfrtp_1
X_21391_ _21401_/CLK _21391_/D repeater241/X vssd1 vssd1 vccd1 vccd1 _21391_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18921__S _18926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20342_ _20949_/CLK _20342_/D repeater269/X vssd1 vssd1 vccd1 vccd1 _20342_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_190_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20273_ _20293_/CLK _20273_/D repeater263/X vssd1 vssd1 vccd1 vccd1 _20273_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__19986__RESET_B repeater185/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19915__RESET_B repeater225/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_144_HCLK_A clkbuf_4_3_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15121__B1 _15097_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17949__B1 _18521_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18368__S _18617_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13435__B1 _13313_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10790_ _10790_/A vssd1 vssd1 vccd1 vccd1 _10790_/Y sky130_fd_sc_hd__inv_2
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12460_ _12423_/A _12423_/B _12453_/X _12458_/Y vssd1 vssd1 vccd1 vccd1 _20934_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_130_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11411_ _11411_/A _11776_/B _11786_/C vssd1 vssd1 vccd1 vccd1 _11412_/D sky130_fd_sc_hd__or3_2
X_12391_ _12453_/A vssd1 vssd1 vccd1 vccd1 _12445_/A sky130_fd_sc_hd__clkbuf_2
X_20609_ _20657_/CLK _20609_/D repeater198/X vssd1 vssd1 vccd1 vccd1 _20609_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__18831__S _18927_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11342_ _11342_/A vssd1 vssd1 vccd1 vccd1 _11412_/C sky130_fd_sc_hd__inv_2
X_14130_ _20558_/Q vssd1 vssd1 vccd1 vccd1 _14130_/Y sky130_fd_sc_hd__inv_2
XFILLER_192_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__21261__RESET_B repeater233/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11273_ _20910_/Q _20909_/Q _20912_/Q _20911_/Q vssd1 vssd1 vccd1 vccd1 _12505_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_106_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14061_ _20267_/Q vssd1 vssd1 vccd1 vccd1 _14078_/A sky130_fd_sc_hd__inv_2
XFILLER_152_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13012_ _13012_/A vssd1 vssd1 vccd1 vccd1 _13012_/X sky130_fd_sc_hd__buf_1
XANTENNA_input50_A HWDATA[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10224_ _10224_/A vssd1 vssd1 vccd1 vccd1 _10227_/A sky130_fd_sc_hd__inv_2
XFILLER_79_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17820_ _17820_/A vssd1 vssd1 vccd1 vccd1 _17951_/A sky130_fd_sc_hd__clkbuf_2
X_10155_ _10155_/A _10155_/B vssd1 vssd1 vccd1 vccd1 _10187_/A sky130_fd_sc_hd__or2_1
XFILLER_0_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17751_ _19781_/Q vssd1 vssd1 vccd1 vccd1 _17751_/Y sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_66_HCLK_A clkbuf_4_11_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14963_ _14963_/A _14963_/B _14963_/C _14963_/D vssd1 vssd1 vccd1 vccd1 _14965_/C
+ sky130_fd_sc_hd__or4_4
X_10086_ _20804_/Q vssd1 vssd1 vccd1 vccd1 _10086_/Y sky130_fd_sc_hd__inv_2
XFILLER_47_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output137_A _20043_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16702_ _16720_/A vssd1 vssd1 vccd1 vccd1 _16709_/A sky130_fd_sc_hd__buf_1
XFILLER_208_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17404__A2 _17324_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13914_ _13914_/A _13914_/B _13914_/C _13914_/D vssd1 vssd1 vccd1 vccd1 _13962_/A
+ sky130_fd_sc_hd__and4_1
X_17682_ _19604_/Q _17829_/B vssd1 vssd1 vccd1 vccd1 _17682_/X sky130_fd_sc_hd__and2_1
X_14894_ _14894_/A _14894_/B _14892_/X _14893_/X vssd1 vssd1 vccd1 vccd1 _14901_/B
+ sky130_fd_sc_hd__or4bb_1
XFILLER_90_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19421_ _19828_/CLK _19421_/D vssd1 vssd1 vccd1 vccd1 _19421_/Q sky130_fd_sc_hd__dfxtp_1
X_16633_ _21074_/Q vssd1 vssd1 vccd1 vccd1 _16633_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13845_ _20315_/Q vssd1 vssd1 vccd1 vccd1 _13891_/A sky130_fd_sc_hd__inv_2
XFILLER_223_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20143__RESET_B repeater249/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11524__A _17290_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19352_ _20137_/CLK _19352_/D vssd1 vssd1 vccd1 vccd1 _19352_/Q sky130_fd_sc_hd__dfxtp_1
X_16564_ _16564_/A _16564_/B vssd1 vssd1 vccd1 vccd1 _16564_/X sky130_fd_sc_hd__or2_1
X_13776_ _20204_/Q vssd1 vssd1 vccd1 vccd1 _14593_/A sky130_fd_sc_hd__inv_2
XFILLER_200_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10988_ _21018_/Q vssd1 vssd1 vccd1 vccd1 _10988_/X sky130_fd_sc_hd__buf_1
XFILLER_204_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18303_ _17079_/Y _15255_/Y _18908_/S vssd1 vssd1 vccd1 vccd1 _18303_/X sky130_fd_sc_hd__mux2_1
XFILLER_203_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15515_ _19762_/Q _15507_/X _15514_/X _15509_/X vssd1 vssd1 vccd1 vccd1 _19762_/D
+ sky130_fd_sc_hd__a22o_1
X_12727_ _13329_/A vssd1 vssd1 vccd1 vccd1 _13108_/B sky130_fd_sc_hd__buf_4
X_19283_ _19765_/Q _19757_/Q _19749_/Q _19741_/Q _19285_/S0 _21017_/Q vssd1 vssd1
+ vccd1 vccd1 _19283_/X sky130_fd_sc_hd__mux4_1
X_16495_ _21095_/Q vssd1 vssd1 vccd1 vccd1 _16495_/Y sky130_fd_sc_hd__inv_2
XFILLER_204_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18234_ _20858_/Q input7/X _18236_/S vssd1 vssd1 vccd1 vccd1 _18234_/X sky130_fd_sc_hd__mux2_1
X_15446_ _19790_/Q _15441_/X _15431_/X _15442_/X vssd1 vssd1 vccd1 vccd1 _19790_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12658_ input59/X vssd1 vssd1 vccd1 vccd1 _12658_/X sky130_fd_sc_hd__clkbuf_4
XPHY_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__21349__RESET_B repeater210/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19407__CLK _19813_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18165_ _18164_/X _14101_/Y _18904_/S vssd1 vssd1 vccd1 vccd1 _18165_/X sky130_fd_sc_hd__mux2_1
X_11609_ _21260_/Q _11596_/A _21113_/Q _11605_/X vssd1 vssd1 vccd1 vccd1 _21113_/D
+ sky130_fd_sc_hd__a22o_1
X_15377_ _15377_/A vssd1 vssd1 vccd1 vccd1 _15657_/A sky130_fd_sc_hd__clkbuf_2
X_12589_ _12601_/A vssd1 vssd1 vccd1 vccd1 _12589_/X sky130_fd_sc_hd__buf_1
XANTENNA__18741__S _18875_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17116_ _19317_/Q vssd1 vssd1 vccd1 vccd1 _17116_/Y sky130_fd_sc_hd__inv_2
X_14328_ _14328_/A vssd1 vssd1 vccd1 vccd1 _14378_/A sky130_fd_sc_hd__buf_1
XFILLER_172_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_opt_1_HCLK clkbuf_opt_1_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_opt_1_HCLK/X
+ sky130_fd_sc_hd__clkbuf_16
X_18096_ _18630_/X _17219_/X _18653_/X _18064_/X _18095_/X vssd1 vssd1 vccd1 vccd1
+ _18097_/C sky130_fd_sc_hd__o221a_1
XFILLER_144_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14154__A1 _20540_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17047_ _11457_/A _19287_/Q _11459_/A vssd1 vssd1 vccd1 vccd1 _17048_/B sky130_fd_sc_hd__o21a_1
XFILLER_132_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14259_ _14267_/A vssd1 vssd1 vccd1 vccd1 _14268_/A sky130_fd_sc_hd__inv_2
XANTENNA__19093__A1 _21085_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18998_ _17006_/Y _20425_/Q _19026_/S vssd1 vssd1 vccd1 vccd1 _19978_/D sky130_fd_sc_hd__mux2_1
Xrepeater201 repeater205/X vssd1 vssd1 vccd1 vccd1 repeater201/X sky130_fd_sc_hd__buf_4
XANTENNA__20913__RESET_B repeater218/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater212 repeater215/X vssd1 vssd1 vccd1 vccd1 repeater212/X sky130_fd_sc_hd__buf_8
Xrepeater223 repeater224/X vssd1 vssd1 vccd1 vccd1 repeater223/X sky130_fd_sc_hd__buf_6
XFILLER_112_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18188__S _18617_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13665__B1 _13545_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17949_ _18532_/X _17947_/X _18521_/X _17948_/X vssd1 vssd1 vccd1 vccd1 _17957_/A
+ sky130_fd_sc_hd__o22ai_2
Xrepeater234 repeater236/X vssd1 vssd1 vccd1 vccd1 repeater234/X sky130_fd_sc_hd__buf_8
Xrepeater245 repeater246/X vssd1 vssd1 vccd1 vccd1 repeater245/X sky130_fd_sc_hd__buf_8
XFILLER_94_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater256 repeater257/X vssd1 vssd1 vccd1 vccd1 repeater256/X sky130_fd_sc_hd__buf_8
XFILLER_238_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20960_ _20981_/CLK _20960_/D repeater186/X vssd1 vssd1 vccd1 vccd1 _20960_/Q sky130_fd_sc_hd__dfrtp_1
Xrepeater267 repeater268/X vssd1 vssd1 vccd1 vccd1 repeater267/X sky130_fd_sc_hd__buf_8
Xrepeater278 repeater279/X vssd1 vssd1 vccd1 vccd1 repeater278/X sky130_fd_sc_hd__buf_6
XANTENNA__15832__C _15832_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19619_ _21453_/CLK _19619_/D vssd1 vssd1 vccd1 vccd1 _19619_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17800__C1 _17799_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20891_ _21449_/CLK _20891_/D repeater248/X vssd1 vssd1 vccd1 vccd1 _20891_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_3709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21443_ _21444_/CLK _21443_/D repeater246/X vssd1 vssd1 vccd1 vccd1 _21443_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_21_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12265__A _20499_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18651__S _18886_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21019__RESET_B repeater238/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21374_ _21374_/CLK _21374_/D repeater257/X vssd1 vssd1 vccd1 vccd1 _21374_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_119_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20325_ _20326_/CLK _20325_/D repeater250/X vssd1 vssd1 vccd1 vccd1 _20325_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_123_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15342__B1 _14264_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20256_ _20256_/CLK _20256_/D repeater217/X vssd1 vssd1 vccd1 vccd1 _20256_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_1_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20187_ _20623_/CLK _20187_/D repeater194/X vssd1 vssd1 vccd1 vccd1 _20187_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__10513__A _20691_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09998_ _17036_/A vssd1 vssd1 vccd1 vccd1 _09998_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13656__B1 _13454_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11960_ _21001_/Q _21000_/Q vssd1 vssd1 vccd1 vccd1 _13185_/B sky130_fd_sc_hd__nand2_1
XFILLER_57_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10911_ _20702_/Q vssd1 vssd1 vccd1 vccd1 _12750_/A sky130_fd_sc_hd__inv_2
XFILLER_233_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18826__S _18927_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11891_ _21022_/Q _11883_/X _11877_/A _11890_/X vssd1 vssd1 vccd1 vccd1 _21022_/D
+ sky130_fd_sc_hd__a31o_1
X_13630_ _20380_/Q _13625_/X _13489_/X _13626_/X vssd1 vssd1 vccd1 vccd1 _20380_/D
+ sky130_fd_sc_hd__a22o_1
X_10842_ _10842_/A _20033_/Q vssd1 vssd1 vccd1 vccd1 _14307_/C sky130_fd_sc_hd__nor2_1
XFILLER_44_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18898__A1 _14566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13561_ _13567_/A vssd1 vssd1 vccd1 vccd1 _13561_/X sky130_fd_sc_hd__buf_1
X_10773_ _10773_/A _10773_/B vssd1 vssd1 vccd1 vccd1 _10804_/A sky130_fd_sc_hd__or2_1
XFILLER_201_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15300_ _15302_/A vssd1 vssd1 vccd1 vccd1 _15305_/A sky130_fd_sc_hd__inv_2
XFILLER_197_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12512_ _12512_/A vssd1 vssd1 vccd1 vccd1 _12512_/Y sky130_fd_sc_hd__inv_2
XFILLER_201_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16280_ _19397_/Q _16276_/X _16277_/X _16279_/X vssd1 vssd1 vccd1 vccd1 _19397_/D
+ sky130_fd_sc_hd__a22o_1
X_13492_ _13514_/A vssd1 vssd1 vccd1 vccd1 _13492_/X sky130_fd_sc_hd__buf_1
XFILLER_13_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21442__RESET_B repeater245/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15231_ _20477_/Q _15070_/A _20465_/Q _15059_/A _15230_/X vssd1 vssd1 vccd1 vccd1
+ _15232_/D sky130_fd_sc_hd__o221a_1
XFILLER_60_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12443_ _12443_/A vssd1 vssd1 vccd1 vccd1 _12443_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18561__S _18897_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15581__B1 _15550_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15162_ _15185_/A vssd1 vssd1 vccd1 vccd1 _15193_/A sky130_fd_sc_hd__inv_2
XFILLER_138_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12374_ _20961_/Q _12376_/B _12373_/X _12315_/B vssd1 vssd1 vccd1 vccd1 _20961_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_126_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14113_ _20554_/Q vssd1 vssd1 vccd1 vccd1 _18031_/A sky130_fd_sc_hd__inv_2
X_11325_ _19844_/Q vssd1 vssd1 vccd1 vccd1 _11371_/A sky130_fd_sc_hd__inv_2
XANTENNA__15333__B1 _13557_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14390__A _20031_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19970_ _20422_/CLK _19970_/D repeater184/X vssd1 vssd1 vccd1 vccd1 _19970_/Q sky130_fd_sc_hd__dfrtp_1
X_15093_ _15093_/A vssd1 vssd1 vccd1 vccd1 _15093_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_5_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20557__CLK _20592_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11256_ _19908_/Q vssd1 vssd1 vccd1 vccd1 _16689_/A sky130_fd_sc_hd__buf_1
XANTENNA__19075__A1 _20900_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18921_ _17132_/Y _17131_/Y _18926_/S vssd1 vssd1 vccd1 vccd1 _18921_/X sky130_fd_sc_hd__mux2_1
XFILLER_69_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14044_ _20284_/Q vssd1 vssd1 vccd1 vccd1 _14094_/A sky130_fd_sc_hd__inv_2
XANTENNA__19170__S1 _20122_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold9_A hold9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10207_ _10207_/A _10207_/B vssd1 vssd1 vccd1 vccd1 _10207_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_repeater202_A repeater203/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18852_ _18851_/X _15154_/Y _18906_/S vssd1 vssd1 vccd1 vccd1 _18852_/X sky130_fd_sc_hd__mux2_1
X_11187_ _11187_/A vssd1 vssd1 vccd1 vccd1 _17133_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_122_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17803_ _18378_/X _17856_/A _18141_/X _17480_/X vssd1 vssd1 vccd1 vccd1 _17803_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_94_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10138_ _10185_/A vssd1 vssd1 vccd1 vccd1 _10260_/B sky130_fd_sc_hd__inv_2
XFILLER_227_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18783_ _17079_/Y _15243_/Y _18908_/S vssd1 vssd1 vccd1 vccd1 _18783_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15995_ _19537_/Q _15993_/X _15944_/X _15994_/X vssd1 vssd1 vccd1 vccd1 _19537_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13647__B1 _13506_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20324__RESET_B repeater250/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17734_ _18694_/X _17839_/A _18697_/X _17869_/A _17733_/X vssd1 vssd1 vccd1 vccd1
+ _17734_/X sky130_fd_sc_hd__o221a_2
X_14946_ _20580_/Q _14962_/A _14945_/Y _20107_/Q vssd1 vssd1 vccd1 vccd1 _14946_/X
+ sky130_fd_sc_hd__o22a_1
X_10069_ _21399_/Q vssd1 vssd1 vccd1 vccd1 _10160_/A sky130_fd_sc_hd__inv_2
XFILLER_48_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17665_ _17548_/X _17646_/X _17560_/X _17655_/X _17664_/X vssd1 vssd1 vccd1 vccd1
+ _17665_/Y sky130_fd_sc_hd__o221ai_4
XANTENNA__12870__A1 _20744_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14877_ _14963_/C _14977_/A vssd1 vssd1 vccd1 vccd1 _14878_/B sky130_fd_sc_hd__or2_1
XFILLER_223_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18736__S _18926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16616_ _16616_/A _16616_/B vssd1 vssd1 vccd1 vccd1 _16616_/Y sky130_fd_sc_hd__nor2_1
X_19404_ _21011_/CLK _19404_/D vssd1 vssd1 vccd1 vccd1 _19404_/Q sky130_fd_sc_hd__dfxtp_1
X_13828_ _20607_/Q _14574_/A _20624_/Q _14590_/A vssd1 vssd1 vccd1 vccd1 _13828_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_211_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17596_ _19523_/Q vssd1 vssd1 vccd1 vccd1 _17596_/Y sky130_fd_sc_hd__inv_2
X_16547_ _21149_/Q vssd1 vssd1 vccd1 vccd1 _16547_/Y sky130_fd_sc_hd__inv_2
X_19335_ _20172_/CLK _19335_/D vssd1 vssd1 vccd1 vccd1 _19335_/Q sky130_fd_sc_hd__dfxtp_1
X_13759_ _18081_/A _20205_/Q _20606_/Q _14573_/A vssd1 vssd1 vccd1 vccd1 _13759_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17010__B1 _16984_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19266_ _19262_/X _19263_/X _19264_/X _19265_/X _21005_/Q _21006_/Q vssd1 vssd1 vccd1
+ vccd1 _19266_/X sky130_fd_sc_hd__mux4_2
XANTENNA__09659__A _12863_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16478_ _19292_/Q _16473_/X _16295_/X _16474_/X vssd1 vssd1 vccd1 vccd1 _19292_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__21183__RESET_B repeater216/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18217_ _21040_/Q input70/X _18242_/S vssd1 vssd1 vccd1 vccd1 _18217_/X sky130_fd_sc_hd__mux2_1
X_15429_ _15429_/A vssd1 vssd1 vccd1 vccd1 _15429_/X sky130_fd_sc_hd__clkbuf_2
X_19197_ _17757_/Y _17758_/Y _17759_/Y _17760_/Y _20130_/Q _20131_/Q vssd1 vssd1 vccd1
+ vccd1 _19197_/X sky130_fd_sc_hd__mux4_1
XANTENNA__18471__S _18680_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18148_ _18003_/Y _20656_/Q _18903_/S vssd1 vssd1 vccd1 vccd1 _18148_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18079_ _18079_/A vssd1 vssd1 vccd1 vccd1 _18083_/B sky130_fd_sc_hd__buf_2
XANTENNA__12813__A _12815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20110_ _21433_/CLK _20110_/D repeater234/X vssd1 vssd1 vccd1 vccd1 _20110_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_236_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09921_ _21437_/Q _21438_/Q _09924_/S vssd1 vssd1 vccd1 vccd1 _21438_/D sky130_fd_sc_hd__mux2_1
XANTENNA__19066__A1 _21127_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21090_ _21424_/CLK _21090_/D repeater230/X vssd1 vssd1 vccd1 vccd1 _21090_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_131_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20041_ _20042_/CLK _20041_/D repeater219/X vssd1 vssd1 vccd1 vccd1 _20041_/Q sky130_fd_sc_hd__dfstp_1
X_09852_ _09864_/A vssd1 vssd1 vccd1 vccd1 _09852_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09783_ _09783_/A vssd1 vssd1 vccd1 vccd1 _16619_/B sky130_fd_sc_hd__buf_1
XANTENNA__13638__B1 _13426_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18577__A0 _18848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_215_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20943_ _20943_/CLK _20943_/D repeater275/X vssd1 vssd1 vccd1 vccd1 _20943_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_215_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18646__S _18875_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11164__A _16616_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18329__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20874_ _21459_/CLK _20874_/D repeater244/X vssd1 vssd1 vccd1 vccd1 _20874_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_54_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18381__S _18908_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21426_ _21429_/CLK _21426_/D repeater229/X vssd1 vssd1 vccd1 vccd1 _21426_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_136_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19930__RESET_B repeater251/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21357_ _21357_/CLK _21357_/D repeater199/X vssd1 vssd1 vccd1 vccd1 _21357_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_162_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11110_ _11105_/B _11109_/Y _11051_/X _11101_/X _11053_/A vssd1 vssd1 vccd1 vccd1
+ _11111_/A sky130_fd_sc_hd__o32a_1
XFILLER_146_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20308_ _20316_/CLK _20308_/D repeater196/X vssd1 vssd1 vccd1 vccd1 _20308_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__20835__RESET_B repeater257/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12090_ _20380_/Q vssd1 vssd1 vccd1 vccd1 _12090_/Y sky130_fd_sc_hd__inv_2
X_21288_ _21306_/CLK _21288_/D repeater207/X vssd1 vssd1 vccd1 vccd1 _21288_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_146_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11041_ _19977_/Q _19976_/Q _11041_/C _16989_/B vssd1 vssd1 vccd1 vccd1 _17004_/A
+ sky130_fd_sc_hd__or4_4
X_20239_ _21481_/CLK _20239_/D repeater206/X vssd1 vssd1 vccd1 vccd1 _20239_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__19152__S1 _21017_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14800_ _14800_/A _14800_/B vssd1 vssd1 vccd1 vccd1 _14800_/Y sky130_fd_sc_hd__nand2_1
XFILLER_18_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15780_ _15787_/A vssd1 vssd1 vccd1 vccd1 _15789_/A sky130_fd_sc_hd__inv_2
XANTENNA__18568__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12992_ _20695_/Q _12983_/X _12991_/X _12987_/X vssd1 vssd1 vccd1 vccd1 _20695_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input13_A HADDR[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14731_ _14732_/A vssd1 vssd1 vccd1 vccd1 _14731_/X sky130_fd_sc_hd__buf_1
X_11943_ _11943_/A vssd1 vssd1 vccd1 vccd1 _11943_/X sky130_fd_sc_hd__buf_1
XANTENNA__18556__S _18928_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17450_ _20776_/Q vssd1 vssd1 vccd1 vccd1 _17450_/Y sky130_fd_sc_hd__inv_2
XFILLER_189_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14662_ _20129_/Q _16482_/A vssd1 vssd1 vccd1 vccd1 _14663_/B sky130_fd_sc_hd__or2_1
XFILLER_33_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11874_ _21022_/Q vssd1 vssd1 vccd1 vccd1 _11874_/Y sky130_fd_sc_hd__inv_2
XFILLER_233_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16401_ _19336_/Q _16399_/X _16335_/X _16400_/X vssd1 vssd1 vccd1 vccd1 _19336_/D
+ sky130_fd_sc_hd__a22o_1
X_13613_ _13625_/A vssd1 vssd1 vccd1 vccd1 _13613_/X sky130_fd_sc_hd__buf_1
X_17381_ _17390_/A vssd1 vssd1 vccd1 vccd1 _17381_/X sky130_fd_sc_hd__buf_1
X_10825_ _10825_/A vssd1 vssd1 vccd1 vccd1 _10825_/Y sky130_fd_sc_hd__inv_2
X_14593_ _14593_/A _14593_/B vssd1 vssd1 vccd1 vccd1 _14602_/A sky130_fd_sc_hd__or2_1
XANTENNA__12604__B2 _12601_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19120_ _19125_/S _14275_/Y _19126_/S vssd1 vssd1 vccd1 vccd1 _19120_/X sky130_fd_sc_hd__mux2_2
X_16332_ _16332_/A vssd1 vssd1 vccd1 vccd1 _16332_/X sky130_fd_sc_hd__clkbuf_2
X_13544_ _20427_/Q _13537_/X _13543_/X _13541_/X vssd1 vssd1 vccd1 vccd1 _20427_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_185_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10756_ _10756_/A _10756_/B vssd1 vssd1 vccd1 vccd1 _10836_/A sky130_fd_sc_hd__or2_1
XFILLER_187_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19051_ _16780_/X _20818_/Q _19058_/S vssd1 vssd1 vccd1 vccd1 _19925_/D sky130_fd_sc_hd__mux2_1
XFILLER_13_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16263_ _16269_/A vssd1 vssd1 vccd1 vccd1 _16270_/A sky130_fd_sc_hd__inv_2
XANTENNA__18291__S _18787_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13475_ input52/X vssd1 vssd1 vccd1 vccd1 _13475_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_repeater152_A _18902_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10687_ _10687_/A vssd1 vssd1 vccd1 vccd1 _10687_/Y sky130_fd_sc_hd__inv_2
XFILLER_185_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18002_ _18033_/A vssd1 vssd1 vccd1 vccd1 _18006_/B sky130_fd_sc_hd__buf_2
X_15214_ _15214_/A vssd1 vssd1 vccd1 vccd1 _15214_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_185_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12426_ _12426_/A _12455_/A vssd1 vssd1 vccd1 vccd1 _12427_/B sky130_fd_sc_hd__or2_1
X_16194_ _16405_/A _16419_/B _16194_/C vssd1 vssd1 vccd1 vccd1 _16206_/A sky130_fd_sc_hd__or3_4
X_15145_ _20436_/Q vssd1 vssd1 vccd1 vccd1 _15145_/Y sky130_fd_sc_hd__inv_2
X_12357_ _12105_/X _12323_/B _12350_/X _12355_/Y vssd1 vssd1 vccd1 vccd1 _20970_/D
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__17846__A2 _17214_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output81_A _17874_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11308_ _11544_/A vssd1 vssd1 vccd1 vccd1 _11312_/A sky130_fd_sc_hd__inv_2
XFILLER_153_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15076_ _15076_/A _15076_/B vssd1 vssd1 vccd1 vccd1 _15184_/A sky130_fd_sc_hd__or2_1
X_19953_ _21234_/CLK _19953_/D repeater188/X vssd1 vssd1 vccd1 vccd1 _19953_/Q sky130_fd_sc_hd__dfrtp_1
X_12288_ _12432_/A _20523_/Q _20936_/Q _12284_/Y _12287_/X vssd1 vssd1 vccd1 vccd1
+ _12301_/B sky130_fd_sc_hd__o221a_1
Xclkbuf_leaf_10_HCLK clkbuf_opt_2_HCLK/X vssd1 vssd1 vccd1 vccd1 _20432_/CLK sky130_fd_sc_hd__clkbuf_16
X_18904_ _18903_/X _14070_/A _18904_/S vssd1 vssd1 vccd1 vccd1 _18904_/X sky130_fd_sc_hd__mux2_1
XANTENNA__19143__S1 _21017_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14027_ _20296_/Q _14026_/Y _14013_/B _13965_/X vssd1 vssd1 vccd1 vccd1 _20296_/D
+ sky130_fd_sc_hd__o211a_1
X_11239_ _11241_/A _11251_/A vssd1 vssd1 vccd1 vccd1 _11239_/X sky130_fd_sc_hd__or2_1
X_19884_ _21338_/CLK _19884_/D repeater221/X vssd1 vssd1 vccd1 vccd1 _19884_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_68_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18835_ _17281_/X _17284_/Y _18835_/S vssd1 vssd1 vccd1 vccd1 _18835_/X sky130_fd_sc_hd__mux2_1
XFILLER_121_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15978_ _15978_/A vssd1 vssd1 vccd1 vccd1 _15978_/X sky130_fd_sc_hd__buf_1
XFILLER_36_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18766_ _18765_/X _19236_/X _18930_/S vssd1 vssd1 vccd1 vccd1 _18766_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_152_HCLK clkbuf_opt_1_HCLK/X vssd1 vssd1 vccd1 vccd1 _20890_/CLK sky130_fd_sc_hd__clkbuf_16
X_17717_ _16519_/Y _17378_/A _17716_/Y _17390_/X vssd1 vssd1 vccd1 vccd1 _17717_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_64_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14929_ _20582_/Q vssd1 vssd1 vccd1 vccd1 _14929_/Y sky130_fd_sc_hd__inv_2
XFILLER_82_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18466__S _18928_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18697_ _18696_/X _14923_/Y _18907_/S vssd1 vssd1 vccd1 vccd1 _18697_/X sky130_fd_sc_hd__mux2_1
X_17648_ _20898_/Q vssd1 vssd1 vccd1 vccd1 _17648_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__21364__RESET_B repeater254/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17579_ _18756_/X _17472_/A _18755_/X _17474_/A vssd1 vssd1 vccd1 vccd1 _17579_/X
+ sky130_fd_sc_hd__o22a_2
X_19318_ _19961_/CLK _19318_/D vssd1 vssd1 vccd1 vccd1 _19318_/Q sky130_fd_sc_hd__dfxtp_1
X_20590_ _20590_/CLK _20590_/D repeater259/X vssd1 vssd1 vccd1 vccd1 _20590_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_188_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19249_ _17358_/Y _17359_/Y _17360_/Y _17361_/Y _20130_/Q _20131_/Q vssd1 vssd1 vccd1
+ vccd1 _19249_/X sky130_fd_sc_hd__mux4_1
XANTENNA__13384__D_N _20872_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21211_ _21401_/CLK _21211_/D repeater241/X vssd1 vssd1 vccd1 vccd1 _21211_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__20872__CLK _21452_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21142_ _21191_/CLK _21142_/D repeater192/X vssd1 vssd1 vccd1 vccd1 _21142_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_160_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19134__S1 _21017_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09904_ _09904_/A vssd1 vssd1 vccd1 vccd1 _17021_/A sky130_fd_sc_hd__inv_2
X_21073_ _21424_/CLK _21073_/D repeater230/X vssd1 vssd1 vccd1 vccd1 _21073_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_101_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20024_ _21424_/CLK input72/X repeater229/X vssd1 vssd1 vccd1 vccd1 _20024_/Q sky130_fd_sc_hd__dfrtp_1
X_09835_ _15879_/A vssd1 vssd1 vccd1 vccd1 _09835_/X sky130_fd_sc_hd__buf_1
XANTENNA_input5_A HADDR[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09766_ _11055_/A _20150_/Q _21230_/Q _09765_/Y vssd1 vssd1 vccd1 vccd1 _09766_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_73_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12834__A1 _20762_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_227_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18376__S _18748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09697_ _15523_/A vssd1 vssd1 vccd1 vccd1 _10898_/A sky130_fd_sc_hd__buf_1
XPHY_4026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20926_ _20929_/CLK _20926_/D repeater266/X vssd1 vssd1 vccd1 vccd1 _20926_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_215_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20857_ _20857_/CLK _20857_/D repeater243/X vssd1 vssd1 vccd1 vccd1 _20857_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__21034__RESET_B repeater242/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10610_ _20748_/Q vssd1 vssd1 vccd1 vccd1 _10610_/Y sky130_fd_sc_hd__inv_2
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18722__A0 _18848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11590_ _11590_/A _11590_/B vssd1 vssd1 vccd1 vccd1 _11591_/B sky130_fd_sc_hd__nand2_1
XPHY_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20788_ _21390_/CLK _20788_/D repeater240/X vssd1 vssd1 vccd1 vccd1 _20788_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10541_ _21317_/Q vssd1 vssd1 vccd1 vccd1 _10705_/A sky130_fd_sc_hd__inv_2
XPHY_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19000__S _19019_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13260_ _13254_/X _20562_/Q _13260_/S vssd1 vssd1 vccd1 vccd1 _20562_/D sky130_fd_sc_hd__mux2_1
XFILLER_210_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10472_ _20687_/Q vssd1 vssd1 vccd1 vccd1 _10472_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_33_HCLK clkbuf_opt_4_HCLK/A vssd1 vssd1 vccd1 vccd1 _21001_/CLK sky130_fd_sc_hd__clkbuf_16
X_12211_ _20935_/Q vssd1 vssd1 vccd1 vccd1 _12424_/A sky130_fd_sc_hd__inv_2
XANTENNA__13549__A _13566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21409_ _21433_/CLK _21409_/D repeater233/X vssd1 vssd1 vccd1 vccd1 _21409_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_170_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13191_ _13225_/A vssd1 vssd1 vccd1 vccd1 _13215_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_191_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12770__B1 _12670_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12142_ _20959_/Q _12140_/Y _20979_/Q _18077_/A vssd1 vssd1 vccd1 vccd1 _12142_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_190_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16950_ _16958_/C vssd1 vssd1 vccd1 vccd1 _16950_/Y sky130_fd_sc_hd__inv_2
X_12073_ _20951_/Q vssd1 vssd1 vccd1 vccd1 _12073_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_151_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10128__A2 _10126_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11024_ _20808_/Q vssd1 vssd1 vccd1 vccd1 _11024_/Y sky130_fd_sc_hd__inv_2
X_15901_ _19582_/Q _15896_/X _15795_/X _15897_/X vssd1 vssd1 vccd1 vccd1 _19582_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_103_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16881_ _20809_/Q vssd1 vssd1 vccd1 vccd1 _16984_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13284__A input54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18620_ _18845_/A0 _10461_/Y _18896_/S vssd1 vssd1 vccd1 vccd1 _18620_/X sky130_fd_sc_hd__mux2_1
X_15832_ _15832_/A _15832_/B _15832_/C vssd1 vssd1 vccd1 vccd1 _16194_/C sky130_fd_sc_hd__or3_4
XFILLER_206_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15763_ _19644_/Q _15757_/X _15762_/X _15760_/X vssd1 vssd1 vccd1 vccd1 _19644_/D
+ sky130_fd_sc_hd__a22o_1
X_18551_ _18550_/X _10085_/Y _18885_/S vssd1 vssd1 vccd1 vccd1 _18551_/X sky130_fd_sc_hd__mux2_1
XANTENNA__18286__S _18891_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12975_ _12891_/X _20700_/Q _12975_/S vssd1 vssd1 vccd1 vccd1 _20700_/D sky130_fd_sc_hd__mux2_1
XFILLER_245_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14714_ _20154_/Q _14711_/X _12863_/A _14712_/X vssd1 vssd1 vccd1 vccd1 _20154_/D
+ sky130_fd_sc_hd__a22o_1
X_17502_ _17348_/X _17501_/Y _21022_/Q vssd1 vssd1 vccd1 vccd1 _17502_/X sky130_fd_sc_hd__o21a_1
X_11926_ _11926_/A _11926_/B _11926_/C _11926_/D vssd1 vssd1 vccd1 vccd1 _11926_/X
+ sky130_fd_sc_hd__or4_4
X_18482_ _18481_/X _13948_/Y _18903_/S vssd1 vssd1 vccd1 vccd1 _18482_/X sky130_fd_sc_hd__mux2_1
XFILLER_73_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15694_ _15785_/A vssd1 vssd1 vccd1 vccd1 _15694_/X sky130_fd_sc_hd__clkbuf_2
XPHY_4560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17433_ _19609_/Q vssd1 vssd1 vccd1 vccd1 _17433_/Y sky130_fd_sc_hd__inv_2
XPHY_4582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14645_ _14645_/A vssd1 vssd1 vccd1 vccd1 _14645_/Y sky130_fd_sc_hd__inv_2
XPHY_4593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11857_ _11851_/B _11856_/Y _11803_/X _11852_/X _11806_/A vssd1 vssd1 vccd1 vccd1
+ _11858_/A sky130_fd_sc_hd__o32a_1
XFILLER_60_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10808_ _21296_/Q _10807_/Y _10798_/X _10773_/B vssd1 vssd1 vccd1 vccd1 _21296_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_32_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17364_ _19456_/Q vssd1 vssd1 vccd1 vccd1 _17364_/Y sky130_fd_sc_hd__inv_2
XPHY_3892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14576_ _14576_/A _14633_/A vssd1 vssd1 vccd1 vccd1 _14577_/B sky130_fd_sc_hd__or2_2
X_11788_ _21042_/Q _11787_/X _19113_/X vssd1 vssd1 vccd1 vccd1 _21042_/D sky130_fd_sc_hd__mux2_1
XFILLER_220_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18713__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19103_ _16667_/X _21075_/Q _19870_/D vssd1 vssd1 vccd1 vccd1 _19103_/X sky130_fd_sc_hd__mux2_1
X_16315_ _19381_/Q _16312_/X _16231_/X _16314_/X vssd1 vssd1 vccd1 vccd1 _19381_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_119_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13527_ _13527_/A vssd1 vssd1 vccd1 vccd1 _13530_/A sky130_fd_sc_hd__buf_1
X_17295_ _17390_/A vssd1 vssd1 vccd1 vccd1 _17295_/X sky130_fd_sc_hd__buf_1
X_10739_ _19927_/Q _19926_/Q _16777_/A vssd1 vssd1 vccd1 vccd1 _16786_/A sky130_fd_sc_hd__or3_1
XFILLER_185_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19034_ _16854_/X _20835_/Q _19046_/S vssd1 vssd1 vccd1 vccd1 _19942_/D sky130_fd_sc_hd__mux2_1
XFILLER_185_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16246_ _16465_/B vssd1 vssd1 vccd1 vccd1 _16344_/B sky130_fd_sc_hd__buf_1
XANTENNA__13002__A1 _20691_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13458_ _13481_/A vssd1 vssd1 vccd1 vccd1 _13458_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__18034__B _18078_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12409_ _12409_/A vssd1 vssd1 vccd1 vccd1 _12417_/B sky130_fd_sc_hd__inv_2
XANTENNA__11013__B1 _10985_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16177_ _19447_/Q _16173_/X _16147_/X _16174_/X vssd1 vssd1 vccd1 vccd1 _19447_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17819__A2 _17232_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20125__CLK _21452_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput105 _17587_/Y vssd1 vssd1 vccd1 vccd1 HRDATA[4] sky130_fd_sc_hd__clkbuf_2
X_13389_ _13416_/A vssd1 vssd1 vccd1 vccd1 _13410_/A sky130_fd_sc_hd__buf_1
XFILLER_115_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput116 _18118_/LO vssd1 vssd1 vccd1 vccd1 IRQ[13] sky130_fd_sc_hd__clkbuf_2
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput127 _17090_/X vssd1 vssd1 vccd1 vccd1 IRQ[9] sky130_fd_sc_hd__clkbuf_2
XFILLER_99_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12761__B1 _12651_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput138 _18121_/LO vssd1 vssd1 vccd1 vccd1 scl_o_S4 sky130_fd_sc_hd__clkbuf_2
X_15128_ _15128_/A vssd1 vssd1 vccd1 vccd1 _15128_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_3_3_0_HCLK clkbuf_3_3_0_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_7_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_141_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15059_ _15059_/A _15059_/B vssd1 vssd1 vccd1 vccd1 _15214_/A sky130_fd_sc_hd__or2_2
X_19936_ _20159_/CLK _19936_/D repeater251/X vssd1 vssd1 vccd1 vccd1 _19936_/Q sky130_fd_sc_hd__dfrtp_1
X_19867_ _21183_/CLK _19867_/D repeater216/X vssd1 vssd1 vccd1 vccd1 _19867_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_122_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12810__B _13104_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09620_ _09657_/A vssd1 vssd1 vccd1 vccd1 _09620_/X sky130_fd_sc_hd__buf_1
X_18818_ _18817_/X _15115_/Y _18906_/S vssd1 vssd1 vccd1 vccd1 _18818_/X sky130_fd_sc_hd__mux2_2
XFILLER_244_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14266__B1 _13704_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19798_ _19820_/CLK _19798_/D vssd1 vssd1 vccd1 vccd1 _19798_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_209_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18749_ _17541_/Y _20638_/Q _18849_/S vssd1 vssd1 vccd1 vccd1 _18749_/X sky130_fd_sc_hd__mux2_1
XFILLER_237_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18196__S _18891_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20711_ _21367_/CLK _20711_/D repeater254/X vssd1 vssd1 vccd1 vccd1 _20711_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18924__S _18929_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20642_ _20657_/CLK _20642_/D repeater198/X vssd1 vssd1 vccd1 vccd1 _20642_/Q sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_56_HCLK clkbuf_4_12_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _21342_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_149_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20573_ _20946_/CLK _20573_/D repeater266/X vssd1 vssd1 vccd1 vccd1 _20573_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_177_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18180__A1 _13917_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20427__RESET_B repeater270/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20080__RESET_B repeater259/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21125_ _21125_/CLK _21125_/D repeater237/X vssd1 vssd1 vccd1 vccd1 _21125_/Q sky130_fd_sc_hd__dfrtp_1
X_21056_ _21147_/CLK _21056_/D repeater215/X vssd1 vssd1 vccd1 vccd1 _21056_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_132_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20007_ _21223_/CLK _20007_/D repeater238/X vssd1 vssd1 vccd1 vccd1 _20007_/Q sky130_fd_sc_hd__dfrtp_1
X_09818_ _15865_/A vssd1 vssd1 vccd1 vccd1 _09818_/X sky130_fd_sc_hd__buf_1
XFILLER_246_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__21286__RESET_B repeater207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17994__A1 _18344_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_234_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09749_ _11058_/A _20153_/Q _09744_/X _09745_/Y _09748_/X vssd1 vssd1 vccd1 vccd1
+ _09768_/A sky130_fd_sc_hd__o221a_1
XANTENNA__12807__A1 _20774_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12760_ _12778_/A vssd1 vssd1 vccd1 vccd1 _12760_/X sky130_fd_sc_hd__buf_1
XFILLER_160_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ _17553_/A vssd1 vssd1 vccd1 vccd1 _14256_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_242_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20909_ _20915_/CLK _20909_/D repeater218/X vssd1 vssd1 vccd1 vccd1 _20909_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12691_ _20824_/Q _12686_/X _09649_/X _12688_/X vssd1 vssd1 vccd1 vccd1 _20824_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18834__S _18930_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14430_ _21480_/Q vssd1 vssd1 vccd1 vccd1 _14430_/Y sky130_fd_sc_hd__inv_2
XPHY_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11642_ _11646_/A vssd1 vssd1 vccd1 vccd1 _11642_/X sky130_fd_sc_hd__clkbuf_2
XPHY_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14361_ _14503_/A _14502_/A _14361_/C _14504_/A vssd1 vssd1 vccd1 vccd1 _14362_/D
+ sky130_fd_sc_hd__or4_4
XFILLER_168_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11573_ _11743_/A vssd1 vssd1 vccd1 vccd1 _11573_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16100_ _19482_/Q _16094_/X _15873_/X _16096_/X vssd1 vssd1 vccd1 vccd1 _19482_/D
+ sky130_fd_sc_hd__a22o_1
Xinput18 HADDR[25] vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__buf_1
XPHY_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13312_ _20539_/Q _13307_/X _13311_/X _13308_/X vssd1 vssd1 vccd1 vccd1 _20539_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_167_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10524_ _10785_/A vssd1 vssd1 vccd1 vccd1 _10827_/A sky130_fd_sc_hd__buf_1
Xinput29 HADDR[6] vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__buf_1
XANTENNA__20850__RESET_B repeater243/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17080_ _17080_/A vssd1 vssd1 vccd1 vccd1 _18079_/A sky130_fd_sc_hd__buf_1
X_14292_ _20127_/Q vssd1 vssd1 vccd1 vccd1 _14292_/X sky130_fd_sc_hd__buf_1
XPHY_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16031_ _19520_/Q _16028_/X _15772_/X _16029_/X vssd1 vssd1 vccd1 vccd1 _19520_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__20168__RESET_B repeater190/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13243_ _14262_/A vssd1 vssd1 vccd1 vccd1 _13243_/X sky130_fd_sc_hd__buf_2
X_10455_ _21303_/Q vssd1 vssd1 vccd1 vccd1 _10779_/A sky130_fd_sc_hd__inv_2
XFILLER_184_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13174_ _20599_/Q _13165_/X _13173_/X _13167_/X vssd1 vssd1 vccd1 vccd1 _20599_/D
+ sky130_fd_sc_hd__a22o_1
X_10386_ _21365_/Q _10385_/Y _10373_/X _10281_/B vssd1 vssd1 vccd1 vccd1 _21365_/D
+ sky130_fd_sc_hd__o211a_1
X_12125_ _20369_/Q vssd1 vssd1 vccd1 vccd1 _12125_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17982_ _17982_/A _18001_/B vssd1 vssd1 vccd1 vccd1 _17982_/Y sky130_fd_sc_hd__nor2_1
X_19721_ _19774_/CLK _19721_/D vssd1 vssd1 vccd1 vccd1 _19721_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12056_ _20957_/Q vssd1 vssd1 vccd1 vccd1 _12311_/A sky130_fd_sc_hd__inv_2
X_16933_ _19962_/Q vssd1 vssd1 vccd1 vccd1 _16933_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11007_ _21013_/Q vssd1 vssd1 vccd1 vccd1 _15413_/A sky130_fd_sc_hd__inv_2
X_19652_ _19820_/CLK _19652_/D vssd1 vssd1 vccd1 vccd1 _19652_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16864_ _16862_/Y _16863_/Y _16848_/X vssd1 vssd1 vccd1 vccd1 _16864_/X sky130_fd_sc_hd__o21a_1
XFILLER_203_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18603_ _17830_/X _09731_/Y _18928_/S vssd1 vssd1 vccd1 vccd1 _18603_/X sky130_fd_sc_hd__mux2_1
X_15815_ _15815_/A _20134_/Q _16484_/B vssd1 vssd1 vccd1 vccd1 _16419_/C sky130_fd_sc_hd__or3_4
X_16795_ _16795_/A _16795_/B vssd1 vssd1 vccd1 vccd1 _16795_/Y sky130_fd_sc_hd__nor2_1
X_19583_ _21021_/CLK _19583_/D vssd1 vssd1 vccd1 vccd1 _19583_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_225_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_219_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17214__A _18045_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15746_ _19653_/Q _15743_/X _15725_/X _15745_/X vssd1 vssd1 vccd1 vccd1 _19653_/D
+ sky130_fd_sc_hd__a22o_1
X_18534_ _18533_/X _20276_/Q _18904_/S vssd1 vssd1 vccd1 vccd1 _18534_/X sky130_fd_sc_hd__mux2_1
XANTENNA__19282__S0 _19285_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12958_ _20708_/Q _12948_/X _12957_/X _12951_/X vssd1 vssd1 vccd1 vccd1 _20708_/D
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_79_HCLK clkbuf_4_13_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20623_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__17737__B2 _17728_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18029__B _18032_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11909_ _15559_/A _11909_/B vssd1 vssd1 vccd1 vccd1 _11910_/B sky130_fd_sc_hd__or2_1
XFILLER_233_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15677_ _19685_/Q _15674_/X _15657_/X _15676_/X vssd1 vssd1 vccd1 vccd1 _19685_/D
+ sky130_fd_sc_hd__a22o_1
X_18465_ _18464_/X _21291_/Q _18617_/S vssd1 vssd1 vccd1 vccd1 _18465_/X sky130_fd_sc_hd__mux2_1
X_12889_ _12809_/X _20737_/Q _12889_/S vssd1 vssd1 vccd1 vccd1 _20737_/D sky130_fd_sc_hd__mux2_1
XANTENNA__18744__S _18841_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14628_ _20191_/Q _14627_/Y _14624_/X _14581_/B vssd1 vssd1 vccd1 vccd1 _20191_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__20938__RESET_B repeater278/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17416_ _19385_/Q vssd1 vssd1 vccd1 vccd1 _17416_/Y sky130_fd_sc_hd__inv_2
X_18396_ _18845_/A0 _10443_/Y _18896_/S vssd1 vssd1 vccd1 vccd1 _18396_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17347_ _19584_/Q vssd1 vssd1 vccd1 vccd1 _17348_/A sky130_fd_sc_hd__inv_2
X_14559_ _20137_/Q vssd1 vssd1 vccd1 vccd1 _16077_/A sky130_fd_sc_hd__inv_2
XFILLER_159_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18045__A _18045_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17278_ _17370_/A vssd1 vssd1 vccd1 vccd1 _17449_/A sky130_fd_sc_hd__buf_1
XFILLER_146_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16229_ _16325_/A _16229_/B _16229_/C vssd1 vssd1 vccd1 vccd1 _16240_/A sky130_fd_sc_hd__or3_4
X_19017_ _16924_/X _20406_/Q _19019_/S vssd1 vssd1 vccd1 vccd1 _19959_/D sky130_fd_sc_hd__mux2_1
XANTENNA__19111__A0 _17064_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11537__A1 _21138_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12821__A _12841_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19919_ _21379_/CLK _19919_/D repeater213/X vssd1 vssd1 vccd1 vccd1 _19919_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_69_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_216_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09603_ _10975_/A vssd1 vssd1 vccd1 vccd1 _14304_/A sky130_fd_sc_hd__buf_2
XFILLER_84_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19273__S0 _19275_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_224_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18654__S _18908_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_104_HCLK_A clkbuf_4_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10597__A2_N _20762_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_167_HCLK_A clkbuf_opt_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20625_ _20697_/CLK _20625_/D repeater193/X vssd1 vssd1 vccd1 vccd1 _20625_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_rebuffer3_A _20027_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10579__A2 _20742_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20556_ _20592_/CLK _20556_/D repeater260/X vssd1 vssd1 vccd1 vccd1 _20556_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_192_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20261__RESET_B repeater264/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20487_ _20937_/CLK _20487_/D repeater277/X vssd1 vssd1 vccd1 vccd1 _20487_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_138_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10240_ _21363_/Q vssd1 vssd1 vccd1 vccd1 _10278_/A sky130_fd_sc_hd__inv_2
XFILLER_105_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10171_ _21404_/Q _10169_/X _10170_/X _10164_/A vssd1 vssd1 vccd1 vccd1 _21404_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__21467__RESET_B repeater205/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21108_ _21424_/CLK _21108_/D repeater230/X vssd1 vssd1 vccd1 vccd1 _21108_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_154_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18829__S _18930_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13930_ _13922_/X _13930_/B _13930_/C _13930_/D vssd1 vssd1 vccd1 vccd1 _13962_/B
+ sky130_fd_sc_hd__and4b_1
XFILLER_47_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21039_ _21401_/CLK _21039_/D repeater242/X vssd1 vssd1 vccd1 vccd1 _21039_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_208_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13861_ _20295_/Q vssd1 vssd1 vccd1 vccd1 _14011_/A sky130_fd_sc_hd__inv_2
XFILLER_170_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15600_ _19724_/Q _15596_/X _15473_/X _15598_/X vssd1 vssd1 vccd1 vccd1 _19724_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_216_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12812_ _20771_/Q vssd1 vssd1 vccd1 vccd1 _16779_/A sky130_fd_sc_hd__buf_2
X_16580_ _16580_/A vssd1 vssd1 vccd1 vccd1 _19917_/D sky130_fd_sc_hd__inv_2
XFILLER_170_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13792_ _20620_/Q _14586_/A _20616_/Q _14582_/A _13791_/X vssd1 vssd1 vccd1 vccd1
+ _13811_/A sky130_fd_sc_hd__o221a_1
XANTENNA__19264__S0 _19275_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15531_ _15537_/A vssd1 vssd1 vccd1 vccd1 _15531_/X sky130_fd_sc_hd__buf_1
X_12743_ _12743_/A _12743_/B _18971_/X _18975_/X vssd1 vssd1 vccd1 vccd1 _12743_/X
+ sky130_fd_sc_hd__or4b_4
XFILLER_31_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18564__S _18680_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_242_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18250_ _17976_/Y _20453_/Q _18784_/S vssd1 vssd1 vccd1 vccd1 _18250_/X sky130_fd_sc_hd__mux2_1
XFILLER_63_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15462_ _19784_/Q _15459_/X _15427_/X _15460_/X vssd1 vssd1 vccd1 vccd1 _19784_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_188_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12674_ _12680_/A vssd1 vssd1 vccd1 vccd1 _12674_/X sky130_fd_sc_hd__buf_1
XPHY_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17201_ _17201_/A vssd1 vssd1 vccd1 vccd1 _17575_/A sky130_fd_sc_hd__buf_1
X_14413_ _14409_/Y _20211_/Q _14410_/Y _20028_/Q _14412_/X vssd1 vssd1 vccd1 vccd1
+ _14420_/C sky130_fd_sc_hd__o221a_1
Xclkbuf_leaf_8_HCLK clkbuf_opt_2_HCLK/A vssd1 vssd1 vccd1 vccd1 _21222_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11625_ _21109_/Q _11625_/B _14813_/C vssd1 vssd1 vccd1 vccd1 _11638_/A sky130_fd_sc_hd__or3b_4
XPHY_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11216__B1 _09659_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18181_ _18180_/X _14088_/A _18904_/S vssd1 vssd1 vccd1 vccd1 _18181_/X sky130_fd_sc_hd__mux2_1
XPHY_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15393_ _19815_/Q _15389_/X _15352_/X _15390_/X vssd1 vssd1 vccd1 vccd1 _19815_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_26_HCLK_A clkbuf_opt_4_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17132_ _19309_/Q _17369_/B vssd1 vssd1 vccd1 vccd1 _17132_/Y sky130_fd_sc_hd__nor2_1
XPHY_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12964__B1 _12881_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14344_ _20222_/Q vssd1 vssd1 vccd1 vccd1 _14460_/C sky130_fd_sc_hd__inv_2
XFILLER_184_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11556_ _21133_/Q _11552_/X _10886_/X _11554_/X vssd1 vssd1 vccd1 vccd1 _21133_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_89_HCLK_A clkbuf_4_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17063_ _16548_/A _17062_/Y _16585_/A vssd1 vssd1 vccd1 vccd1 _19877_/D sky130_fd_sc_hd__o21ai_1
X_10507_ _20693_/Q vssd1 vssd1 vccd1 vccd1 _10507_/Y sky130_fd_sc_hd__inv_2
XFILLER_183_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14275_ _20242_/Q vssd1 vssd1 vccd1 vccd1 _14275_/Y sky130_fd_sc_hd__inv_2
X_11487_ _19111_/X vssd1 vssd1 vccd1 vccd1 _11487_/X sky130_fd_sc_hd__buf_1
XFILLER_137_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16014_ _16340_/A vssd1 vssd1 vccd1 vccd1 _16014_/X sky130_fd_sc_hd__clkbuf_2
X_13226_ _13248_/A vssd1 vssd1 vccd1 vccd1 _13226_/X sky130_fd_sc_hd__buf_1
XFILLER_170_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10438_ _21306_/Q _18082_/A _10777_/A _20690_/Q vssd1 vssd1 vccd1 vccd1 _10438_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_170_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17209__A _17209_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13157_ _20607_/Q _13150_/X _13032_/X _13152_/X vssd1 vssd1 vccd1 vccd1 _20607_/D
+ sky130_fd_sc_hd__a22o_1
X_10369_ _10369_/A vssd1 vssd1 vccd1 vccd1 _10369_/Y sky130_fd_sc_hd__inv_2
X_12108_ _20954_/Q vssd1 vssd1 vccd1 vccd1 _12308_/A sky130_fd_sc_hd__inv_2
XANTENNA__13456__B _13456_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17965_ _18524_/X _17931_/X _18201_/X _17932_/X _17964_/X vssd1 vssd1 vccd1 vccd1
+ _17966_/C sky130_fd_sc_hd__o221a_1
XFILLER_100_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13088_ _20645_/Q _13086_/X _12860_/X _13087_/X vssd1 vssd1 vccd1 vccd1 _20645_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18739__S _18930_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19704_ _19706_/CLK _19704_/D vssd1 vssd1 vccd1 vccd1 _19704_/Q sky130_fd_sc_hd__dfxtp_1
X_16916_ _16913_/Y _16914_/Y _16915_/X vssd1 vssd1 vccd1 vccd1 _16916_/X sky130_fd_sc_hd__o21a_1
X_12039_ _20950_/Q vssd1 vssd1 vccd1 vccd1 _12304_/A sky130_fd_sc_hd__inv_2
XFILLER_238_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17896_ _17896_/A _17898_/B vssd1 vssd1 vccd1 vccd1 _17896_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__13692__A1 _20344_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09950__A _09957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_238_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19635_ _20142_/CLK _19635_/D vssd1 vssd1 vccd1 vccd1 _19635_/Q sky130_fd_sc_hd__dfxtp_1
X_16847_ _19941_/Q vssd1 vssd1 vccd1 vccd1 _16847_/Y sky130_fd_sc_hd__inv_2
XFILLER_226_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13472__A _13481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_241_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19255__S0 _19275_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19566_ _19812_/CLK _19566_/D vssd1 vssd1 vccd1 vccd1 _19566_/Q sky130_fd_sc_hd__dfxtp_1
X_16778_ _16778_/A _16778_/B vssd1 vssd1 vccd1 vccd1 _16778_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__18907__A0 _18906_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19886__SET_B repeater217/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18517_ _18516_/X _21294_/Q _18617_/S vssd1 vssd1 vccd1 vccd1 _18517_/X sky130_fd_sc_hd__mux2_1
XFILLER_80_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15729_ input66/X vssd1 vssd1 vccd1 vccd1 _16235_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__18474__S _18898_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19497_ _20326_/CLK _19497_/D vssd1 vssd1 vccd1 vccd1 _19497_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18448_ _18447_/X _10768_/A _18841_/S vssd1 vssd1 vccd1 vccd1 _18448_/X sky130_fd_sc_hd__mux2_1
XFILLER_194_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_221_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20701__RESET_B repeater190/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18379_ _17281_/X _17779_/Y _18835_/S vssd1 vssd1 vccd1 vccd1 _18379_/X sky130_fd_sc_hd__mux2_1
X_20410_ _20413_/CLK _20410_/D repeater185/X vssd1 vssd1 vccd1 vccd1 _20410_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12955__B1 _12954_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21390_ _21390_/CLK _21390_/D repeater240/X vssd1 vssd1 vccd1 vccd1 _21390_/Q sky130_fd_sc_hd__dfrtp_1
X_20341_ _20951_/CLK _20341_/D repeater269/X vssd1 vssd1 vccd1 vccd1 _20341_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_162_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20272_ _20724_/CLK _20272_/D repeater264/X vssd1 vssd1 vccd1 vccd1 _20272_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__13380__B1 _13169_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20003__SET_B repeater190/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18649__S _18907_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_229_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_245_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09639__B1 _09638_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19246__S0 _21005_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_231_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18384__S _18908_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_231_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16693__A _16720_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13199__B1 _12993_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12726__A _12898_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11410_ _11410_/A _11410_/B _11410_/C vssd1 vssd1 vccd1 vccd1 _11786_/C sky130_fd_sc_hd__or3_1
XFILLER_166_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12946__B1 _12697_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20608_ _20622_/CLK _20608_/D repeater195/X vssd1 vssd1 vccd1 vccd1 _20608_/Q sky130_fd_sc_hd__dfrtp_1
X_12390_ _12073_/X _12389_/Y _12359_/A _12306_/B vssd1 vssd1 vccd1 vccd1 _20951_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_123_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11341_ _11357_/A _11341_/B vssd1 vssd1 vccd1 vccd1 _11342_/A sky130_fd_sc_hd__or2_2
X_20539_ _20592_/CLK _20539_/D repeater267/X vssd1 vssd1 vccd1 vccd1 _20539_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_165_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14060_ _20268_/Q vssd1 vssd1 vccd1 vccd1 _14103_/A sky130_fd_sc_hd__inv_2
X_11272_ _11272_/A _11272_/B vssd1 vssd1 vccd1 vccd1 _11545_/B sky130_fd_sc_hd__nand2_1
XFILLER_152_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13011_ _20686_/Q _13005_/X _12922_/X _13007_/X vssd1 vssd1 vccd1 vccd1 _20686_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13557__A input54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10223_ _10223_/A _10223_/B _10227_/C vssd1 vssd1 vccd1 vccd1 _21379_/D sky130_fd_sc_hd__nor3_1
XANTENNA_input43_A HWDATA[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10154_ _10154_/A _10190_/A vssd1 vssd1 vccd1 vccd1 _10155_/B sky130_fd_sc_hd__or2_1
XFILLER_79_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18559__S _18680_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13123__B1 _12999_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21230__RESET_B repeater249/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14962_ _14962_/A _14962_/B _14962_/C _14962_/D vssd1 vssd1 vccd1 vccd1 _14963_/B
+ sky130_fd_sc_hd__or4_4
X_17750_ _19717_/Q vssd1 vssd1 vccd1 vccd1 _17750_/Y sky130_fd_sc_hd__inv_2
XFILLER_248_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10085_ _20784_/Q vssd1 vssd1 vccd1 vccd1 _10085_/Y sky130_fd_sc_hd__inv_2
XFILLER_248_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16701_ _19895_/Q _14235_/B _14236_/B vssd1 vssd1 vccd1 vccd1 _16701_/X sky130_fd_sc_hd__a21bo_1
XFILLER_235_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13913_ _20660_/Q _13893_/C _20644_/Q _14017_/A _13912_/X vssd1 vssd1 vccd1 vccd1
+ _13914_/D sky130_fd_sc_hd__o221a_1
X_14893_ _20590_/Q _14965_/A _20579_/Q _14845_/A vssd1 vssd1 vccd1 vccd1 _14893_/X
+ sky130_fd_sc_hd__o22a_1
X_17681_ _19404_/Q vssd1 vssd1 vccd1 vccd1 _17681_/Y sky130_fd_sc_hd__inv_2
XFILLER_208_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19420_ _19828_/CLK _19420_/D vssd1 vssd1 vccd1 vccd1 _19420_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16632_ _16632_/A _16632_/B _16632_/C vssd1 vssd1 vccd1 vccd1 _19843_/D sky130_fd_sc_hd__nor3_1
XFILLER_63_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13844_ _20316_/Q vssd1 vssd1 vccd1 vccd1 _13893_/A sky130_fd_sc_hd__inv_2
XFILLER_223_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19237__S0 _20130_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19351_ _19961_/CLK _19351_/D vssd1 vssd1 vccd1 vccd1 _19351_/Q sky130_fd_sc_hd__dfxtp_1
X_16563_ _16583_/A _16539_/A _16561_/Y _16547_/Y _16562_/X vssd1 vssd1 vccd1 vccd1
+ _16564_/B sky130_fd_sc_hd__o32a_1
X_13775_ _20618_/Q vssd1 vssd1 vccd1 vccd1 _13775_/Y sky130_fd_sc_hd__inv_2
X_10987_ _15653_/A vssd1 vssd1 vccd1 vccd1 _15375_/A sky130_fd_sc_hd__buf_1
XANTENNA__18294__S _18904_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_231_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18302_ _18301_/X _16830_/A _18667_/S vssd1 vssd1 vccd1 vccd1 _18302_/X sky130_fd_sc_hd__mux2_1
XFILLER_200_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12726_ _12898_/A _17153_/A vssd1 vssd1 vccd1 vccd1 _13329_/A sky130_fd_sc_hd__or2_2
X_15514_ _15785_/A vssd1 vssd1 vccd1 vccd1 _15514_/X sky130_fd_sc_hd__buf_1
XFILLER_204_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16494_ _16516_/A _16681_/B vssd1 vssd1 vccd1 vccd1 _16494_/X sky130_fd_sc_hd__or2_2
XFILLER_203_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19282_ _19685_/Q _19813_/Q _19805_/Q _19797_/Q _19285_/S0 _21017_/Q vssd1 vssd1
+ vccd1 vccd1 _19282_/X sky130_fd_sc_hd__mux4_2
XFILLER_188_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18233_ _20857_/Q input6/X _18236_/S vssd1 vssd1 vccd1 vccd1 _18233_/X sky130_fd_sc_hd__mux2_1
X_15445_ _19791_/Q _15441_/X _15429_/X _15442_/X vssd1 vssd1 vccd1 vccd1 _19791_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12657_ _20841_/Q _12650_/X _12656_/X _12654_/X vssd1 vssd1 vccd1 vccd1 _20841_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_150_HCLK_A clkbuf_opt_1_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11608_ _18992_/X _11598_/A _21114_/Q _11605_/X vssd1 vssd1 vccd1 vccd1 _21114_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_30_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15376_ _15389_/A vssd1 vssd1 vccd1 vccd1 _15376_/X sky130_fd_sc_hd__buf_1
X_18164_ _18163_/X _13904_/Y _18903_/S vssd1 vssd1 vccd1 vccd1 _18164_/X sky130_fd_sc_hd__mux2_1
X_12588_ _12600_/A vssd1 vssd1 vccd1 vccd1 _12588_/X sky130_fd_sc_hd__buf_1
Xclkbuf_leaf_109_HCLK clkbuf_opt_3_HCLK/A vssd1 vssd1 vccd1 vccd1 _20075_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14327_ _20235_/Q vssd1 vssd1 vccd1 vccd1 _14328_/A sky130_fd_sc_hd__inv_2
X_17115_ _19446_/Q vssd1 vssd1 vccd1 vccd1 _17115_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14273__D _14273_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11539_ _21136_/Q _11534_/X _10900_/X _11535_/X vssd1 vssd1 vccd1 vccd1 _21136_/D
+ sky130_fd_sc_hd__a22o_1
X_18095_ _18645_/X _17862_/A _18651_/X _18065_/X vssd1 vssd1 vccd1 vccd1 _18095_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_209_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17046_ _17046_/A _17046_/B vssd1 vssd1 vccd1 vccd1 _19842_/D sky130_fd_sc_hd__and2_1
X_14258_ _14258_/A vssd1 vssd1 vccd1 vccd1 _14258_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__18042__B _18042_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13467__A _13483_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13209_ input52/X vssd1 vssd1 vccd1 vccd1 _13209_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__13362__B1 _13144_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14189_ _14093_/A _14093_/B _14187_/Y _14215_/B vssd1 vssd1 vccd1 vccd1 _20283_/D
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__18469__S _18898_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18997_ _17010_/X _20426_/Q _19026_/S vssd1 vssd1 vccd1 vccd1 _19979_/D sky130_fd_sc_hd__mux2_1
XFILLER_97_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater202 repeater203/X vssd1 vssd1 vccd1 vccd1 repeater202/X sky130_fd_sc_hd__buf_8
XFILLER_140_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater213 repeater215/X vssd1 vssd1 vccd1 vccd1 repeater213/X sky130_fd_sc_hd__buf_8
X_17948_ _18064_/A vssd1 vssd1 vccd1 vccd1 _17948_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_227_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater224 repeater226/X vssd1 vssd1 vccd1 vccd1 repeater224/X sky130_fd_sc_hd__buf_8
XANTENNA__13665__A1 _20361_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater235 repeater237/X vssd1 vssd1 vccd1 vccd1 repeater235/X sky130_fd_sc_hd__buf_8
Xrepeater246 repeater247/X vssd1 vssd1 vccd1 vccd1 repeater246/X sky130_fd_sc_hd__buf_6
XFILLER_39_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09680__A input65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater257 repeater268/X vssd1 vssd1 vccd1 vccd1 repeater257/X sky130_fd_sc_hd__buf_8
Xrepeater268 repeater269/X vssd1 vssd1 vccd1 vccd1 repeater268/X sky130_fd_sc_hd__buf_6
XFILLER_66_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17879_ _18501_/X _17857_/X _18492_/X _17869_/X vssd1 vssd1 vccd1 vccd1 _17879_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_238_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater279 repeater280/X vssd1 vssd1 vccd1 vccd1 repeater279/X sky130_fd_sc_hd__buf_6
XFILLER_65_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20953__RESET_B repeater187/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19618_ _21449_/CLK _19618_/D vssd1 vssd1 vccd1 vccd1 _19618_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19228__S0 _20130_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20890_ _20890_/CLK _20890_/D repeater185/X vssd1 vssd1 vccd1 vccd1 _20890_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_38_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19549_ _19789_/CLK _19549_/D vssd1 vssd1 vccd1 vccd1 _19549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21442_ _21445_/CLK _21442_/D repeater245/X vssd1 vssd1 vccd1 vccd1 _21442_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_181_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12980__S _12980_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21373_ _21375_/CLK _21373_/D repeater257/X vssd1 vssd1 vccd1 vccd1 _21373_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA_clkbuf_leaf_72_HCLK_A clkbuf_opt_7_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20324_ _20326_/CLK _20324_/D repeater250/X vssd1 vssd1 vccd1 vccd1 _20324_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_116_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12156__B2 _20344_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13353__B1 _13216_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20255_ _20256_/CLK _20255_/D repeater217/X vssd1 vssd1 vccd1 vccd1 _20255_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_103_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20186_ _21483_/CLK _20186_/D repeater193/X vssd1 vssd1 vccd1 vccd1 _20186_/Q sky130_fd_sc_hd__dfrtp_1
X_09997_ _20020_/Q _10013_/A _09985_/A vssd1 vssd1 vccd1 vccd1 _17036_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__18379__S _18835_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15592__A _15592_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10910_ _09931_/X _21246_/Q _10910_/S vssd1 vssd1 vccd1 vccd1 _21246_/D sky130_fd_sc_hd__mux2_1
XFILLER_205_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20694__RESET_B repeater193/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19219__S0 _20130_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11890_ _11885_/A _11885_/B _11886_/A _11889_/X vssd1 vssd1 vccd1 vccd1 _11890_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_71_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_232_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10841_ _21277_/Q _10677_/A _10812_/A _10839_/A vssd1 vssd1 vccd1 vccd1 _21277_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_44_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19003__S _19019_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13560_ input53/X vssd1 vssd1 vccd1 vccd1 _13560_/X sky130_fd_sc_hd__buf_4
XFILLER_240_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10772_ _10772_/A _10807_/A vssd1 vssd1 vccd1 vccd1 _10773_/B sky130_fd_sc_hd__or2_2
XFILLER_197_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12511_ _19908_/Q _12515_/A vssd1 vssd1 vccd1 vccd1 _12511_/Y sky130_fd_sc_hd__nor2_1
XFILLER_201_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13491_ _13491_/A vssd1 vssd1 vccd1 vccd1 _13514_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18842__S _18896_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15230_ _18001_/A _20066_/Q _20487_/Q _15129_/X vssd1 vssd1 vccd1 vccd1 _15230_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_9_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12919__B1 _12918_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12442_ _20944_/Q _12437_/C _12438_/X _12440_/A vssd1 vssd1 vccd1 vccd1 _20944_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_100_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17966__B _17966_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21134__CLK _21134_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13592__B1 _13511_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15161_ _20075_/Q _15089_/Y _15090_/Y _15089_/A _15160_/X vssd1 vssd1 vccd1 vccd1
+ _20075_/D sky130_fd_sc_hd__o221a_1
X_12373_ _12373_/A vssd1 vssd1 vccd1 vccd1 _12373_/X sky130_fd_sc_hd__buf_1
XANTENNA__21482__RESET_B repeater200/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14112_ _20557_/Q vssd1 vssd1 vccd1 vccd1 _14112_/Y sky130_fd_sc_hd__inv_2
X_11324_ _19870_/Q vssd1 vssd1 vccd1 vccd1 _15310_/A sky130_fd_sc_hd__buf_1
XFILLER_5_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15333__A1 _20025_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15092_ _20053_/Q vssd1 vssd1 vccd1 vccd1 _15092_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_114_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13344__B1 _13284_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13287__A input53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14043_ _20285_/Q vssd1 vssd1 vccd1 vccd1 _14095_/A sky130_fd_sc_hd__inv_2
X_18920_ _18919_/X _21268_/Q _18920_/S vssd1 vssd1 vccd1 vccd1 _18920_/X sky130_fd_sc_hd__mux2_1
X_11255_ _19066_/X _11250_/X _21186_/Q _11251_/X vssd1 vssd1 vccd1 vccd1 _21186_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_107_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10206_ _10206_/A _10210_/A vssd1 vssd1 vccd1 vccd1 _10207_/B sky130_fd_sc_hd__or2_2
X_18851_ _17079_/Y _15234_/Y _18908_/S vssd1 vssd1 vccd1 vccd1 _18851_/X sky130_fd_sc_hd__mux2_1
X_11186_ _11179_/X _11180_/X _11186_/S vssd1 vssd1 vccd1 vccd1 _21218_/D sky130_fd_sc_hd__mux2_1
XFILLER_121_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18289__S _18680_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17802_ _18395_/X _17839_/A _18392_/X _17869_/A _17801_/X vssd1 vssd1 vccd1 vccd1
+ _17802_/X sky130_fd_sc_hd__o221a_2
X_10137_ _10137_/A _10137_/B _10137_/C _10137_/D vssd1 vssd1 vccd1 vccd1 _10185_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_122_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18782_ _18781_/X _14073_/A _18850_/S vssd1 vssd1 vccd1 vccd1 _18782_/X sky130_fd_sc_hd__mux2_1
XFILLER_209_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15994_ _15994_/A vssd1 vssd1 vccd1 vccd1 _15994_/X sky130_fd_sc_hd__buf_1
XFILLER_248_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17733_ _18700_/X _17401_/X _18703_/X _17226_/A vssd1 vssd1 vccd1 vccd1 _17733_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_94_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14945_ _20596_/Q vssd1 vssd1 vccd1 vccd1 _14945_/Y sky130_fd_sc_hd__inv_2
X_10068_ _10152_/A _10151_/A _10068_/C _10068_/D vssd1 vssd1 vccd1 vccd1 _10075_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_235_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17664_ _12606_/A _17656_/X _17658_/X _17661_/X _17663_/X vssd1 vssd1 vccd1 vccd1
+ _17664_/X sky130_fd_sc_hd__o2111a_1
X_14876_ _14963_/D _14876_/B vssd1 vssd1 vccd1 vccd1 _14977_/A sky130_fd_sc_hd__or2_1
XFILLER_211_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19403_ _21009_/CLK _19403_/D vssd1 vssd1 vccd1 vccd1 _19403_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_235_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16615_ _16585_/A _16558_/X _16614_/X vssd1 vssd1 vccd1 vccd1 _19988_/D sky130_fd_sc_hd__a21bo_1
X_13827_ _20201_/Q vssd1 vssd1 vccd1 vccd1 _14590_/A sky130_fd_sc_hd__inv_2
XFILLER_51_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17595_ _19411_/Q vssd1 vssd1 vccd1 vccd1 _17595_/Y sky130_fd_sc_hd__inv_2
X_19334_ _20172_/CLK _19334_/D vssd1 vssd1 vccd1 vccd1 _19334_/Q sky130_fd_sc_hd__dfxtp_1
X_16546_ _16546_/A vssd1 vssd1 vccd1 vccd1 _16738_/B sky130_fd_sc_hd__buf_1
X_13758_ _20183_/Q vssd1 vssd1 vccd1 vccd1 _14573_/A sky130_fd_sc_hd__inv_2
XFILLER_62_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18037__B _18084_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12709_ _20814_/Q _12707_/X _11736_/X _12708_/X vssd1 vssd1 vccd1 vccd1 _20814_/D
+ sky130_fd_sc_hd__a22o_1
X_19265_ _17248_/Y _17249_/Y _17250_/Y _17251_/Y _19275_/S0 _21004_/Q vssd1 vssd1
+ vccd1 vccd1 _19265_/X sky130_fd_sc_hd__mux4_2
X_13689_ _20347_/Q _13686_/X _12849_/A _13688_/X vssd1 vssd1 vccd1 vccd1 _20347_/D
+ sky130_fd_sc_hd__a22o_1
X_16477_ _19293_/Q _16473_/X _16293_/X _16474_/X vssd1 vssd1 vccd1 vccd1 _19293_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18752__S _18907_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18216_ _18215_/X _14090_/A _18904_/S vssd1 vssd1 vccd1 vccd1 _18216_/X sky130_fd_sc_hd__mux2_1
X_15428_ _19800_/Q _15423_/X _15427_/X _15425_/X vssd1 vssd1 vccd1 vccd1 _19800_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_176_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19196_ _19192_/X _19193_/X _19194_/X _19195_/X _20123_/Q _20124_/Q vssd1 vssd1 vccd1
+ vccd1 _19196_/X sky130_fd_sc_hd__mux4_2
XFILLER_163_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13583__B1 _13432_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15359_ _15366_/A vssd1 vssd1 vccd1 vccd1 _15359_/X sky130_fd_sc_hd__buf_1
X_18147_ _18146_/X _10280_/A _18886_/S vssd1 vssd1 vccd1 vccd1 _18147_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18078_ _18078_/A _18078_/B vssd1 vssd1 vccd1 vccd1 _18078_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__12813__B _13106_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13335__B1 _13265_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09920_ _09925_/A vssd1 vssd1 vccd1 vccd1 _09924_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_171_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17029_ _21251_/Q vssd1 vssd1 vccd1 vccd1 _17029_/Y sky130_fd_sc_hd__inv_2
XFILLER_236_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10614__A _20764_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20040_ _21183_/CLK _20040_/D repeater216/X vssd1 vssd1 vccd1 vccd1 _20040_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__18274__A0 _18273_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09851_ _10843_/B vssd1 vssd1 vccd1 vccd1 _09851_/X sky130_fd_sc_hd__buf_1
XANTENNA__18199__S _18667_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09782_ _21460_/Q _09781_/Y _09777_/X vssd1 vssd1 vccd1 vccd1 _21460_/D sky130_fd_sc_hd__o21a_1
XFILLER_105_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18927__S _18927_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_227_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20942_ _20950_/CLK _20942_/D repeater278/X vssd1 vssd1 vccd1 vccd1 _20942_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_4219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20873_ _21459_/CLK _20873_/D repeater244/X vssd1 vssd1 vccd1 vccd1 _20873_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_54_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13810__A1 _20609_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18662__S _18910_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21425_ _21429_/CLK _21425_/D repeater231/X vssd1 vssd1 vccd1 vccd1 _21425_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_163_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14118__A2 _20288_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21356_ _21367_/CLK _21356_/D repeater254/X vssd1 vssd1 vccd1 vccd1 _21356_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_135_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12723__B _13106_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13326__B1 _13173_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20307_ _20693_/CLK _20307_/D repeater196/X vssd1 vssd1 vccd1 vccd1 _20307_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_150_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21287_ _21306_/CLK _21287_/D repeater207/X vssd1 vssd1 vccd1 vccd1 _21287_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_146_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19970__RESET_B repeater184/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18265__A0 _18848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11040_ _16949_/B _11040_/B vssd1 vssd1 vccd1 vccd1 _16989_/B sky130_fd_sc_hd__or2_2
X_20238_ _21481_/CLK _20238_/D repeater205/X vssd1 vssd1 vccd1 vccd1 _20238_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_76_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20169_ _21125_/CLK _20169_/D repeater190/X vssd1 vssd1 vccd1 vccd1 _20169_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_190_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20804__RESET_B repeater252/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12991_ input59/X vssd1 vssd1 vccd1 vccd1 _12991_/X sky130_fd_sc_hd__buf_2
XFILLER_217_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18837__S _18879_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14730_ _17774_/B _14730_/B vssd1 vssd1 vccd1 vccd1 _14732_/A sky130_fd_sc_hd__or2_2
XFILLER_85_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11942_ _21010_/Q _11941_/X _21010_/Q _11941_/X vssd1 vssd1 vccd1 vccd1 _21010_/D
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_245_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14661_ _16484_/A _14661_/B vssd1 vssd1 vccd1 vccd1 _16482_/A sky130_fd_sc_hd__or2_1
X_11873_ _10934_/X _11816_/Y _11817_/X _11864_/X vssd1 vssd1 vccd1 vccd1 _21024_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_189_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13612_ _20392_/Q _13605_/X _13547_/X _13608_/X vssd1 vssd1 vccd1 vccd1 _20392_/D
+ sky130_fd_sc_hd__a22o_1
X_16400_ _16400_/A vssd1 vssd1 vccd1 vccd1 _16400_/X sky130_fd_sc_hd__buf_1
X_10824_ _10824_/A _10824_/B _10824_/C vssd1 vssd1 vccd1 vccd1 _21287_/D sky130_fd_sc_hd__nor3_1
XFILLER_72_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17380_ _21046_/Q vssd1 vssd1 vccd1 vccd1 _17380_/Y sky130_fd_sc_hd__inv_2
X_14592_ _14592_/A _14605_/A vssd1 vssd1 vccd1 vccd1 _14593_/B sky130_fd_sc_hd__or2_2
XFILLER_44_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12604__A2 _12600_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16331_ _19371_/Q _16326_/X _16237_/X _16328_/X vssd1 vssd1 vccd1 vccd1 _19371_/D
+ sky130_fd_sc_hd__a22o_1
X_13543_ input61/X vssd1 vssd1 vccd1 vccd1 _13543_/X sky130_fd_sc_hd__clkbuf_4
X_10755_ _10755_/A _10839_/A vssd1 vssd1 vccd1 vccd1 _10756_/B sky130_fd_sc_hd__or2_2
XANTENNA__12186__A _20341_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18572__S _18667_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19050_ _16784_/Y _20819_/Q _19058_/S vssd1 vssd1 vccd1 vccd1 _19926_/D sky130_fd_sc_hd__mux2_1
X_16262_ _16269_/A vssd1 vssd1 vccd1 vccd1 _16262_/X sky130_fd_sc_hd__buf_1
X_13474_ _20456_/Q _13472_/X _13287_/X _13473_/X vssd1 vssd1 vccd1 vccd1 _20456_/D
+ sky130_fd_sc_hd__a22o_1
X_10686_ _10659_/A _10659_/B _10685_/X _10683_/Y vssd1 vssd1 vccd1 vccd1 _21330_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_40_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12368__A1 _12036_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18001_ _18001_/A _18001_/B vssd1 vssd1 vccd1 vccd1 _18001_/Y sky130_fd_sc_hd__nor2_1
X_15213_ _15061_/A _15061_/B _15211_/Y _15179_/A vssd1 vssd1 vccd1 vccd1 _20046_/D
+ sky130_fd_sc_hd__a211oi_2
X_12425_ _12425_/A _12425_/B vssd1 vssd1 vccd1 vccd1 _12455_/A sky130_fd_sc_hd__or2_1
X_16193_ _20136_/Q vssd1 vssd1 vccd1 vccd1 _16419_/B sky130_fd_sc_hd__buf_1
X_15144_ _15131_/X _15144_/B _15144_/C _15144_/D vssd1 vssd1 vccd1 vccd1 _15144_/X
+ sky130_fd_sc_hd__and4b_1
X_12356_ _20971_/Q _12355_/Y _12344_/X _12325_/B vssd1 vssd1 vccd1 vccd1 _20971_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__13317__B1 _13240_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11307_ _11543_/A _11307_/B _11307_/C _11543_/C vssd1 vssd1 vccd1 vccd1 _11544_/A
+ sky130_fd_sc_hd__or4_4
X_15075_ _15075_/A _15188_/A vssd1 vssd1 vccd1 vccd1 _15076_/B sky130_fd_sc_hd__or2_2
X_19952_ _20809_/CLK _19952_/D repeater270/X vssd1 vssd1 vccd1 vccd1 _19952_/Q sky130_fd_sc_hd__dfrtp_1
X_12287_ _12396_/A _20501_/Q _12425_/A _20516_/Q vssd1 vssd1 vccd1 vccd1 _12287_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_206_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18256__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18903_ _18902_/X _13907_/Y _18903_/S vssd1 vssd1 vccd1 vccd1 _18903_/X sky130_fd_sc_hd__mux2_1
X_14026_ _14026_/A vssd1 vssd1 vccd1 vccd1 _14026_/Y sky130_fd_sc_hd__inv_2
X_11238_ _11250_/A vssd1 vssd1 vccd1 vccd1 _11251_/A sky130_fd_sc_hd__inv_2
XFILLER_106_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19883_ _21338_/CLK _19883_/D repeater221/X vssd1 vssd1 vccd1 vccd1 _19883_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_95_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18834_ _18833_/X _19256_/X _18930_/S vssd1 vssd1 vccd1 vccd1 _18834_/X sky130_fd_sc_hd__mux2_1
X_11169_ _11176_/A _15594_/A vssd1 vssd1 vccd1 vccd1 _11170_/A sky130_fd_sc_hd__or2_1
XANTENNA__20545__RESET_B repeater263/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18765_ _18764_/X _17505_/X _18929_/S vssd1 vssd1 vccd1 vccd1 _18765_/X sky130_fd_sc_hd__mux2_1
XANTENNA__18747__S _18897_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15977_ _19546_/Q _15968_/X _15941_/X _15971_/X vssd1 vssd1 vccd1 vccd1 _19546_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_209_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17716_ _21050_/Q vssd1 vssd1 vccd1 vccd1 _17716_/Y sky130_fd_sc_hd__inv_2
X_14928_ _14926_/Y _20083_/Q _20572_/Q _15003_/A _14927_/X vssd1 vssd1 vccd1 vccd1
+ _14933_/C sky130_fd_sc_hd__o221a_1
X_18696_ _18695_/X _15111_/Y _18906_/S vssd1 vssd1 vccd1 vccd1 _18696_/X sky130_fd_sc_hd__mux2_2
XFILLER_36_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17647_ _21132_/Q vssd1 vssd1 vccd1 vccd1 _17647_/Y sky130_fd_sc_hd__inv_2
X_14859_ _20085_/Q vssd1 vssd1 vccd1 vccd1 _15005_/A sky130_fd_sc_hd__inv_2
XANTENNA__18048__A _18048_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17578_ _18742_/X _17933_/A _18766_/X _17854_/A _17577_/Y vssd1 vssd1 vccd1 vccd1
+ _17578_/X sky130_fd_sc_hd__o221a_1
XFILLER_177_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19317_ _19961_/CLK _19317_/D vssd1 vssd1 vccd1 vccd1 _19317_/Q sky130_fd_sc_hd__dfxtp_1
X_16529_ _16519_/Y _16680_/B _19998_/Q vssd1 vssd1 vccd1 vccd1 _16688_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__11712__B _15312_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18482__S _18903_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19248_ _17354_/Y _17355_/Y _17356_/Y _17357_/Y _20130_/Q _20131_/Q vssd1 vssd1 vccd1
+ vccd1 _19248_/X sky130_fd_sc_hd__mux4_2
XANTENNA__21333__RESET_B repeater204/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13556__B1 _13555_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19179_ _19729_/Q _19369_/Q _19785_/Q _19769_/Q _19280_/S0 _20122_/Q vssd1 vssd1
+ vccd1 vccd1 _19179_/X sky130_fd_sc_hd__mux4_2
XANTENNA__12824__A _12842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18495__A0 _18494_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21210_ _21401_/CLK _21210_/D repeater241/X vssd1 vssd1 vccd1 vccd1 _21210_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_117_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21141_ _21141_/CLK _21141_/D repeater192/X vssd1 vssd1 vccd1 vccd1 _21141_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_160_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09903_ _09898_/X _09899_/X _09898_/X _09899_/X vssd1 vssd1 vccd1 vccd1 _09904_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_132_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21072_ _21424_/CLK _21072_/D repeater230/X vssd1 vssd1 vccd1 vccd1 _21072_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_116_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20023_ _21421_/CLK _20023_/D repeater232/X vssd1 vssd1 vccd1 vccd1 _20023_/Q sky130_fd_sc_hd__dfrtp_1
X_09834_ _21447_/Q vssd1 vssd1 vccd1 vccd1 _15881_/A sky130_fd_sc_hd__buf_1
XFILLER_246_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20286__RESET_B repeater262/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09765_ _20150_/Q vssd1 vssd1 vccd1 vccd1 _09765_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18657__S _18669_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14284__A1 _20123_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20215__RESET_B repeater202/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09696_ input49/X vssd1 vssd1 vccd1 vccd1 _15523_/A sky130_fd_sc_hd__clkbuf_4
XPHY_4016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20258__SET_B repeater217/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_227_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20925_ _20930_/CLK _20925_/D repeater268/X vssd1 vssd1 vccd1 vccd1 _20925_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_4049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_230_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20856_ _21459_/CLK _20856_/D repeater243/X vssd1 vssd1 vccd1 vccd1 _20856_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18392__S _18907_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10519__A _20690_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20787_ _21390_/CLK _20787_/D repeater240/X vssd1 vssd1 vccd1 vccd1 _20787_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10540_ _10540_/A _10540_/B _10723_/C vssd1 vssd1 vccd1 vccd1 _10701_/C sky130_fd_sc_hd__or3_1
XFILLER_10_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17930__C1 _17929_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10471_ _10452_/X _10471_/B _10471_/C _10471_/D vssd1 vssd1 vccd1 vccd1 _10523_/B
+ sky130_fd_sc_hd__and4b_1
XFILLER_10_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__21003__RESET_B repeater235/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18486__A0 _18485_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12210_ _20922_/Q vssd1 vssd1 vccd1 vccd1 _12470_/A sky130_fd_sc_hd__inv_2
XFILLER_108_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21408_ _21433_/CLK _21408_/D repeater236/X vssd1 vssd1 vccd1 vccd1 _21408_/Q sky130_fd_sc_hd__dfrtp_2
X_13190_ _13329_/A _13456_/B vssd1 vssd1 vccd1 vccd1 _13225_/A sky130_fd_sc_hd__or2_2
XFILLER_203_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12141_ _20393_/Q vssd1 vssd1 vccd1 vccd1 _18077_/A sky130_fd_sc_hd__inv_2
X_21339_ _21341_/CLK _21339_/D repeater222/X vssd1 vssd1 vccd1 vccd1 _21339_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_2_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12072_ _20965_/Q _12067_/Y _12332_/A _20393_/Q _12071_/X vssd1 vssd1 vccd1 vccd1
+ _12087_/B sky130_fd_sc_hd__o221a_1
XFILLER_89_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15900_ _19583_/Q _15896_/X _15793_/X _15897_/X vssd1 vssd1 vccd1 vccd1 _19583_/D
+ sky130_fd_sc_hd__a22o_1
X_11023_ _11596_/A _11022_/X _21243_/Q vssd1 vssd1 vccd1 vccd1 _21243_/D sky130_fd_sc_hd__mux2_1
XFILLER_77_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16880_ _10752_/B _16879_/X _16848_/X vssd1 vssd1 vccd1 vccd1 _16880_/X sky130_fd_sc_hd__o21a_1
XFILLER_131_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15831_ _16419_/A vssd1 vssd1 vccd1 vccd1 _16093_/A sky130_fd_sc_hd__buf_1
XFILLER_66_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18567__S _18907_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18550_ _18845_/A0 _10313_/Y _18884_/S vssd1 vssd1 vccd1 vccd1 _18550_/X sky130_fd_sc_hd__mux2_1
X_15762_ _15762_/A vssd1 vssd1 vccd1 vccd1 _15762_/X sky130_fd_sc_hd__buf_1
X_12974_ _17178_/A _12981_/A vssd1 vssd1 vccd1 vccd1 _12975_/S sky130_fd_sc_hd__or2_1
X_17501_ _11878_/Y _19583_/Q _17500_/X vssd1 vssd1 vccd1 vccd1 _17501_/Y sky130_fd_sc_hd__o21ai_1
X_14713_ _20155_/Q _14711_/X _12860_/A _14712_/X vssd1 vssd1 vccd1 vccd1 _20155_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_17_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11925_ _21006_/Q _11924_/X _21006_/Q _11924_/X vssd1 vssd1 vccd1 vccd1 _11926_/D
+ sky130_fd_sc_hd__a2bb2o_1
X_18481_ _18848_/A0 _14143_/Y _18884_/S vssd1 vssd1 vccd1 vccd1 _18481_/X sky130_fd_sc_hd__mux2_1
XANTENNA_output112_A _18109_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15693_ _19675_/Q _15688_/X _15663_/X _15690_/X vssd1 vssd1 vccd1 vccd1 _19675_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17432_ _19625_/Q vssd1 vssd1 vccd1 vccd1 _17432_/Y sky130_fd_sc_hd__inv_2
XPHY_4583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14644_ _14572_/A _14572_/B _14639_/X _14641_/Y vssd1 vssd1 vccd1 vccd1 _20182_/D
+ sky130_fd_sc_hd__a211oi_2
X_11856_ _21029_/Q _11856_/B vssd1 vssd1 vccd1 vccd1 _11856_/Y sky130_fd_sc_hd__nor2_1
XPHY_4594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10807_ _10807_/A vssd1 vssd1 vccd1 vccd1 _10807_/Y sky130_fd_sc_hd__inv_2
XFILLER_220_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14575_ _14575_/A _14575_/B _14637_/A vssd1 vssd1 vccd1 vccd1 _14633_/A sky130_fd_sc_hd__or3_1
X_17363_ _19440_/Q vssd1 vssd1 vccd1 vccd1 _17363_/Y sky130_fd_sc_hd__inv_2
X_11787_ _19874_/Q _16596_/D _16597_/A _16596_/C vssd1 vssd1 vccd1 vccd1 _11787_/X
+ sky130_fd_sc_hd__a211o_1
XPHY_3893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_repeater262_A repeater263/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19102_ _16668_/X _21076_/Q _19870_/D vssd1 vssd1 vccd1 vccd1 _19102_/X sky130_fd_sc_hd__mux2_1
XFILLER_159_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16314_ _16320_/A vssd1 vssd1 vccd1 vccd1 _16314_/X sky130_fd_sc_hd__buf_1
X_10738_ _19925_/Q _16773_/A vssd1 vssd1 vccd1 vccd1 _16777_/A sky130_fd_sc_hd__or2_4
X_13526_ _13526_/A vssd1 vssd1 vccd1 vccd1 _20432_/D sky130_fd_sc_hd__inv_2
XFILLER_186_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17294_ _21045_/Q vssd1 vssd1 vccd1 vccd1 _17294_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19033_ _16859_/X _20836_/Q _19046_/S vssd1 vssd1 vccd1 vccd1 _19943_/D sky130_fd_sc_hd__mux2_1
XFILLER_146_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16245_ _19414_/Q _16240_/X _16016_/X _16241_/X vssd1 vssd1 vccd1 vccd1 _19414_/D
+ sky130_fd_sc_hd__a22o_1
X_13457_ _13491_/A vssd1 vssd1 vccd1 vccd1 _13481_/A sky130_fd_sc_hd__clkbuf_2
X_10669_ _21337_/Q _21336_/Q _10669_/C vssd1 vssd1 vccd1 vccd1 _10669_/X sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_opt_0_HCLK_A clkbuf_opt_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12644__A _13046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12408_ _12408_/A _12490_/B _12408_/C vssd1 vssd1 vccd1 vccd1 _12409_/A sky130_fd_sc_hd__or3_4
X_16176_ _19448_/Q _16173_/X _16145_/X _16174_/X vssd1 vssd1 vccd1 vccd1 _19448_/D
+ sky130_fd_sc_hd__a22o_1
X_13388_ _17080_/A _13456_/B vssd1 vssd1 vccd1 vccd1 _13416_/A sky130_fd_sc_hd__or2_2
XFILLER_154_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput106 _17665_/Y vssd1 vssd1 vccd1 vccd1 HRDATA[5] sky130_fd_sc_hd__clkbuf_2
XFILLER_126_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput117 _18119_/LO vssd1 vssd1 vccd1 vccd1 IRQ[14] sky130_fd_sc_hd__clkbuf_2
XFILLER_115_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput128 _21120_/Q vssd1 vssd1 vccd1 vccd1 MSO_S2 sky130_fd_sc_hd__clkbuf_2
X_12339_ _12339_/A vssd1 vssd1 vccd1 vccd1 _12339_/Y sky130_fd_sc_hd__inv_2
X_15127_ _20443_/Q vssd1 vssd1 vccd1 vccd1 _15127_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15955__A _15961_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20797__RESET_B repeater255/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput139 _18122_/LO vssd1 vssd1 vccd1 vccd1 scl_o_S5 sky130_fd_sc_hd__clkbuf_2
XFILLER_217_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15058_ _20044_/Q vssd1 vssd1 vccd1 vccd1 _15059_/A sky130_fd_sc_hd__inv_2
X_19935_ _21242_/CLK _19935_/D repeater189/X vssd1 vssd1 vccd1 vccd1 _19935_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__20726__RESET_B repeater254/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14009_ _14009_/A vssd1 vssd1 vccd1 vccd1 _14031_/B sky130_fd_sc_hd__buf_1
XANTENNA__13475__A input52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19866_ _21182_/CLK input75/X repeater217/X vssd1 vssd1 vccd1 vccd1 _19867_/D sky130_fd_sc_hd__dfrtp_1
XANTENNA__20897__SET_B repeater212/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18817_ _17079_/Y _15237_/Y _18908_/S vssd1 vssd1 vccd1 vccd1 _18817_/X sky130_fd_sc_hd__mux2_1
X_19797_ _19811_/CLK _19797_/D vssd1 vssd1 vccd1 vccd1 _19797_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__18477__S _18904_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_244_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18748_ _18747_/X _20180_/Q _18748_/S vssd1 vssd1 vccd1 vccd1 _18748_/X sky130_fd_sc_hd__mux2_2
XFILLER_36_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18679_ _17281_/X _17710_/Y _18835_/S vssd1 vssd1 vccd1 vccd1 _18679_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12819__A _17083_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18952__A1 _21084_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20710_ _21357_/CLK _20710_/D repeater210/X vssd1 vssd1 vccd1 vccd1 _20710_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_24_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20641_ _20657_/CLK _20641_/D repeater198/X vssd1 vssd1 vccd1 vccd1 _20641_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_177_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19101__S _19870_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20572_ _20590_/CLK _20572_/D repeater258/X vssd1 vssd1 vccd1 vccd1 _20572_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18940__S _18946_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21124_ _21125_/CLK _21124_/D repeater190/X vssd1 vssd1 vccd1 vccd1 _21124_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_105_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13701__B1 _13506_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_127_HCLK_A clkbuf_4_4_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13385__A _13601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21055_ _21055_/CLK _21055_/D repeater220/X vssd1 vssd1 vccd1 vccd1 _21055_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_99_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18640__A0 _17079_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20006_ _21438_/CLK _20006_/D repeater240/X vssd1 vssd1 vccd1 vccd1 _20006_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_246_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09817_ _21452_/Q vssd1 vssd1 vccd1 vccd1 _15869_/A sky130_fd_sc_hd__buf_1
XANTENNA__18387__S _18908_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09748_ _21225_/Q _09746_/Y _21233_/Q _09747_/Y vssd1 vssd1 vccd1 vccd1 _09748_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_27_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09679_ _21469_/Q _09673_/X _09676_/X _09678_/X vssd1 vssd1 vccd1 vccd1 _21469_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_36_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11710_ _21071_/Q vssd1 vssd1 vccd1 vccd1 _16663_/A sky130_fd_sc_hd__clkbuf_2
XPHY_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20908_ _20908_/CLK _20908_/D repeater217/X vssd1 vssd1 vccd1 vccd1 _20908_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_36_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12690_ _20825_/Q _12686_/X _09645_/X _12688_/X vssd1 vssd1 vccd1 vccd1 _20825_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11641_ _11641_/A vssd1 vssd1 vccd1 vccd1 _11646_/A sky130_fd_sc_hd__inv_2
XPHY_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20839_ _20841_/CLK _20839_/D repeater256/X vssd1 vssd1 vccd1 vccd1 _20839_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19011__S _19019_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14360_ _20219_/Q vssd1 vssd1 vccd1 vccd1 _14504_/A sky130_fd_sc_hd__inv_2
XANTENNA__17320__A _17320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11572_ _21128_/Q _11562_/X _11571_/X _11566_/X vssd1 vssd1 vccd1 vccd1 _21128_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13311_ _13311_/A vssd1 vssd1 vccd1 vccd1 _13311_/X sky130_fd_sc_hd__buf_2
X_10523_ _10523_/A _10523_/B _10523_/C _10523_/D vssd1 vssd1 vccd1 vccd1 _10785_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_10_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput19 HADDR[26] vssd1 vssd1 vccd1 vccd1 input19/X sky130_fd_sc_hd__buf_1
XPHY_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14291_ _14779_/B _14288_/X _15335_/B _20121_/Q _14290_/Y vssd1 vssd1 vccd1 vccd1
+ _14302_/B sky130_fd_sc_hd__a221o_1
XPHY_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18850__S _18850_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13242_ _20572_/Q _13239_/X _13240_/X _13241_/X vssd1 vssd1 vccd1 vccd1 _20572_/D
+ sky130_fd_sc_hd__a22o_1
X_16030_ _19521_/Q _16028_/X _15769_/X _16029_/X vssd1 vssd1 vccd1 vccd1 _19521_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_input73_A RsRx_S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10454_ _20696_/Q vssd1 vssd1 vccd1 vccd1 _10454_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_142_HCLK clkbuf_4_3_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _21239_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__19120__A1 _14275_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20890__RESET_B repeater185/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13173_ _13714_/A vssd1 vssd1 vccd1 vccd1 _13173_/X sky130_fd_sc_hd__clkbuf_4
X_10385_ _10385_/A vssd1 vssd1 vccd1 vccd1 _10385_/Y sky130_fd_sc_hd__inv_2
X_12124_ _12119_/X _20388_/Q _12329_/A _20390_/Q _12123_/X vssd1 vssd1 vccd1 vccd1
+ _12144_/A sky130_fd_sc_hd__o221a_1
XANTENNA__19735__CLK _19765_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17981_ _17981_/A _18001_/B vssd1 vssd1 vccd1 vccd1 _17981_/Y sky130_fd_sc_hd__nor2_1
X_19720_ _20326_/CLK _19720_/D vssd1 vssd1 vccd1 vccd1 _19720_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20137__RESET_B repeater248/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16932_ _16930_/Y _16931_/Y _16915_/X vssd1 vssd1 vccd1 vccd1 _16932_/X sky130_fd_sc_hd__o21a_1
X_12055_ _20364_/Q vssd1 vssd1 vccd1 vccd1 _12055_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18631__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11006_ _21013_/Q vssd1 vssd1 vccd1 vccd1 _15505_/A sky130_fd_sc_hd__buf_1
X_19651_ _19821_/CLK _19651_/D vssd1 vssd1 vccd1 vccd1 _19651_/Q sky130_fd_sc_hd__dfxtp_1
X_16863_ _16863_/A _16863_/B vssd1 vssd1 vccd1 vccd1 _16863_/Y sky130_fd_sc_hd__nor2_1
XFILLER_238_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18297__S _18644_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14248__B2 _18946_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_49_HCLK_A clkbuf_4_9_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18602_ _18601_/X _14103_/X _18904_/S vssd1 vssd1 vccd1 vccd1 _18602_/X sky130_fd_sc_hd__mux2_1
XFILLER_203_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15814_ _20136_/Q vssd1 vssd1 vccd1 vccd1 _16165_/B sky130_fd_sc_hd__buf_1
X_19582_ _19821_/CLK _19582_/D vssd1 vssd1 vccd1 vccd1 _19582_/Q sky130_fd_sc_hd__dfxtp_1
X_16794_ _16794_/A vssd1 vssd1 vccd1 vccd1 _16794_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18533_ _17940_/Y _20651_/Q _18903_/S vssd1 vssd1 vccd1 vccd1 _18533_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15745_ _15751_/A vssd1 vssd1 vccd1 vccd1 _15745_/X sky130_fd_sc_hd__buf_1
XFILLER_234_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12957_ _14264_/A vssd1 vssd1 vccd1 vccd1 _12957_/X sky130_fd_sc_hd__buf_2
XFILLER_61_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19282__S1 _21017_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17737__A2 _17719_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18934__A1 _21142_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11908_ _21014_/Q vssd1 vssd1 vccd1 vccd1 _15559_/A sky130_fd_sc_hd__inv_2
X_18464_ _17900_/Y _20752_/Q _18775_/S vssd1 vssd1 vccd1 vccd1 _18464_/X sky130_fd_sc_hd__mux2_1
X_15676_ _15682_/A vssd1 vssd1 vccd1 vccd1 _15676_/X sky130_fd_sc_hd__buf_1
XPHY_4380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12888_ _17178_/A _12899_/A vssd1 vssd1 vccd1 vccd1 _12889_/S sky130_fd_sc_hd__or2_1
XPHY_4391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17415_ _19521_/Q vssd1 vssd1 vccd1 vccd1 _17415_/Y sky130_fd_sc_hd__inv_2
XFILLER_221_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14627_ _14627_/A vssd1 vssd1 vccd1 vccd1 _14627_/Y sky130_fd_sc_hd__inv_2
X_11839_ _11833_/B _11827_/X _11838_/Y _11834_/X _11811_/A vssd1 vssd1 vccd1 vccd1
+ _11840_/A sky130_fd_sc_hd__o32a_1
X_18395_ _18394_/X _14077_/A _18850_/S vssd1 vssd1 vccd1 vccd1 _18395_/X sky130_fd_sc_hd__mux2_1
XPHY_3690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18698__A0 _17079_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17346_ _21215_/Q vssd1 vssd1 vccd1 vccd1 _17346_/Y sky130_fd_sc_hd__inv_2
X_14558_ _16405_/B vssd1 vssd1 vccd1 vccd1 _15833_/B sky130_fd_sc_hd__buf_1
X_13509_ _14262_/A vssd1 vssd1 vccd1 vccd1 _13509_/X sky130_fd_sc_hd__buf_2
XFILLER_146_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17277_ _19310_/Q _17533_/B vssd1 vssd1 vccd1 vccd1 _17277_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__18760__S _18929_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14489_ _14461_/D _14368_/B _14486_/Y _14488_/X vssd1 vssd1 vccd1 vccd1 _20225_/D
+ sky130_fd_sc_hd__a211oi_2
X_19016_ _16928_/X _20407_/Q _19019_/S vssd1 vssd1 vccd1 vccd1 _19960_/D sky130_fd_sc_hd__mux2_1
X_16228_ _19422_/Q _16223_/X _16127_/X _16224_/X vssd1 vssd1 vccd1 vccd1 _19422_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__20907__RESET_B repeater217/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19111__A1 _20251_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20242__CLK _21452_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16159_ _16159_/A vssd1 vssd1 vccd1 vccd1 _16159_/X sky130_fd_sc_hd__buf_1
XFILLER_170_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15684__B1 _15588_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19918_ _21406_/CLK _19918_/D repeater213/X vssd1 vssd1 vccd1 vccd1 _19918_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_244_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_228_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19849_ _21183_/CLK _19849_/D repeater219/X vssd1 vssd1 vccd1 vccd1 _19851_/D sky130_fd_sc_hd__dfstp_1
XFILLER_84_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_228_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09602_ _20891_/Q _19986_/Q vssd1 vssd1 vccd1 vccd1 _10975_/A sky130_fd_sc_hd__nand2_1
XFILLER_243_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_23_HCLK clkbuf_4_9_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _21390_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_25_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18935__S _18946_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19273__S1 _21004_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18925__A1 _19271_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_224_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18689__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20624_ _20697_/CLK _20624_/D repeater193/X vssd1 vssd1 vccd1 vccd1 _20624_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_165_HCLK clkbuf_opt_0_HCLK/A vssd1 vssd1 vccd1 vccd1 _21445_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_149_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20555_ _20592_/CLK _20555_/D repeater260/X vssd1 vssd1 vccd1 vccd1 _20555_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__18670__S _18748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19758__CLK _21009_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20486_ _20937_/CLK _20486_/D repeater277/X vssd1 vssd1 vccd1 vccd1 _20486_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_192_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10170_ _10183_/A vssd1 vssd1 vccd1 vccd1 _10170_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_160_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_248_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20230__RESET_B repeater203/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21107_ _21424_/CLK _21107_/D repeater231/X vssd1 vssd1 vccd1 vccd1 _21107_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_154_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18613__A0 _18848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21038_ _21401_/CLK _21038_/D repeater242/X vssd1 vssd1 vccd1 vccd1 _21038_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_208_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19006__S _19019_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13860_ _20563_/Q vssd1 vssd1 vccd1 vccd1 _14030_/A sky130_fd_sc_hd__inv_2
XFILLER_170_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12811_ _12809_/X _20772_/Q _12811_/S vssd1 vssd1 vccd1 vccd1 _20772_/D sky130_fd_sc_hd__mux2_1
XFILLER_34_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13791_ _13789_/Y _20191_/Q _20614_/Q _14580_/A vssd1 vssd1 vccd1 vccd1 _13791_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__18845__S _18896_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19264__S1 _21004_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_231_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15530_ _15536_/A vssd1 vssd1 vccd1 vccd1 _15537_/A sky130_fd_sc_hd__inv_2
XFILLER_188_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12742_ _12742_/A vssd1 vssd1 vccd1 vccd1 _12743_/B sky130_fd_sc_hd__inv_2
XANTENNA__12661__B1 _12660_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_242_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15461_ _19785_/Q _15459_/X _15424_/X _15460_/X vssd1 vssd1 vccd1 vccd1 _19785_/D
+ sky130_fd_sc_hd__a22o_1
X_12673_ input53/X vssd1 vssd1 vccd1 vccd1 _12673_/X sky130_fd_sc_hd__buf_4
XFILLER_63_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17200_ _17933_/A vssd1 vssd1 vccd1 vccd1 _17200_/X sky130_fd_sc_hd__clkbuf_2
XPHY_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14412_ _14395_/Y _20225_/Q _14411_/Y _20230_/Q vssd1 vssd1 vccd1 vccd1 _14412_/X
+ sky130_fd_sc_hd__o22a_1
X_11624_ _21104_/Q vssd1 vssd1 vccd1 vccd1 _14813_/C sky130_fd_sc_hd__buf_1
XPHY_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18180_ _18179_/X _13917_/Y _18903_/S vssd1 vssd1 vccd1 vccd1 _18180_/X sky130_fd_sc_hd__mux2_1
XPHY_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15392_ _19816_/Q _15389_/X _15350_/X _15390_/X vssd1 vssd1 vccd1 vccd1 _19816_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17131_ _19333_/Q vssd1 vssd1 vccd1 vccd1 _17131_/Y sky130_fd_sc_hd__inv_2
XPHY_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14343_ _14343_/A vssd1 vssd1 vccd1 vccd1 _14462_/B sky130_fd_sc_hd__clkbuf_2
X_11555_ _21134_/Q _11552_/X _10884_/X _11554_/X vssd1 vssd1 vccd1 vccd1 _21134_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_168_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18580__S _18669_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10506_ _20667_/Q vssd1 vssd1 vccd1 vccd1 _10506_/Y sky130_fd_sc_hd__inv_2
X_17062_ _19877_/Q vssd1 vssd1 vccd1 vccd1 _17062_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20389__RESET_B repeater278/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14274_ _13600_/X _20243_/Q _14274_/S vssd1 vssd1 vccd1 vccd1 _20243_/D sky130_fd_sc_hd__mux2_1
XFILLER_10_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11486_ _15377_/A vssd1 vssd1 vccd1 vccd1 _11486_/X sky130_fd_sc_hd__buf_4
XFILLER_171_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16013_ _19528_/Q _16008_/X _16012_/X _16010_/X vssd1 vssd1 vccd1 vccd1 _19528_/D
+ sky130_fd_sc_hd__a22o_1
X_13225_ _13225_/A vssd1 vssd1 vccd1 vccd1 _13248_/A sky130_fd_sc_hd__buf_1
XFILLER_137_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10437_ _21301_/Q vssd1 vssd1 vccd1 vccd1 _10777_/A sky130_fd_sc_hd__inv_2
XANTENNA__20318__RESET_B repeater262/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater225_A repeater226/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12922__A input50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13156_ _20608_/Q _13150_/X _13030_/X _13152_/X vssd1 vssd1 vccd1 vccd1 _20608_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_88_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10368_ _10289_/A _10289_/B _10290_/Y _10405_/B vssd1 vssd1 vccd1 vccd1 _21374_/D
+ sky130_fd_sc_hd__a211oi_4
X_12107_ _20370_/Q vssd1 vssd1 vccd1 vccd1 _12107_/Y sky130_fd_sc_hd__inv_2
X_17964_ _18194_/X _17963_/X _18199_/X _17947_/A vssd1 vssd1 vccd1 vccd1 _17964_/X
+ sky130_fd_sc_hd__o22a_1
X_13087_ _13099_/A vssd1 vssd1 vccd1 vccd1 _13087_/X sky130_fd_sc_hd__buf_1
X_10299_ _20717_/Q vssd1 vssd1 vccd1 vccd1 _17901_/A sky130_fd_sc_hd__inv_2
XFILLER_214_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18604__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19703_ _19828_/CLK _19703_/D vssd1 vssd1 vccd1 vccd1 _19703_/Q sky130_fd_sc_hd__dfxtp_1
X_16915_ _16915_/A vssd1 vssd1 vccd1 vccd1 _16915_/X sky130_fd_sc_hd__buf_1
X_12038_ _20391_/Q vssd1 vssd1 vccd1 vccd1 _12038_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_46_HCLK _20004_/CLK vssd1 vssd1 vccd1 vccd1 _21151_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_clkbuf_leaf_110_HCLK_A clkbuf_opt_3_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17895_ _17895_/A _17898_/B vssd1 vssd1 vccd1 vccd1 _17895_/Y sky130_fd_sc_hd__nor2_1
XFILLER_77_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17225__A _17320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19634_ _20142_/CLK _19634_/D vssd1 vssd1 vccd1 vccd1 _19634_/Q sky130_fd_sc_hd__dfxtp_1
X_16846_ _16844_/Y _16845_/X _16831_/X vssd1 vssd1 vccd1 vccd1 _16846_/X sky130_fd_sc_hd__o21a_1
XFILLER_225_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__21177__RESET_B repeater216/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19565_ _19706_/CLK _19565_/D vssd1 vssd1 vccd1 vccd1 _19565_/Q sky130_fd_sc_hd__dfxtp_1
X_16777_ _16777_/A vssd1 vssd1 vccd1 vccd1 _16777_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19255__S1 _21004_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13989_ _20314_/Q _13986_/Y _13891_/B _13988_/X vssd1 vssd1 vccd1 vccd1 _20314_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_241_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18516_ _17942_/Y _20755_/Q _18775_/S vssd1 vssd1 vccd1 vccd1 _18516_/X sky130_fd_sc_hd__mux2_1
X_15728_ _19661_/Q _15723_/X _15725_/X _15727_/X vssd1 vssd1 vccd1 vccd1 _19661_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_179_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19496_ _20326_/CLK _19496_/D vssd1 vssd1 vccd1 vccd1 _19496_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_234_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18447_ _18446_/X _10635_/Y _18885_/S vssd1 vssd1 vccd1 vccd1 _18447_/X sky130_fd_sc_hd__mux2_1
XFILLER_221_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15659_ _15667_/A vssd1 vssd1 vccd1 vccd1 _15659_/X sky130_fd_sc_hd__buf_1
XFILLER_33_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09678__A _15330_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18378_ _18377_/X _16778_/A _18880_/S vssd1 vssd1 vccd1 vccd1 _18378_/X sky130_fd_sc_hd__mux2_1
XFILLER_221_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17895__A _17895_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17329_ _17158_/X _17298_/X _17170_/X _17309_/X _17328_/X vssd1 vssd1 vccd1 vccd1
+ _17329_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_146_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18490__S _18908_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14157__B1 _20550_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20741__RESET_B repeater207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20340_ _20949_/CLK _20340_/D repeater269/X vssd1 vssd1 vccd1 vccd1 _20340_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_107_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20059__RESET_B repeater281/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20271_ _20724_/CLK _20271_/D repeater263/X vssd1 vssd1 vccd1 vccd1 _20271_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_108_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19191__S0 _20123_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15409__B1 _15352_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_229_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11694__A1 _21080_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_32_HCLK_A clkbuf_opt_4_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18665__S _18884_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19246__S1 _21006_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19995__RESET_B repeater218/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_95_HCLK_A clkbuf_4_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11183__A _15884_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_213_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19924__RESET_B repeater212/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20829__RESET_B repeater251/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12726__B _17153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20607_ _20622_/CLK _20607_/D repeater195/X vssd1 vssd1 vccd1 vccd1 _20607_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_193_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11340_ _11340_/A vssd1 vssd1 vccd1 vccd1 _11341_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_165_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20538_ _20592_/CLK _20538_/D repeater267/X vssd1 vssd1 vccd1 vccd1 _20538_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_193_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11271_ _12506_/A _20912_/Q _11271_/C _11286_/C vssd1 vssd1 vccd1 vccd1 _11272_/B
+ sky130_fd_sc_hd__or4b_4
XFILLER_192_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20411__RESET_B repeater185/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20469_ _20470_/CLK _20469_/D repeater279/X vssd1 vssd1 vccd1 vccd1 _20469_/Q sky130_fd_sc_hd__dfrtp_1
X_13010_ _20687_/Q _13005_/X _12920_/X _13007_/X vssd1 vssd1 vccd1 vccd1 _20687_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19182__S0 _19280_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10222_ _10041_/B _10224_/A _10041_/A vssd1 vssd1 vccd1 vccd1 _10223_/B sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_69_HCLK clkbuf_opt_7_HCLK/A vssd1 vssd1 vccd1 vccd1 _20220_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_79_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10153_ _10153_/A _10153_/B vssd1 vssd1 vccd1 vccd1 _10190_/A sky130_fd_sc_hd__or2_1
XFILLER_160_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input36_A HTRANS[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14961_ _14961_/A _14961_/B _14961_/C _14961_/D vssd1 vssd1 vccd1 vccd1 _14962_/D
+ sky130_fd_sc_hd__or4_4
X_10084_ _21403_/Q _10080_/Y _21382_/Q _10081_/Y _10083_/X vssd1 vssd1 vccd1 vccd1
+ _10098_/A sky130_fd_sc_hd__o221a_1
Xhold8 hold8/A vssd1 vssd1 vccd1 vccd1 hold8/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_248_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16700_ _16700_/A _18942_/X vssd1 vssd1 vccd1 vccd1 _19894_/D sky130_fd_sc_hd__and2_1
XANTENNA__13573__A _13594_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13912_ _20650_/Q _13883_/A _13911_/Y _20307_/Q vssd1 vssd1 vccd1 vccd1 _13912_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11685__A1 _21086_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10488__A2 _20691_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17680_ _19298_/Q vssd1 vssd1 vccd1 vccd1 _17680_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12882__B1 _12881_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14892_ _14891_/Y _14883_/A _20595_/Q _20106_/Q vssd1 vssd1 vccd1 vccd1 _14892_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_235_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16631_ _16631_/A _17162_/A vssd1 vssd1 vccd1 vccd1 _19876_/D sky130_fd_sc_hd__nor2_1
XFILLER_74_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13843_ _20318_/Q vssd1 vssd1 vccd1 vccd1 _13894_/B sky130_fd_sc_hd__inv_2
XANTENNA__18575__S _18903_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19237__S1 _20131_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19350_ _20137_/CLK _19350_/D vssd1 vssd1 vccd1 vccd1 _19350_/Q sky130_fd_sc_hd__dfxtp_1
X_16562_ _16548_/A _19913_/Q _16553_/A _16556_/A _16556_/B vssd1 vssd1 vccd1 vccd1
+ _16562_/X sky130_fd_sc_hd__o32a_1
XFILLER_16_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13774_ _20176_/Q vssd1 vssd1 vccd1 vccd1 _14566_/A sky130_fd_sc_hd__inv_2
X_10986_ _21015_/Q vssd1 vssd1 vccd1 vccd1 _15653_/A sky130_fd_sc_hd__inv_2
XFILLER_216_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18301_ _18848_/A0 _17967_/Y _18666_/S vssd1 vssd1 vccd1 vccd1 _18301_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15513_ input64/X vssd1 vssd1 vccd1 vccd1 _15785_/A sky130_fd_sc_hd__buf_1
X_19281_ _19277_/X _19278_/X _19279_/X _19280_/X _20123_/Q _20124_/Q vssd1 vssd1 vccd1
+ vccd1 _19281_/X sky130_fd_sc_hd__mux4_2
X_12725_ _17060_/A _12725_/B _17140_/B _13383_/A vssd1 vssd1 vccd1 vccd1 _17153_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_231_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16493_ _19843_/Q vssd1 vssd1 vccd1 vccd1 _16681_/B sky130_fd_sc_hd__buf_1
XFILLER_70_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_repeater175_A _18644_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18232_ _20856_/Q input5/X _18236_/S vssd1 vssd1 vccd1 vccd1 _18232_/X sky130_fd_sc_hd__mux2_1
XFILLER_231_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15444_ _19792_/Q _15441_/X _15427_/X _15442_/X vssd1 vssd1 vccd1 vccd1 _19792_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_31_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12656_ input61/X vssd1 vssd1 vccd1 vccd1 _12656_/X sky130_fd_sc_hd__clkbuf_4
XPHY_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18163_ _18848_/A0 _14102_/Y _18902_/S vssd1 vssd1 vccd1 vccd1 _18163_/X sky130_fd_sc_hd__mux2_1
X_11607_ _18991_/X _11598_/A _21115_/Q _11605_/X vssd1 vssd1 vccd1 vccd1 _21115_/D
+ sky130_fd_sc_hd__a22o_1
X_12587_ _20881_/Q _12581_/X _18233_/X _12583_/X vssd1 vssd1 vccd1 vccd1 _20881_/D
+ sky130_fd_sc_hd__a22o_1
X_15375_ _15375_/A _15542_/B _15708_/C vssd1 vssd1 vccd1 vccd1 _15389_/A sky130_fd_sc_hd__or3_4
XFILLER_156_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17114_ _19478_/Q vssd1 vssd1 vccd1 vccd1 _17114_/Y sky130_fd_sc_hd__inv_2
XPHY_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14326_ _20239_/Q vssd1 vssd1 vccd1 vccd1 _14382_/A sky130_fd_sc_hd__inv_2
X_11538_ _21137_/Q _11534_/X _10898_/X _11535_/X vssd1 vssd1 vccd1 vccd1 _21137_/D
+ sky130_fd_sc_hd__a22o_1
X_18094_ _18642_/X _17858_/X _18639_/X _17211_/X _18093_/X vssd1 vssd1 vccd1 vccd1
+ _18097_/B sky130_fd_sc_hd__o221a_2
XFILLER_156_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17045_ _21095_/Q _17044_/Y _16684_/A vssd1 vssd1 vccd1 vccd1 _19839_/D sky130_fd_sc_hd__o21ai_1
X_11469_ _11481_/A vssd1 vssd1 vccd1 vccd1 _11469_/X sky130_fd_sc_hd__buf_1
X_14257_ _14267_/A vssd1 vssd1 vccd1 vccd1 _14257_/X sky130_fd_sc_hd__buf_1
XANTENNA__19173__S0 _19280_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13208_ _20588_/Q _13206_/X _13006_/X _13207_/X vssd1 vssd1 vccd1 vccd1 _20588_/D
+ sky130_fd_sc_hd__a22o_1
X_14188_ _20284_/Q _14187_/Y _14183_/X _14095_/B vssd1 vssd1 vccd1 vccd1 _20284_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_140_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13139_ _13165_/A vssd1 vssd1 vccd1 vccd1 _13139_/X sky130_fd_sc_hd__buf_1
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18996_ _17013_/Y _20427_/Q _19026_/S vssd1 vssd1 vccd1 vccd1 _19980_/D sky130_fd_sc_hd__mux2_1
XFILLER_100_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21358__RESET_B repeater254/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater203 repeater204/X vssd1 vssd1 vccd1 vccd1 repeater203/X sky130_fd_sc_hd__clkbuf_8
X_17947_ _17947_/A vssd1 vssd1 vccd1 vccd1 _17947_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_97_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrepeater214 repeater215/X vssd1 vssd1 vccd1 vccd1 repeater214/X sky130_fd_sc_hd__buf_6
Xrepeater225 repeater226/X vssd1 vssd1 vccd1 vccd1 repeater225/X sky130_fd_sc_hd__clkbuf_8
XFILLER_227_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13483__A _13483_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater236 repeater237/X vssd1 vssd1 vccd1 vccd1 repeater236/X sky130_fd_sc_hd__buf_6
XANTENNA__11676__A1 _21088_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater247 repeater248/X vssd1 vssd1 vccd1 vccd1 repeater247/X sky130_fd_sc_hd__buf_8
XANTENNA__12873__B1 _12872_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17878_ _18543_/X _17853_/X _18556_/X _17854_/X vssd1 vssd1 vccd1 vccd1 _17878_/X
+ sky130_fd_sc_hd__o22a_1
Xrepeater258 repeater266/X vssd1 vssd1 vccd1 vccd1 repeater258/X sky130_fd_sc_hd__buf_4
XFILLER_226_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater269 repeater270/X vssd1 vssd1 vccd1 vccd1 repeater269/X sky130_fd_sc_hd__clkbuf_8
XFILLER_65_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19617_ _21449_/CLK _19617_/D vssd1 vssd1 vccd1 vccd1 _19617_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16829_ _16829_/A vssd1 vssd1 vccd1 vccd1 _16829_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17800__B2 _18048_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19228__S1 _20131_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18485__S _18784_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19548_ _21459_/CLK _19548_/D vssd1 vssd1 vccd1 vccd1 _19548_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_207_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19479_ _19961_/CLK _19479_/D vssd1 vssd1 vccd1 vccd1 _19479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21441_ _21445_/CLK _21441_/D repeater244/X vssd1 vssd1 vccd1 vccd1 _21441_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_159_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21372_ _21372_/CLK _21372_/D repeater257/X vssd1 vssd1 vccd1 vccd1 _21372_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_134_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20323_ _21480_/CLK _20323_/D repeater206/X vssd1 vssd1 vccd1 vccd1 _20323_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_79_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19164__S0 _19280_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20254_ _20908_/CLK _20254_/D repeater217/X vssd1 vssd1 vccd1 vccd1 _20254_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_116_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20185_ _20623_/CLK _20185_/D repeater194/X vssd1 vssd1 vccd1 vccd1 _20185_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_135_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09996_ _21419_/Q vssd1 vssd1 vccd1 vccd1 _09996_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12864__B1 _12863_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19219__S1 _20131_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18395__S _18850_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10840_ _21278_/Q _10839_/Y _10830_/X _10756_/B vssd1 vssd1 vccd1 vccd1 _21278_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_232_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20923__CLK _20930_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10771_ _10771_/A _10771_/B vssd1 vssd1 vccd1 vccd1 _10807_/A sky130_fd_sc_hd__or2_1
XFILLER_44_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12510_ _12510_/A vssd1 vssd1 vccd1 vccd1 _20917_/D sky130_fd_sc_hd__inv_2
XFILLER_44_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13490_ _20449_/Q _13481_/X _13489_/X _13483_/X vssd1 vssd1 vccd1 vccd1 _20449_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_40_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12441_ _20945_/Q _12440_/Y _12395_/B _12440_/A _12411_/X vssd1 vssd1 vccd1 vccd1
+ _20945_/D sky130_fd_sc_hd__o221a_1
XFILLER_40_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15160_ _15177_/A vssd1 vssd1 vccd1 vccd1 _15160_/X sky130_fd_sc_hd__clkbuf_2
X_12372_ _12372_/A vssd1 vssd1 vccd1 vccd1 _12376_/B sky130_fd_sc_hd__inv_2
XFILLER_138_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11323_ _21185_/Q _11322_/B _16564_/A _11322_/Y vssd1 vssd1 vccd1 vccd1 _21185_/D
+ sky130_fd_sc_hd__a211o_1
X_14111_ _20548_/Q _14087_/A _14108_/Y _20282_/Q _14110_/X vssd1 vssd1 vccd1 vccd1
+ _14120_/B sky130_fd_sc_hd__o221a_1
XFILLER_153_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15091_ _20442_/Q vssd1 vssd1 vccd1 vccd1 _15091_/Y sky130_fd_sc_hd__inv_2
XFILLER_181_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19155__S0 _19285_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11254_ _19065_/X _11250_/X _21187_/Q _11251_/X vssd1 vssd1 vccd1 vccd1 _21187_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_141_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14042_ _20286_/Q vssd1 vssd1 vccd1 vccd1 _14096_/A sky130_fd_sc_hd__inv_2
XANTENNA__17982__B _18001_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10205_ _10205_/A _10205_/B vssd1 vssd1 vccd1 vccd1 _10210_/A sky130_fd_sc_hd__or2_1
XFILLER_192_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18850_ _18849_/X _14071_/A _18850_/S vssd1 vssd1 vccd1 vccd1 _18850_/X sky130_fd_sc_hd__mux2_1
X_11185_ _15885_/A _17684_/A vssd1 vssd1 vccd1 vccd1 _11186_/S sky130_fd_sc_hd__or2_1
XANTENNA__21451__RESET_B repeater247/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17801_ _18138_/X _17581_/A _18673_/X _17226_/A vssd1 vssd1 vccd1 vccd1 _17801_/X
+ sky130_fd_sc_hd__o22a_1
X_10136_ _10125_/X _10136_/B _10136_/C _10136_/D vssd1 vssd1 vccd1 vccd1 _10137_/D
+ sky130_fd_sc_hd__and4b_1
X_18781_ _18780_/X _13943_/Y _18849_/S vssd1 vssd1 vccd1 vccd1 _18781_/X sky130_fd_sc_hd__mux2_1
X_15993_ _15993_/A vssd1 vssd1 vccd1 vccd1 _15993_/X sky130_fd_sc_hd__buf_1
XFILLER_95_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17732_ _17732_/A vssd1 vssd1 vccd1 vccd1 _17869_/A sky130_fd_sc_hd__buf_1
X_14944_ _20567_/Q _14853_/B _20594_/Q _14882_/A _14943_/X vssd1 vssd1 vccd1 vccd1
+ _14948_/C sky130_fd_sc_hd__o221a_1
X_10067_ _10155_/A _10154_/A _10156_/A _10153_/A vssd1 vssd1 vccd1 vccd1 _10068_/D
+ sky130_fd_sc_hd__or4_4
XFILLER_248_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16046__B1 _16014_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17663_ _18712_/X _17856_/A _18721_/X _17480_/X vssd1 vssd1 vccd1 vccd1 _17663_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_208_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14875_ _14960_/A _14981_/A vssd1 vssd1 vccd1 vccd1 _14876_/B sky130_fd_sc_hd__or2_2
XFILLER_75_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19402_ _21009_/CLK _19402_/D vssd1 vssd1 vccd1 vccd1 _19402_/Q sky130_fd_sc_hd__dfxtp_1
X_16614_ _16613_/Y _16605_/X _16539_/X _16541_/X vssd1 vssd1 vccd1 vccd1 _16614_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_211_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13826_ _20184_/Q vssd1 vssd1 vccd1 vccd1 _14574_/A sky130_fd_sc_hd__inv_2
XANTENNA__12607__B1 _18221_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17594_ _19395_/Q vssd1 vssd1 vccd1 vccd1 _17594_/Y sky130_fd_sc_hd__inv_2
XFILLER_235_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19333_ _20172_/CLK _19333_/D vssd1 vssd1 vccd1 vccd1 _19333_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_232_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16545_ _16545_/A vssd1 vssd1 vccd1 vccd1 _16689_/B sky130_fd_sc_hd__buf_1
X_13757_ _20628_/Q vssd1 vssd1 vccd1 vccd1 _18081_/A sky130_fd_sc_hd__inv_2
X_10969_ _10969_/A _10969_/B _10969_/C _10969_/D vssd1 vssd1 vccd1 vccd1 _10970_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_203_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12708_ _12708_/A vssd1 vssd1 vccd1 vccd1 _12708_/X sky130_fd_sc_hd__buf_1
XFILLER_31_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19264_ _17244_/Y _17245_/Y _17246_/Y _17247_/Y _19275_/S0 _21004_/Q vssd1 vssd1
+ vccd1 vccd1 _19264_/X sky130_fd_sc_hd__mux4_2
X_16476_ _19294_/Q _16473_/X _16291_/X _16474_/X vssd1 vssd1 vccd1 vccd1 _19294_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_203_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13688_ _13708_/A vssd1 vssd1 vccd1 vccd1 _13688_/X sky130_fd_sc_hd__buf_1
X_18215_ _18214_/X _17990_/Y _18903_/S vssd1 vssd1 vccd1 vccd1 _18215_/X sky130_fd_sc_hd__mux2_1
XFILLER_176_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20333__RESET_B repeater270/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15427_ _15588_/A vssd1 vssd1 vccd1 vccd1 _15427_/X sky130_fd_sc_hd__clkbuf_2
X_12639_ input27/X _12637_/X _20847_/Q _12638_/X vssd1 vssd1 vccd1 vccd1 _20847_/D
+ sky130_fd_sc_hd__o22a_1
XPHY_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19195_ _19306_/Q _19828_/Q _19836_/Q _19420_/Q _19280_/S0 _20122_/Q vssd1 vssd1
+ vccd1 vccd1 _19195_/X sky130_fd_sc_hd__mux4_2
XFILLER_145_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18146_ _18145_/X _10090_/Y _18644_/S vssd1 vssd1 vccd1 vccd1 _18146_/X sky130_fd_sc_hd__mux2_1
X_15358_ _15448_/A _15967_/B _16325_/C vssd1 vssd1 vccd1 vccd1 _15366_/A sky130_fd_sc_hd__or3_4
X_14309_ _14309_/A _14309_/B vssd1 vssd1 vccd1 vccd1 _16481_/B sky130_fd_sc_hd__nand2_2
XFILLER_171_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18077_ _18077_/A _18078_/B vssd1 vssd1 vccd1 vccd1 _18077_/Y sky130_fd_sc_hd__nor2_1
X_15289_ _19855_/Q _15289_/B vssd1 vssd1 vccd1 vccd1 _15290_/B sky130_fd_sc_hd__or2_1
XFILLER_171_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17028_ _21248_/Q vssd1 vssd1 vccd1 vccd1 _17028_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09850_ _20033_/Q vssd1 vssd1 vccd1 vccd1 _10843_/B sky130_fd_sc_hd__buf_1
XFILLER_86_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09691__A input60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17482__C1 _17479_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09781_ _16620_/A _09781_/B vssd1 vssd1 vccd1 vccd1 _09781_/Y sky130_fd_sc_hd__nor2_1
X_18979_ _21427_/Q _21100_/Q _18983_/S vssd1 vssd1 vccd1 vccd1 _18979_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12846__B1 _09638_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10630__A _20767_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_227_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20941_ _20950_/CLK _20941_/D repeater272/X vssd1 vssd1 vccd1 vccd1 _20941_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_227_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19104__S _19870_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_214_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20872_ _21452_/CLK _20872_/D repeater247/X vssd1 vssd1 vccd1 vccd1 _20872_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_42_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18943__S _18946_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13271__B1 _13270_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_210_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19985__D _19985_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20074__RESET_B repeater276/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13023__B1 _12853_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21424_ _21424_/CLK _21424_/D repeater231/X vssd1 vssd1 vccd1 vccd1 _21424_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_148_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13388__A _17080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21355_ _21407_/CLK _21355_/D repeater252/X vssd1 vssd1 vccd1 vccd1 _21355_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__19137__S0 _19285_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20306_ _20693_/CLK _20306_/D repeater196/X vssd1 vssd1 vccd1 vccd1 _20306_/Q sky130_fd_sc_hd__dfrtp_4
X_21286_ _21306_/CLK _21286_/D repeater207/X vssd1 vssd1 vccd1 vccd1 _21286_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_190_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21209__RESET_B repeater242/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20237_ _21477_/CLK _20237_/D repeater204/X vssd1 vssd1 vccd1 vccd1 _20237_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_150_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20168_ _21125_/CLK _20168_/D repeater190/X vssd1 vssd1 vccd1 vccd1 _20168_/Q sky130_fd_sc_hd__dfrtp_1
X_09979_ _21415_/Q _09975_/X _09688_/X _09976_/X vssd1 vssd1 vccd1 vccd1 _21415_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12837__B1 _12673_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12990_ _20696_/Q _12983_/X _12989_/X _12987_/X vssd1 vssd1 vccd1 vccd1 _20696_/D
+ sky130_fd_sc_hd__a22o_1
X_20099_ _20101_/CLK _20099_/D repeater259/X vssd1 vssd1 vccd1 vccd1 _20099_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_183_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11941_ _11165_/X _11940_/B _19116_/S _11940_/Y _11917_/X vssd1 vssd1 vccd1 vccd1
+ _11941_/X sky130_fd_sc_hd__o221a_1
XANTENNA__16579__A1 _16495_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_217_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19014__S _19019_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_232_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20844__RESET_B repeater243/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14660_ _14660_/A vssd1 vssd1 vccd1 vccd1 _14660_/Y sky130_fd_sc_hd__inv_2
XFILLER_72_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11872_ _11180_/X _11863_/X _11822_/B _11871_/X vssd1 vssd1 vccd1 vccd1 _21025_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_205_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13611_ _20393_/Q _13605_/X _13545_/X _13608_/X vssd1 vssd1 vccd1 vccd1 _20393_/D
+ sky130_fd_sc_hd__a22o_1
X_10823_ _10505_/X _10825_/A _10763_/A vssd1 vssd1 vccd1 vccd1 _10824_/C sky130_fd_sc_hd__o21a_1
X_14591_ _14591_/A _14591_/B vssd1 vssd1 vccd1 vccd1 _14605_/A sky130_fd_sc_hd__or2_1
XFILLER_25_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12065__B2 _20395_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18853__S _18907_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16330_ _19372_/Q _16326_/X _16235_/X _16328_/X vssd1 vssd1 vccd1 vccd1 _19372_/D
+ sky130_fd_sc_hd__a22o_1
X_13542_ _20428_/Q _13537_/X _13538_/X _13541_/X vssd1 vssd1 vccd1 vccd1 _20428_/D
+ sky130_fd_sc_hd__a22o_1
X_10754_ _10754_/A _10754_/B vssd1 vssd1 vccd1 vccd1 _10839_/A sky130_fd_sc_hd__or2_2
XFILLER_111_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17977__B _17978_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16261_ _16297_/A _16344_/B _16261_/C vssd1 vssd1 vccd1 vccd1 _16269_/A sky130_fd_sc_hd__or3_4
X_10685_ _10685_/A vssd1 vssd1 vccd1 vccd1 _10685_/X sky130_fd_sc_hd__buf_2
XANTENNA__13014__B1 _12925_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13473_ _13483_/A vssd1 vssd1 vccd1 vccd1 _13473_/X sky130_fd_sc_hd__buf_1
X_18000_ _18000_/A _18001_/B vssd1 vssd1 vccd1 vccd1 _18000_/Y sky130_fd_sc_hd__nor2_1
X_15212_ _20047_/Q _15211_/Y _15177_/A _15063_/B vssd1 vssd1 vccd1 vccd1 _20047_/D
+ sky130_fd_sc_hd__o211a_1
X_12424_ _12424_/A _12458_/A vssd1 vssd1 vccd1 vccd1 _12425_/B sky130_fd_sc_hd__or2_2
XFILLER_127_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16192_ _19438_/Q _16187_/X _16163_/X _16188_/X vssd1 vssd1 vccd1 vccd1 _19438_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_5_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15143_ _20454_/Q _15079_/A _20450_/Q _15075_/A _15142_/X vssd1 vssd1 vccd1 vccd1
+ _15144_/D sky130_fd_sc_hd__o221a_1
X_12355_ _12355_/A vssd1 vssd1 vccd1 vccd1 _12355_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19128__S0 _19285_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11306_ _11311_/A _11306_/B _11306_/C vssd1 vssd1 vccd1 vccd1 _11543_/C sky130_fd_sc_hd__or3_1
XFILLER_181_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15074_ _15074_/A _15074_/B vssd1 vssd1 vccd1 vccd1 _15188_/A sky130_fd_sc_hd__or2_1
X_12286_ _20936_/Q vssd1 vssd1 vccd1 vccd1 _12425_/A sky130_fd_sc_hd__inv_2
X_19951_ _21234_/CLK _19951_/D repeater270/X vssd1 vssd1 vccd1 vccd1 _19951_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11925__A1_N _21006_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11237_ _19911_/Q _19910_/Q vssd1 vssd1 vccd1 vccd1 _11250_/A sky130_fd_sc_hd__or2_2
X_18902_ _18901_/X _14146_/Y _18902_/S vssd1 vssd1 vccd1 vccd1 _18902_/X sky130_fd_sc_hd__mux2_1
X_14025_ _14013_/A _14013_/B _14023_/Y _14004_/A vssd1 vssd1 vccd1 vccd1 _20297_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_206_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19882_ _21334_/CLK _19882_/D repeater221/X vssd1 vssd1 vccd1 vccd1 _19882_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12930__A input46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18833_ _18832_/X _11916_/Y _18929_/S vssd1 vssd1 vccd1 vccd1 _18833_/X sky130_fd_sc_hd__mux2_1
X_11168_ _19110_/X vssd1 vssd1 vccd1 vccd1 _11176_/A sky130_fd_sc_hd__inv_2
XFILLER_121_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10119_ _20803_/Q vssd1 vssd1 vccd1 vccd1 _10119_/Y sky130_fd_sc_hd__inv_2
X_18764_ _18763_/X _10922_/Y _18928_/S vssd1 vssd1 vccd1 vccd1 _18764_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12828__B1 _12660_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15976_ _19547_/Q _15968_/X _15975_/X _15971_/X vssd1 vssd1 vccd1 vccd1 _19547_/D
+ sky130_fd_sc_hd__a22o_1
X_11099_ _21230_/Q _11099_/B vssd1 vssd1 vccd1 vccd1 _11099_/Y sky130_fd_sc_hd__nor2_1
XFILLER_222_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17715_ _21086_/Q vssd1 vssd1 vccd1 vccd1 _17715_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14927_ _20577_/Q _14960_/D _20570_/Q _15001_/A vssd1 vssd1 vccd1 vccd1 _14927_/X
+ sky130_fd_sc_hd__o22a_1
X_18695_ _17079_/Y _15261_/Y _18908_/S vssd1 vssd1 vccd1 vccd1 _18695_/X sky130_fd_sc_hd__mux2_1
XFILLER_224_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17646_ _17637_/Y _17301_/X _17640_/X _17645_/X vssd1 vssd1 vccd1 vccd1 _17646_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_36_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14858_ _15003_/A _15002_/A _15001_/A _14998_/A vssd1 vssd1 vccd1 vccd1 _14864_/C
+ sky130_fd_sc_hd__or4_4
XFILLER_212_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13809_ _20621_/Q _14587_/A _18004_/A _20198_/Q vssd1 vssd1 vccd1 vccd1 _13809_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__13253__B1 _13173_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17577_ _18746_/X _17907_/A _18744_/X _17908_/A vssd1 vssd1 vccd1 vccd1 _17577_/Y
+ sky130_fd_sc_hd__a22oi_4
XFILLER_16_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14789_ _19126_/X _14280_/X _14788_/X vssd1 vssd1 vccd1 vccd1 _20122_/D sky130_fd_sc_hd__a21oi_1
XANTENNA__18763__S _18927_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19316_ _20142_/CLK _19316_/D vssd1 vssd1 vccd1 vccd1 _19316_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_177_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16528_ _19984_/D vssd1 vssd1 vccd1 vccd1 _19986_/D sky130_fd_sc_hd__buf_1
XANTENNA__18192__A0 _18848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19247_ _17350_/Y _17351_/Y _17352_/Y _17353_/Y _20130_/Q _20131_/Q vssd1 vssd1 vccd1
+ vccd1 _19247_/X sky130_fd_sc_hd__mux4_1
XFILLER_177_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16459_ _16459_/A vssd1 vssd1 vccd1 vccd1 _16459_/X sky130_fd_sc_hd__buf_1
XFILLER_176_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18064__A _18064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19178_ _19545_/Q _19537_/Q _19529_/Q _19513_/Q _19280_/S0 _20122_/Q vssd1 vssd1
+ vccd1 vccd1 _19178_/X sky130_fd_sc_hd__mux4_1
XFILLER_129_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18129_ _18128_/X _12198_/Y _18909_/S vssd1 vssd1 vccd1 vccd1 _18129_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21140_ _21141_/CLK _21140_/D repeater192/X vssd1 vssd1 vccd1 vccd1 _21140_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__13001__A input55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21373__RESET_B repeater257/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21302__RESET_B repeater208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09902_ _21254_/Q vssd1 vssd1 vccd1 vccd1 _09902_/Y sky130_fd_sc_hd__inv_2
X_21071_ _21087_/CLK _21071_/D repeater227/X vssd1 vssd1 vccd1 vccd1 _21071_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__13936__A _20638_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16312__A _16319_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20022_ _21421_/CLK _20022_/D repeater214/X vssd1 vssd1 vccd1 vccd1 _20022_/Q sky130_fd_sc_hd__dfrtp_1
X_09833_ _15879_/A _09827_/X _09832_/X _09829_/X vssd1 vssd1 vccd1 vccd1 _21448_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_58_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18938__S _18946_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09764_ _21230_/Q vssd1 vssd1 vccd1 vccd1 _11055_/A sky130_fd_sc_hd__inv_2
XFILLER_100_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09695_ _21465_/Q _09690_/X _09693_/X _09694_/X vssd1 vssd1 vccd1 vccd1 _21465_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_2_0_0_HCLK_A clkbuf_2_1_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20924_ _20929_/CLK _20924_/D repeater267/X vssd1 vssd1 vccd1 vccd1 _20924_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_199_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_242_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20855_ _20857_/CLK _20855_/D repeater243/X vssd1 vssd1 vccd1 vccd1 _20855_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_42_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18673__S _18930_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13244__B1 _13243_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20786_ _21390_/CLK _20786_/D repeater239/X vssd1 vssd1 vccd1 vccd1 _20786_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09596__A _20889_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10470_ _10771_/A _20684_/Q _21283_/Q _10466_/Y _10469_/X vssd1 vssd1 vccd1 vccd1
+ _10471_/D sky130_fd_sc_hd__o221a_1
XFILLER_108_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21407_ _21407_/CLK _21407_/D repeater252/X vssd1 vssd1 vccd1 vccd1 _21407_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_135_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12140_ _20373_/Q vssd1 vssd1 vccd1 vccd1 _12140_/Y sky130_fd_sc_hd__inv_2
X_21338_ _21338_/CLK _21338_/D repeater221/X vssd1 vssd1 vccd1 vccd1 _21338_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_150_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12071_ _12316_/A _20377_/Q _12307_/A _20367_/Q vssd1 vssd1 vccd1 vccd1 _12071_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__19009__S _19019_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21269_ _21273_/CLK _21269_/D repeater246/X vssd1 vssd1 vccd1 vccd1 _21269_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_104_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11022_ _11590_/A _11022_/B vssd1 vssd1 vccd1 vccd1 _11022_/X sky130_fd_sc_hd__and2_1
XFILLER_238_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18848__S _18902_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15830_ _20137_/Q vssd1 vssd1 vccd1 vccd1 _16419_/A sky130_fd_sc_hd__buf_1
XFILLER_77_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15761_ _19645_/Q _15757_/X _15758_/X _15760_/X vssd1 vssd1 vccd1 vccd1 _19645_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_46_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12973_ _12973_/A vssd1 vssd1 vccd1 vccd1 _12981_/A sky130_fd_sc_hd__buf_1
X_17500_ _21020_/Q _17110_/Y _11878_/Y _19583_/Q vssd1 vssd1 vccd1 vccd1 _17500_/X
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__13581__A _13595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14712_ _14724_/A vssd1 vssd1 vccd1 vccd1 _14712_/X sky130_fd_sc_hd__buf_1
X_11924_ _16344_/A _11173_/B _16344_/A _11173_/B vssd1 vssd1 vccd1 vccd1 _11924_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_18480_ _18479_/X _14082_/A _18904_/S vssd1 vssd1 vccd1 vccd1 _18480_/X sky130_fd_sc_hd__mux2_1
X_15692_ _19676_/Q _15688_/X _15661_/X _15690_/X vssd1 vssd1 vccd1 vccd1 _19676_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17431_ _19344_/Q vssd1 vssd1 vccd1 vccd1 _17431_/Y sky130_fd_sc_hd__inv_2
XFILLER_82_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14643_ _20183_/Q _14641_/Y _14642_/X _14574_/B vssd1 vssd1 vccd1 vccd1 _20183_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_4573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13235__B1 _13151_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11855_ _11855_/A vssd1 vssd1 vccd1 vccd1 _11856_/B sky130_fd_sc_hd__inv_2
XANTENNA__18583__S _18885_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output105_A _17587_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10806_ _10773_/A _10773_/B _10795_/X _10804_/Y vssd1 vssd1 vccd1 vccd1 _21297_/D
+ sky130_fd_sc_hd__a211oi_2
X_17362_ _19327_/Q vssd1 vssd1 vccd1 vccd1 _17362_/Y sky130_fd_sc_hd__inv_2
XPHY_3872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14574_ _14574_/A _14574_/B vssd1 vssd1 vccd1 vccd1 _14637_/A sky130_fd_sc_hd__or2_2
XANTENNA__18174__A0 _17281_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11786_ _11786_/A _11786_/B _11786_/C vssd1 vssd1 vccd1 vccd1 _16596_/C sky130_fd_sc_hd__or3_1
XPHY_3883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19101_ _16669_/X _21077_/Q _19870_/D vssd1 vssd1 vccd1 vccd1 _19101_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16313_ _16319_/A vssd1 vssd1 vccd1 vccd1 _16320_/A sky130_fd_sc_hd__inv_2
X_13525_ _16515_/A _13182_/C _13530_/B _11160_/D _13524_/Y vssd1 vssd1 vccd1 vccd1
+ _13526_/A sky130_fd_sc_hd__o32a_1
X_17293_ _19841_/Q vssd1 vssd1 vccd1 vccd1 _17293_/Y sky130_fd_sc_hd__inv_2
XFILLER_159_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10737_ _19924_/Q _16769_/A vssd1 vssd1 vccd1 vccd1 _16773_/A sky130_fd_sc_hd__or2_1
XFILLER_13_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12925__A input48/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19032_ _16864_/X _20837_/Q _19046_/S vssd1 vssd1 vccd1 vccd1 _19944_/D sky130_fd_sc_hd__mux2_1
X_16244_ _19415_/Q _16240_/X _16014_/X _16241_/X vssd1 vssd1 vccd1 vccd1 _19415_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14735__B1 _13707_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13456_ _13657_/A _13456_/B vssd1 vssd1 vccd1 vccd1 _13491_/A sky130_fd_sc_hd__or2_2
X_10668_ _10668_/A _10668_/B vssd1 vssd1 vccd1 vccd1 _10669_/C sky130_fd_sc_hd__nor2_1
X_12407_ _12432_/C _12433_/A _12407_/C _12436_/A vssd1 vssd1 vccd1 vccd1 _12408_/C
+ sky130_fd_sc_hd__or4_4
X_16175_ _19449_/Q _16173_/X _16142_/X _16174_/X vssd1 vssd1 vccd1 vccd1 _19449_/D
+ sky130_fd_sc_hd__a22o_1
X_10599_ _10655_/A _20754_/Q _10660_/A _20759_/Q vssd1 vssd1 vccd1 vccd1 _10599_/X
+ sky130_fd_sc_hd__o22a_1
X_13387_ _13254_/X _20497_/Q _13387_/S vssd1 vssd1 vccd1 vccd1 _20497_/D sky130_fd_sc_hd__mux2_1
XFILLER_217_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput107 _17737_/Y vssd1 vssd1 vccd1 vccd1 HRDATA[6] sky130_fd_sc_hd__clkbuf_2
Xoutput118 _18120_/LO vssd1 vssd1 vccd1 vccd1 IRQ[15] sky130_fd_sc_hd__clkbuf_2
X_15126_ _15126_/A _15126_/B _15121_/X _15125_/X vssd1 vssd1 vccd1 vccd1 _15158_/B
+ sky130_fd_sc_hd__or4bb_4
Xoutput129 _21103_/Q vssd1 vssd1 vccd1 vccd1 MSO_S3 sky130_fd_sc_hd__clkbuf_2
X_12338_ _12333_/A _12333_/B _12376_/A _12334_/Y vssd1 vssd1 vccd1 vccd1 _20980_/D
+ sky130_fd_sc_hd__a211oi_4
XFILLER_99_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15057_ _20045_/Q vssd1 vssd1 vccd1 vccd1 _15060_/A sky130_fd_sc_hd__inv_2
X_19934_ _20841_/CLK _19934_/D repeater251/X vssd1 vssd1 vccd1 vccd1 _19934_/Q sky130_fd_sc_hd__dfrtp_1
X_12269_ _20948_/Q vssd1 vssd1 vccd1 vccd1 _12408_/A sky130_fd_sc_hd__inv_2
XANTENNA__12660__A input58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19861__RESET_B repeater226/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14008_ _13972_/C _13879_/B _14006_/Y _14004_/X vssd1 vssd1 vccd1 vccd1 _20303_/D
+ sky130_fd_sc_hd__a211oi_2
X_19865_ _21167_/CLK _19865_/D repeater225/X vssd1 vssd1 vccd1 vccd1 _19865_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_110_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18758__S _18927_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17988__B1 _18376_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18816_ _18815_/X _14072_/A _18850_/S vssd1 vssd1 vccd1 vccd1 _18816_/X sky130_fd_sc_hd__mux2_1
XFILLER_233_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19796_ _19820_/CLK _19796_/D vssd1 vssd1 vccd1 vccd1 _19796_/Q sky130_fd_sc_hd__dfxtp_1
X_18747_ _17542_/Y _21467_/Q _18897_/S vssd1 vssd1 vccd1 vccd1 _18747_/X sky130_fd_sc_hd__mux2_1
X_15959_ _19555_/Q _15954_/X _15893_/X _15956_/X vssd1 vssd1 vccd1 vccd1 _19555_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_95_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13474__B1 _13287_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18678_ _17754_/X _19589_/Q _18926_/S vssd1 vssd1 vccd1 vccd1 _18678_/X sky130_fd_sc_hd__mux2_1
XFILLER_224_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17629_ _20174_/Q _17368_/X _20175_/Q _17446_/X vssd1 vssd1 vccd1 vccd1 _17629_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_23_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18493__S _18908_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20640_ _20657_/CLK _20640_/D repeater198/X vssd1 vssd1 vccd1 vccd1 _20640_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_196_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11788__A0 _21042_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_220_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20571_ _20590_/CLK _20571_/D repeater258/X vssd1 vssd1 vccd1 vccd1 _20571_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_149_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12835__A _12841_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14726__B1 _13710_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19949__RESET_B repeater255/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21123_ _21125_/CLK _21123_/D repeater190/X vssd1 vssd1 vccd1 vccd1 _21123_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_121_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21054_ _21164_/CLK _21054_/D repeater225/X vssd1 vssd1 vccd1 vccd1 _21054_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_120_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_247_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18668__S _18896_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_219_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20005_ _21125_/CLK _20005_/D repeater190/X vssd1 vssd1 vccd1 vccd1 _20005_/Q sky130_fd_sc_hd__dfrtp_1
X_09816_ _15865_/A _09813_/X input74/X _09815_/X vssd1 vssd1 vccd1 vccd1 _21453_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_143_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_4_5_0_HCLK clkbuf_4_5_0_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_opt_3_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_100_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20436__RESET_B repeater278/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09747_ _20153_/Q vssd1 vssd1 vccd1 vccd1 _09747_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13465__B1 _13274_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19687__CLK _19765_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_227_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09678_ _15330_/A vssd1 vssd1 vccd1 vccd1 _09678_/X sky130_fd_sc_hd__buf_1
XPHY_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20907_ _20915_/CLK _20907_/D repeater217/X vssd1 vssd1 vccd1 vccd1 _20907_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11640_ _11640_/A vssd1 vssd1 vccd1 vccd1 _11640_/X sky130_fd_sc_hd__buf_1
XPHY_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20838_ _20930_/CLK _20838_/D repeater257/X vssd1 vssd1 vccd1 vccd1 _20838_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11571_ _13171_/A vssd1 vssd1 vccd1 vccd1 _11571_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_52_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20769_ _21319_/CLK _20769_/D repeater191/X vssd1 vssd1 vccd1 vccd1 _20769_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_22_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21295__RESET_B repeater208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13310_ _20540_/Q _13307_/X _13154_/X _13308_/X vssd1 vssd1 vccd1 vccd1 _20540_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_168_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10522_ _10522_/A _10522_/B _10522_/C _10522_/D vssd1 vssd1 vccd1 vccd1 _10523_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_52_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14290_ _19107_/X vssd1 vssd1 vccd1 vccd1 _14290_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21224__RESET_B repeater249/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10453_ _21307_/Q vssd1 vssd1 vccd1 vccd1 _10783_/A sky130_fd_sc_hd__inv_2
X_13241_ _13249_/A vssd1 vssd1 vccd1 vccd1 _13241_/X sky130_fd_sc_hd__buf_1
XFILLER_171_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13940__A1 _20638_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13172_ _20600_/Q _13165_/X _13171_/X _13167_/X vssd1 vssd1 vccd1 vccd1 _20600_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_input66_A HWDATA[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10384_ _10281_/A _10281_/B _10380_/Y _10383_/X vssd1 vssd1 vccd1 vccd1 _21366_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_184_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12123_ _20974_/Q _18029_/A _12306_/A _20366_/Q vssd1 vssd1 vccd1 vccd1 _12123_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_184_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17980_ _18033_/A vssd1 vssd1 vccd1 vccd1 _18001_/B sky130_fd_sc_hd__buf_4
XFILLER_97_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12054_ _20385_/Q vssd1 vssd1 vccd1 vccd1 _12054_/Y sky130_fd_sc_hd__inv_2
X_16931_ _16931_/A _16931_/B vssd1 vssd1 vccd1 vccd1 _16931_/Y sky130_fd_sc_hd__nor2_1
XFILLER_77_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18578__S _18667_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11005_ _11003_/X _11004_/Y _11003_/X _11004_/Y vssd1 vssd1 vccd1 vccd1 _11012_/C
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_238_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19650_ _19820_/CLK _19650_/D vssd1 vssd1 vccd1 vccd1 _19650_/Q sky130_fd_sc_hd__dfxtp_1
X_16862_ _16862_/A vssd1 vssd1 vccd1 vccd1 _16862_/Y sky130_fd_sc_hd__inv_2
XFILLER_238_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15813_ _19622_/Q _15807_/X _15812_/X _15808_/X vssd1 vssd1 vccd1 vccd1 _19622_/D
+ sky130_fd_sc_hd__a22o_1
X_18601_ _18600_/X _13925_/Y _18903_/S vssd1 vssd1 vccd1 vccd1 _18601_/X sky130_fd_sc_hd__mux2_1
XANTENNA__20177__RESET_B repeater200/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19581_ _21040_/CLK _19581_/D vssd1 vssd1 vccd1 vccd1 _19581_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16793_ _19929_/Q vssd1 vssd1 vccd1 vccd1 _16795_/A sky130_fd_sc_hd__inv_2
XFILLER_203_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18532_ _17944_/Y _16818_/Y _18875_/S vssd1 vssd1 vccd1 vccd1 _18532_/X sky130_fd_sc_hd__mux2_1
X_15744_ _15750_/A vssd1 vssd1 vccd1 vccd1 _15751_/A sky130_fd_sc_hd__inv_2
XANTENNA__20106__RESET_B repeater259/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12956_ _15385_/A vssd1 vssd1 vccd1 vccd1 _14264_/A sky130_fd_sc_hd__buf_4
XANTENNA__17198__B2 _17169_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_234_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18463_ _18462_/X _10765_/A _18617_/S vssd1 vssd1 vccd1 vccd1 _18463_/X sky130_fd_sc_hd__mux2_1
X_11907_ _21015_/Q vssd1 vssd1 vccd1 vccd1 _15397_/A sky130_fd_sc_hd__buf_1
XFILLER_45_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13208__B1 _13006_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15675_ _15681_/A vssd1 vssd1 vccd1 vccd1 _15682_/A sky130_fd_sc_hd__inv_2
XFILLER_234_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12887_ _12887_/A vssd1 vssd1 vccd1 vccd1 _12899_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_178_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17414_ _19409_/Q vssd1 vssd1 vccd1 vccd1 _17414_/Y sky130_fd_sc_hd__inv_2
XPHY_4392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14626_ _14581_/A _14581_/B _14621_/X _14623_/Y vssd1 vssd1 vccd1 vccd1 _20192_/D
+ sky130_fd_sc_hd__a211oi_2
X_11838_ _21034_/Q _11838_/B vssd1 vssd1 vccd1 vccd1 _11838_/Y sky130_fd_sc_hd__nor2_1
X_18394_ _18393_/X _13919_/Y _18849_/S vssd1 vssd1 vccd1 vccd1 _18394_/X sky130_fd_sc_hd__mux2_1
XFILLER_199_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_221_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17345_ _19400_/Q vssd1 vssd1 vccd1 vccd1 _17345_/Y sky130_fd_sc_hd__inv_2
X_14557_ _14557_/A vssd1 vssd1 vccd1 vccd1 _16405_/B sky130_fd_sc_hd__buf_1
X_11769_ _19086_/X _11764_/X _21048_/Q _11765_/X vssd1 vssd1 vccd1 vccd1 _21048_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_202_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13508_ _20440_/Q _13505_/X _13506_/X _13507_/X vssd1 vssd1 vccd1 vccd1 _20440_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14708__B1 _12853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_opt_4_HCLK clkbuf_opt_4_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_opt_4_HCLK/X
+ sky130_fd_sc_hd__clkbuf_16
X_17276_ _19334_/Q vssd1 vssd1 vccd1 vccd1 _17276_/Y sky130_fd_sc_hd__inv_2
X_14488_ _14488_/A vssd1 vssd1 vccd1 vccd1 _14488_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_leaf_133_HCLK_A clkbuf_4_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19015_ _16932_/X _20408_/Q _19019_/S vssd1 vssd1 vccd1 vccd1 _19961_/D sky130_fd_sc_hd__mux2_1
X_16227_ _19423_/Q _16223_/X _16125_/X _16224_/X vssd1 vssd1 vccd1 vccd1 _19423_/D
+ sky130_fd_sc_hd__a22o_1
X_13439_ _20471_/Q _13436_/X _13243_/X _13437_/X vssd1 vssd1 vccd1 vccd1 _20471_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17658__C1 _17657_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16158_ _16158_/A vssd1 vssd1 vccd1 vccd1 _16158_/X sky130_fd_sc_hd__buf_1
XFILLER_170_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15109_ _15107_/Y _20051_/Q _20438_/Q _15064_/A _15108_/X vssd1 vssd1 vccd1 vccd1
+ _15109_/X sky130_fd_sc_hd__o221a_1
XFILLER_115_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16089_ _19489_/Q _16087_/X _15876_/X _16088_/X vssd1 vssd1 vccd1 vccd1 _19489_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18870__A1 _19266_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19917_ _21055_/CLK _19917_/D repeater220/X vssd1 vssd1 vccd1 vccd1 _19917_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_142_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18488__S _18784_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13695__B1 _12860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19848_ _20042_/CLK _19848_/D repeater219/X vssd1 vssd1 vccd1 vccd1 _19850_/D sky130_fd_sc_hd__dfstp_1
XFILLER_228_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09601_ _12753_/A _10859_/B _14303_/C vssd1 vssd1 vccd1 vccd1 _17204_/A sky130_fd_sc_hd__or3_4
XFILLER_228_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19779_ _21009_/CLK _19779_/D vssd1 vssd1 vccd1 vccd1 _19779_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_243_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18138__A0 _18137_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_13_0_HCLK clkbuf_3_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_13_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_196_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20623_ _20623_/CLK _20623_/D repeater194/X vssd1 vssd1 vccd1 vccd1 _20623_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18951__S _18962_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12565__A _12580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20554_ _20592_/CLK _20554_/D repeater267/X vssd1 vssd1 vccd1 vccd1 _20554_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_164_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20485_ _20937_/CLK _20485_/D repeater277/X vssd1 vssd1 vccd1 vccd1 _20485_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_164_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_55_HCLK_A clkbuf_4_12_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11933__B1 _11932_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21106_ _21424_/CLK _21106_/D repeater230/X vssd1 vssd1 vccd1 vccd1 _21106_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_248_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18398__S _18880_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21037_ _21207_/CLK _21037_/D repeater242/X vssd1 vssd1 vccd1 vccd1 _21037_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20270__RESET_B repeater263/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13438__B1 _13240_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12810_ _12815_/A _13104_/B vssd1 vssd1 vccd1 vccd1 _12811_/S sky130_fd_sc_hd__or2_1
X_13790_ _20191_/Q vssd1 vssd1 vccd1 vccd1 _14580_/A sky130_fd_sc_hd__inv_2
XFILLER_170_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18377__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_216_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0_0_HCLK clkbuf_0_HCLK/X vssd1 vssd1 vccd1 vccd1 clkbuf_1_0_1_HCLK/A sky130_fd_sc_hd__clkbuf_1
X_12741_ _14674_/A vssd1 vssd1 vccd1 vccd1 _12743_/A sky130_fd_sc_hd__inv_2
XFILLER_231_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19022__S _19026_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21476__RESET_B repeater204/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15460_ _15460_/A vssd1 vssd1 vccd1 vccd1 _15460_/X sky130_fd_sc_hd__buf_1
XFILLER_231_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12672_ _12679_/A vssd1 vssd1 vccd1 vccd1 _12672_/X sky130_fd_sc_hd__buf_1
XPHY_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14411_ _21484_/Q vssd1 vssd1 vccd1 vccd1 _14411_/Y sky130_fd_sc_hd__inv_2
XPHY_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21405__RESET_B repeater252/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11623_ _21108_/Q _11623_/B vssd1 vssd1 vccd1 vccd1 _21108_/D sky130_fd_sc_hd__and2_1
XPHY_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15391_ _19817_/Q _15389_/X _15346_/X _15390_/X vssd1 vssd1 vccd1 vccd1 _19817_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13610__B1 _13543_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18861__S _18926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17130_ _20139_/Q vssd1 vssd1 vccd1 vccd1 _18112_/A sky130_fd_sc_hd__inv_2
XPHY_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14342_ _20223_/Q vssd1 vssd1 vccd1 vccd1 _14343_/A sky130_fd_sc_hd__inv_2
XFILLER_7_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11554_ _11566_/A vssd1 vssd1 vccd1 vccd1 _11554_/X sky130_fd_sc_hd__buf_1
XPHY_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19702__CLK _19706_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10505_ _10763_/B vssd1 vssd1 vccd1 vccd1 _10505_/X sky130_fd_sc_hd__buf_1
X_17061_ _20035_/Q _19838_/Q vssd1 vssd1 vccd1 vccd1 _17061_/X sky130_fd_sc_hd__and2_2
XFILLER_183_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15363__B1 _14262_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14273_ _15312_/A _17133_/B _17133_/A _14273_/D vssd1 vssd1 vccd1 vccd1 _14274_/S
+ sky130_fd_sc_hd__or4_4
X_11485_ _19106_/X _11480_/X _21152_/Q _11481_/X vssd1 vssd1 vccd1 vccd1 _21152_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_6_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16012_ _16012_/A vssd1 vssd1 vccd1 vccd1 _16012_/X sky130_fd_sc_hd__clkbuf_2
X_13224_ _20581_/Q _13215_/X _13223_/X _13217_/X vssd1 vssd1 vccd1 vccd1 _20581_/D
+ sky130_fd_sc_hd__a22o_1
X_10436_ _20695_/Q vssd1 vssd1 vccd1 vccd1 _18082_/A sky130_fd_sc_hd__inv_2
XANTENNA__18301__A0 _18848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_3_0_HCLK_A clkbuf_3_3_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13155_ _20609_/Q _13150_/X _13154_/X _13152_/X vssd1 vssd1 vccd1 vccd1 _20609_/D
+ sky130_fd_sc_hd__a22o_1
X_10367_ _10397_/A vssd1 vssd1 vccd1 vccd1 _10405_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA_repeater218_A repeater220/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12106_ _20977_/Q vssd1 vssd1 vccd1 vccd1 _12330_/A sky130_fd_sc_hd__inv_2
XFILLER_124_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17963_ _18048_/A vssd1 vssd1 vccd1 vccd1 _17963_/X sky130_fd_sc_hd__buf_1
XFILLER_88_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10298_ _21362_/Q _10295_/Y _10282_/A _20726_/Q _10297_/X vssd1 vssd1 vccd1 vccd1
+ _10307_/B sky130_fd_sc_hd__o221a_1
X_13086_ _13098_/A vssd1 vssd1 vccd1 vccd1 _13086_/X sky130_fd_sc_hd__buf_1
XFILLER_2_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19702_ _19706_/CLK _19702_/D vssd1 vssd1 vccd1 vccd1 _19702_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_214_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16914_ _16914_/A _16914_/B vssd1 vssd1 vccd1 vccd1 _16914_/Y sky130_fd_sc_hd__nor2_1
X_12037_ _20382_/Q vssd1 vssd1 vccd1 vccd1 _12037_/Y sky130_fd_sc_hd__inv_2
XFILLER_111_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17894_ _17974_/A vssd1 vssd1 vccd1 vccd1 _17898_/B sky130_fd_sc_hd__buf_4
XFILLER_66_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19633_ _21021_/CLK _19633_/D vssd1 vssd1 vccd1 vccd1 _19633_/Q sky130_fd_sc_hd__dfxtp_1
X_16845_ _19939_/Q _16834_/A _16829_/A _19940_/Q vssd1 vssd1 vccd1 vccd1 _16845_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_225_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16776_ _19925_/Q vssd1 vssd1 vccd1 vccd1 _16778_/A sky130_fd_sc_hd__inv_2
XFILLER_19_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19564_ _19706_/CLK _19564_/D vssd1 vssd1 vccd1 vccd1 _19564_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_230_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13988_ _13988_/A vssd1 vssd1 vccd1 vccd1 _13988_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_81_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15727_ _15737_/A vssd1 vssd1 vccd1 vccd1 _15727_/X sky130_fd_sc_hd__buf_1
X_18515_ _18514_/X _14097_/A _18850_/S vssd1 vssd1 vccd1 vccd1 _18515_/X sky130_fd_sc_hd__mux2_1
XFILLER_46_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12939_ _20717_/Q _12935_/X _12853_/X _12937_/X vssd1 vssd1 vccd1 vccd1 _20717_/D
+ sky130_fd_sc_hd__a22o_1
X_19495_ _20326_/CLK _19495_/D vssd1 vssd1 vccd1 vccd1 _19495_/Q sky130_fd_sc_hd__dfxtp_1
X_15658_ _15666_/A vssd1 vssd1 vccd1 vccd1 _15667_/A sky130_fd_sc_hd__inv_2
X_18446_ _18845_/A0 _10475_/Y _18884_/S vssd1 vssd1 vccd1 vccd1 _18446_/X sky130_fd_sc_hd__mux2_1
XFILLER_178_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14609_ _14609_/A vssd1 vssd1 vccd1 vccd1 _14609_/Y sky130_fd_sc_hd__inv_2
X_18377_ _18845_/A0 _17778_/Y _18879_/S vssd1 vssd1 vccd1 vccd1 _18377_/X sky130_fd_sc_hd__mux2_1
X_15589_ _19728_/Q _15584_/X _15588_/X _15586_/X vssd1 vssd1 vccd1 vccd1 _19728_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18771__S _18884_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17328_ _18920_/S _17312_/X _17318_/X _17322_/X _17327_/X vssd1 vssd1 vccd1 vccd1
+ _17328_/X sky130_fd_sc_hd__o2111a_1
XFILLER_193_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17895__B _17898_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17259_ _19318_/Q vssd1 vssd1 vccd1 vccd1 _17259_/Y sky130_fd_sc_hd__inv_2
XFILLER_146_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09694__A _15330_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19096__A1 _21082_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20270_ _20293_/CLK _20270_/D repeater263/X vssd1 vssd1 vccd1 vccd1 _20270_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__15106__B1 _20447_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19191__S1 _20124_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14105__A _20547_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20099__RESET_B repeater259/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20710__RESET_B repeater210/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18056__C1 _18055_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_245_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18946__S _18946_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_132_HCLK clkbuf_4_4_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20949_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_71_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12643__A1 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_213_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18681__S _18879_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19964__RESET_B repeater184/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20606_ _21302_/CLK _20606_/D repeater209/X vssd1 vssd1 vccd1 vccd1 _20606_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_138_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20537_ _20947_/CLK _20537_/D repeater267/X vssd1 vssd1 vccd1 vccd1 _20537_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_181_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19087__A1 _21059_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11270_ _12506_/A _11270_/B _11286_/C _11271_/C vssd1 vssd1 vccd1 vccd1 _11272_/A
+ sky130_fd_sc_hd__or4_4
X_20468_ _20937_/CLK _20468_/D repeater277/X vssd1 vssd1 vccd1 vccd1 _20468_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_106_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19182__S1 _20122_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10221_ _10221_/A _10221_/B _10221_/C vssd1 vssd1 vccd1 vccd1 _10224_/A sky130_fd_sc_hd__or3_4
XANTENNA__18834__A1 _19256_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20399_ _20809_/CLK _20399_/D repeater270/X vssd1 vssd1 vccd1 vccd1 _20399_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_133_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10152_ _10152_/A _10193_/A vssd1 vssd1 vccd1 vccd1 _10153_/B sky130_fd_sc_hd__or2_2
XFILLER_239_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19017__S _19019_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18047__C1 _18046_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17326__A _17928_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14960_ _14960_/A _14960_/B _14960_/C _14960_/D vssd1 vssd1 vccd1 vccd1 _14962_/C
+ sky130_fd_sc_hd__or4_4
X_10083_ _21401_/Q _10082_/Y _10162_/A _20798_/Q vssd1 vssd1 vccd1 vccd1 _10083_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_94_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold9 hold9/A vssd1 vssd1 vccd1 vccd1 hold9/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13911_ _20650_/Q vssd1 vssd1 vccd1 vccd1 _13911_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input29_A HADDR[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14891_ _20595_/Q vssd1 vssd1 vccd1 vccd1 _14891_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18856__S _18910_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16630_ _19880_/Q vssd1 vssd1 vccd1 vccd1 _17162_/A sky130_fd_sc_hd__inv_2
XFILLER_235_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10893__B1 _10892_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13842_ _20319_/Q vssd1 vssd1 vccd1 vccd1 _13894_/A sky130_fd_sc_hd__inv_2
X_16561_ _16561_/A vssd1 vssd1 vccd1 vccd1 _16561_/Y sky130_fd_sc_hd__inv_2
X_13773_ _13768_/Y _20206_/Q _20629_/Q _14595_/A _13772_/X vssd1 vssd1 vccd1 vccd1
+ _13786_/B sky130_fd_sc_hd__o221a_1
X_10985_ _10985_/A vssd1 vssd1 vccd1 vccd1 _10985_/Y sky130_fd_sc_hd__inv_2
X_18300_ _18299_/X _16966_/A _18680_/S vssd1 vssd1 vccd1 vccd1 _18300_/X sky130_fd_sc_hd__mux2_2
X_15512_ _19763_/Q _15507_/X _15456_/X _15509_/X vssd1 vssd1 vccd1 vccd1 _19763_/D
+ sky130_fd_sc_hd__a22o_1
X_19280_ _19307_/Q _19829_/Q _19837_/Q _19421_/Q _19280_/S0 _20122_/Q vssd1 vssd1
+ vccd1 vccd1 _19280_/X sky130_fd_sc_hd__mux4_2
X_12724_ _11179_/X _16915_/A _12724_/S vssd1 vssd1 vccd1 vccd1 _20809_/D sky130_fd_sc_hd__mux2_1
X_16492_ _20001_/Q vssd1 vssd1 vccd1 vccd1 _16503_/A sky130_fd_sc_hd__inv_2
XFILLER_43_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18231_ _20855_/Q input4/X _18236_/S vssd1 vssd1 vccd1 vccd1 _18231_/X sky130_fd_sc_hd__mux2_1
XFILLER_90_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15443_ _19793_/Q _15441_/X _15424_/X _15442_/X vssd1 vssd1 vccd1 vccd1 _19793_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12655_ _20842_/Q _12650_/X _12651_/X _12654_/X vssd1 vssd1 vccd1 vccd1 _20842_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_231_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18591__S _18896_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_repeater168_A _18874_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18162_ _18161_/X _20198_/Q _18748_/S vssd1 vssd1 vccd1 vccd1 _18162_/X sky130_fd_sc_hd__mux2_1
X_11606_ _18990_/X _11598_/A _21116_/Q _11605_/X vssd1 vssd1 vccd1 vccd1 _21116_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15374_ _16594_/B _15374_/B vssd1 vssd1 vccd1 vccd1 _15708_/C sky130_fd_sc_hd__or2_2
X_12586_ _20882_/Q _12581_/X _18234_/X _12583_/X vssd1 vssd1 vccd1 vccd1 _20882_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18522__A0 _17079_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17113_ _19598_/Q _17369_/B vssd1 vssd1 vccd1 vccd1 _17113_/Y sky130_fd_sc_hd__nor2_1
X_14325_ _14313_/Y _19120_/X _14311_/X _14324_/X vssd1 vssd1 vccd1 vccd1 _20241_/D
+ sky130_fd_sc_hd__o22ai_4
XPHY_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18093_ _18633_/X _17205_/X _18636_/X _17861_/A vssd1 vssd1 vccd1 vccd1 _18093_/X
+ sky130_fd_sc_hd__o22a_2
X_11537_ _21138_/Q _11534_/X _10896_/X _11535_/X vssd1 vssd1 vccd1 vccd1 _21138_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17044_ _19839_/Q vssd1 vssd1 vccd1 vccd1 _17044_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14256_ _14256_/A _14256_/B vssd1 vssd1 vccd1 vccd1 _14267_/A sky130_fd_sc_hd__or2_2
XFILLER_143_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output97_A _18059_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11468_ _11480_/A vssd1 vssd1 vccd1 vccd1 _11468_/X sky130_fd_sc_hd__buf_1
XANTENNA__20539__RESET_B repeater267/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_13_HCLK clkbuf_4_3_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _21121_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_125_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11549__A _11549_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13207_ _13217_/A vssd1 vssd1 vccd1 vccd1 _13207_/X sky130_fd_sc_hd__buf_1
XFILLER_171_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19173__S1 _20122_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18042__D _18042_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10419_ _21345_/Q _10418_/Y _10262_/B _10381_/X vssd1 vssd1 vccd1 vccd1 _21345_/D
+ sky130_fd_sc_hd__o211a_1
X_14187_ _14187_/A vssd1 vssd1 vccd1 vccd1 _14187_/Y sky130_fd_sc_hd__inv_2
X_11399_ _11418_/A vssd1 vssd1 vccd1 vccd1 _11402_/B sky130_fd_sc_hd__inv_2
XFILLER_225_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20192__RESET_B repeater200/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13138_ _13138_/A vssd1 vssd1 vccd1 vccd1 _13165_/A sky130_fd_sc_hd__buf_1
X_18995_ _17016_/X _20428_/Q _19026_/S vssd1 vssd1 vccd1 vccd1 _19981_/D sky130_fd_sc_hd__mux2_1
XFILLER_86_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13764__A _20612_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20121__RESET_B repeater247/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_239_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17946_ _20414_/Q _18007_/B vssd1 vssd1 vccd1 vccd1 _17946_/Y sky130_fd_sc_hd__nand2_1
X_13069_ _20656_/Q _13066_/X _12918_/X _13067_/X vssd1 vssd1 vccd1 vccd1 _20656_/D
+ sky130_fd_sc_hd__a22o_1
Xrepeater204 repeater205/X vssd1 vssd1 vccd1 vccd1 repeater204/X sky130_fd_sc_hd__buf_8
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater215 repeater232/X vssd1 vssd1 vccd1 vccd1 repeater215/X sky130_fd_sc_hd__buf_8
Xrepeater226 repeater227/X vssd1 vssd1 vccd1 vccd1 repeater226/X sky130_fd_sc_hd__buf_8
Xclkbuf_leaf_155_HCLK clkbuf_opt_1_HCLK/A vssd1 vssd1 vccd1 vccd1 _21040_/CLK sky130_fd_sc_hd__clkbuf_16
Xrepeater237 repeater238/X vssd1 vssd1 vccd1 vccd1 repeater237/X sky130_fd_sc_hd__buf_8
XFILLER_94_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12873__A1 _20742_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17877_ _20409_/Q vssd1 vssd1 vccd1 vccd1 _17877_/Y sky130_fd_sc_hd__inv_2
Xrepeater248 repeater249/X vssd1 vssd1 vccd1 vccd1 repeater248/X sky130_fd_sc_hd__buf_8
XANTENNA__18766__S _18930_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater259 repeater260/X vssd1 vssd1 vccd1 vccd1 repeater259/X sky130_fd_sc_hd__buf_8
X_19616_ _20137_/CLK _19616_/D vssd1 vssd1 vccd1 vccd1 _19616_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_241_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16828_ _16843_/B vssd1 vssd1 vccd1 vccd1 _16829_/A sky130_fd_sc_hd__buf_1
XANTENNA__17800__A2 _18045_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19547_ _21462_/CLK _19547_/D vssd1 vssd1 vccd1 vccd1 _19547_/Q sky130_fd_sc_hd__dfxtp_1
X_16759_ _19921_/Q vssd1 vssd1 vccd1 vccd1 _16759_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19478_ _19961_/CLK _19478_/D vssd1 vssd1 vccd1 vccd1 _19478_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18429_ _18845_/A0 _10326_/Y _18884_/S vssd1 vssd1 vccd1 vccd1 _18429_/X sky130_fd_sc_hd__mux2_1
XFILLER_221_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21440_ _21459_/CLK _21440_/D repeater244/X vssd1 vssd1 vccd1 vccd1 _21440_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18513__A0 _18848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21371_ _21374_/CLK _21371_/D repeater255/X vssd1 vssd1 vccd1 vccd1 _21371_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__15327__B1 _13547_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20962__RESET_B repeater186/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20322_ _20322_/CLK _20322_/D repeater262/X vssd1 vssd1 vccd1 vccd1 _20322_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__19069__A1 _21141_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20253_ _20908_/CLK _20253_/D repeater217/X vssd1 vssd1 vccd1 vccd1 _20253_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__19164__S1 _20122_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20209__RESET_B repeater203/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20184_ _21483_/CLK _20184_/D repeater194/X vssd1 vssd1 vccd1 vccd1 _20184_/Q sky130_fd_sc_hd__dfrtp_1
X_09995_ _20022_/Q _09988_/B _09994_/Y _20023_/Q _09988_/Y vssd1 vssd1 vccd1 vccd1
+ _20023_/D sky130_fd_sc_hd__a32o_1
XFILLER_142_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17146__A _17290_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13674__A _13680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18676__S _18930_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_217_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10875__B1 _09698_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09599__A _19982_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10770_ _10770_/A _10811_/A vssd1 vssd1 vccd1 vccd1 _10771_/B sky130_fd_sc_hd__or2_2
XANTENNA__18752__A0 _18751_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_213_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15566__B1 _15550_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12440_ _12440_/A vssd1 vssd1 vccd1 vccd1 _12440_/Y sky130_fd_sc_hd__inv_2
XFILLER_166_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_226_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_36_HCLK _20004_/CLK vssd1 vssd1 vccd1 vccd1 _21167_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_166_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12371_ _12093_/X _12315_/B _12364_/X _12369_/Y vssd1 vssd1 vccd1 vccd1 _20962_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_5_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14110_ _20549_/Q _14088_/A _17897_/A _20273_/Q vssd1 vssd1 vccd1 vccd1 _14110_/X
+ sky130_fd_sc_hd__o22a_1
X_11322_ _11322_/A _11322_/B vssd1 vssd1 vccd1 vccd1 _11322_/Y sky130_fd_sc_hd__nor2_1
XFILLER_176_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15090_ _20075_/Q vssd1 vssd1 vccd1 vccd1 _15090_/Y sky130_fd_sc_hd__inv_2
XFILLER_176_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19155__S1 _21017_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14041_ _20287_/Q vssd1 vssd1 vccd1 vccd1 _14097_/A sky130_fd_sc_hd__inv_2
X_11253_ _19064_/X _11250_/X _21188_/Q _11251_/X vssd1 vssd1 vccd1 vccd1 _21188_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_181_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12552__B1 _11733_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10204_ _10204_/A _10213_/A vssd1 vssd1 vccd1 vccd1 _10205_/B sky130_fd_sc_hd__or2_2
XFILLER_79_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11184_ _17290_/A _15847_/A vssd1 vssd1 vccd1 vccd1 _17684_/A sky130_fd_sc_hd__or2_4
XFILLER_121_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13584__A input69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17800_ _18398_/X _18045_/A _18401_/X _18048_/A _17799_/X vssd1 vssd1 vccd1 vccd1
+ _17800_/X sky130_fd_sc_hd__o221a_1
XFILLER_192_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10135_ _10150_/A _20786_/Q _21389_/Q _10132_/Y _10134_/X vssd1 vssd1 vccd1 vccd1
+ _10136_/D sky130_fd_sc_hd__o221a_1
X_15992_ _19538_/Q _15986_/X _15941_/X _15988_/X vssd1 vssd1 vccd1 vccd1 _19538_/D
+ sky130_fd_sc_hd__a22o_1
X_18780_ _18848_/A0 _14156_/Y _18902_/S vssd1 vssd1 vccd1 vccd1 _18780_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14943_ _20593_/Q _14881_/A _14942_/Y _20081_/Q vssd1 vssd1 vccd1 vccd1 _14943_/X
+ sky130_fd_sc_hd__o22a_1
X_10066_ _21392_/Q vssd1 vssd1 vccd1 vccd1 _10153_/A sky130_fd_sc_hd__inv_2
XFILLER_121_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17731_ _18688_/X _17397_/X _18685_/X _17398_/X _17730_/X vssd1 vssd1 vccd1 vccd1
+ _17731_/X sky130_fd_sc_hd__o221a_1
XANTENNA_output135_A _17043_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18586__S _18784_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14874_ _14960_/B _14874_/B vssd1 vssd1 vccd1 vccd1 _14981_/A sky130_fd_sc_hd__or2_1
X_17662_ _18065_/A vssd1 vssd1 vccd1 vccd1 _17856_/A sky130_fd_sc_hd__buf_2
XFILLER_29_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19401_ _19813_/CLK _19401_/D vssd1 vssd1 vccd1 vccd1 _19401_/Q sky130_fd_sc_hd__dfxtp_1
X_16613_ _19988_/Q vssd1 vssd1 vccd1 vccd1 _16613_/Y sky130_fd_sc_hd__inv_2
X_13825_ _20615_/Q vssd1 vssd1 vccd1 vccd1 _13825_/Y sky130_fd_sc_hd__inv_2
XFILLER_235_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12607__A1 _17060_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17593_ _19427_/Q vssd1 vssd1 vccd1 vccd1 _17593_/Y sky130_fd_sc_hd__inv_2
XFILLER_211_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12607__B2 _12601_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12928__A input47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16544_ _21149_/Q _21148_/Q vssd1 vssd1 vccd1 vccd1 _19879_/D sky130_fd_sc_hd__or2_1
X_19332_ _19834_/CLK _19332_/D vssd1 vssd1 vccd1 vccd1 _19332_/Q sky130_fd_sc_hd__dfxtp_1
X_13756_ _20181_/Q vssd1 vssd1 vccd1 vccd1 _14571_/A sky130_fd_sc_hd__inv_2
X_10968_ _10962_/Y _21026_/Q _21199_/Q _10964_/X _10967_/X vssd1 vssd1 vccd1 vccd1
+ _10969_/D sky130_fd_sc_hd__o221a_1
XANTENNA__11551__B _14273_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12707_ _12707_/A vssd1 vssd1 vccd1 vccd1 _12707_/X sky130_fd_sc_hd__buf_1
XFILLER_203_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16475_ _19295_/Q _16473_/X _16288_/X _16474_/X vssd1 vssd1 vccd1 vccd1 _19295_/D
+ sky130_fd_sc_hd__a22o_1
X_19263_ _17240_/Y _17241_/Y _17242_/Y _17243_/Y _19275_/S0 _21004_/Q vssd1 vssd1
+ vccd1 vccd1 _19263_/X sky130_fd_sc_hd__mux4_1
X_13687_ _13687_/A vssd1 vssd1 vccd1 vccd1 _13708_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_188_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10899_ _21251_/Q _10888_/A _10898_/X _10890_/A vssd1 vssd1 vccd1 vccd1 _21251_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_231_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15426_ _19801_/Q _15423_/X _15424_/X _15425_/X vssd1 vssd1 vccd1 vccd1 _19801_/D
+ sky130_fd_sc_hd__a22o_1
X_18214_ _18848_/A0 _14159_/Y _18902_/S vssd1 vssd1 vccd1 vccd1 _18214_/X sky130_fd_sc_hd__mux2_1
X_12638_ _12638_/A vssd1 vssd1 vccd1 vccd1 _12638_/X sky130_fd_sc_hd__buf_1
XPHY_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19194_ _19732_/Q _19372_/Q _19788_/Q _19772_/Q _19280_/S0 _20122_/Q vssd1 vssd1
+ vccd1 vccd1 _19194_/X sky130_fd_sc_hd__mux4_1
XPHY_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15357_ _15574_/A _15357_/B _16481_/A vssd1 vssd1 vccd1 vccd1 _16325_/C sky130_fd_sc_hd__or3_4
X_18145_ _18845_/A0 _10324_/Y _18884_/S vssd1 vssd1 vccd1 vccd1 _18145_/X sky130_fd_sc_hd__mux2_1
X_12569_ _12582_/A vssd1 vssd1 vccd1 vccd1 _12575_/A sky130_fd_sc_hd__buf_1
XANTENNA__12663__A input57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14308_ _14308_/A vssd1 vssd1 vccd1 vccd1 _14309_/B sky130_fd_sc_hd__buf_1
XFILLER_8_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20373__RESET_B repeater186/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18076_ _17925_/A _18076_/B _18076_/C vssd1 vssd1 vccd1 vccd1 _18076_/Y sky130_fd_sc_hd__nand3b_4
X_15288_ _19854_/Q _15288_/B vssd1 vssd1 vccd1 vccd1 _15289_/B sky130_fd_sc_hd__or2_1
X_17027_ _17027_/A _21243_/Q vssd1 vssd1 vccd1 vccd1 _17027_/Y sky130_fd_sc_hd__nor2_1
X_14239_ _19899_/Q _14239_/B vssd1 vssd1 vccd1 vccd1 _14240_/B sky130_fd_sc_hd__or2_1
XFILLER_112_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09780_ _09780_/A vssd1 vssd1 vccd1 vccd1 _16620_/A sky130_fd_sc_hd__buf_1
XFILLER_86_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18978_ _21428_/Q _21101_/Q _18983_/S vssd1 vssd1 vccd1 vccd1 _18978_/X sky130_fd_sc_hd__mux2_1
XFILLER_239_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17929_ _18510_/X _17928_/X _18504_/X _17214_/X vssd1 vssd1 vccd1 vccd1 _17929_/X
+ sky130_fd_sc_hd__o22a_2
XANTENNA__18496__S _18908_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_239_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20940_ _20950_/CLK _20940_/D repeater272/X vssd1 vssd1 vccd1 vccd1 _20940_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_66_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__21161__RESET_B repeater226/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_242_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15796__B1 _15795_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20871_ _21438_/CLK _20871_/D repeater237/X vssd1 vssd1 vccd1 vccd1 _20871_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_81_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_6_0_HCLK_A clkbuf_4_7_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_59_HCLK clkbuf_4_14_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _21306_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_179_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21423_ _21423_/CLK _21423_/D repeater231/X vssd1 vssd1 vccd1 vccd1 _21423_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_175_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12782__B1 _09638_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13388__B _13456_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21354_ _21368_/CLK _21354_/D repeater252/X vssd1 vssd1 vccd1 vccd1 _21354_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_163_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20305_ _20693_/CLK _20305_/D repeater196/X vssd1 vssd1 vccd1 vccd1 _20305_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__19137__S1 _21017_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15884__A _15884_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20043__RESET_B repeater276/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21285_ _21306_/CLK _21285_/D repeater207/X vssd1 vssd1 vccd1 vccd1 _21285_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_190_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20236_ _21477_/CLK _20236_/D repeater204/X vssd1 vssd1 vccd1 vccd1 _20236_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_115_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20167_ _21011_/CLK _20167_/D repeater237/X vssd1 vssd1 vccd1 vccd1 _20167_/Q sky130_fd_sc_hd__dfrtp_1
X_09978_ _21416_/Q _09975_/X _09685_/X _09976_/X vssd1 vssd1 vccd1 vccd1 _21416_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_130_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20098_ _20101_/CLK _20098_/D repeater259/X vssd1 vssd1 vccd1 vccd1 _20098_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_92_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11940_ _11940_/A _11940_/B vssd1 vssd1 vccd1 vccd1 _11940_/Y sky130_fd_sc_hd__nor2_1
XFILLER_176_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11871_ _21025_/Q _10934_/X _11863_/X _11864_/X vssd1 vssd1 vccd1 vccd1 _11871_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_232_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13610_ _20394_/Q _13605_/X _13543_/X _13608_/X vssd1 vssd1 vccd1 vccd1 _20394_/D
+ sky130_fd_sc_hd__a22o_1
X_10822_ _21288_/Q _10824_/B _10812_/X _10765_/B vssd1 vssd1 vccd1 vccd1 _21288_/D
+ sky130_fd_sc_hd__o211a_1
X_14590_ _14590_/A _14609_/A vssd1 vssd1 vccd1 vccd1 _14591_/B sky130_fd_sc_hd__or2_1
XFILLER_26_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18725__A0 _17079_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13541_ _13567_/A vssd1 vssd1 vccd1 vccd1 _13541_/X sky130_fd_sc_hd__buf_1
X_10753_ _21309_/Q _10752_/X _10731_/Y vssd1 vssd1 vccd1 vccd1 _21309_/D sky130_fd_sc_hd__o21a_1
XFILLER_197_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20884__RESET_B repeater243/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19030__S _19046_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16260_ _19406_/Q _16255_/X _16127_/X _16256_/X vssd1 vssd1 vccd1 vccd1 _19406_/D
+ sky130_fd_sc_hd__a22o_1
X_13472_ _13481_/A vssd1 vssd1 vccd1 vccd1 _13472_/X sky130_fd_sc_hd__buf_1
XFILLER_200_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10684_ _21331_/Q _10683_/Y _10680_/X _10661_/B vssd1 vssd1 vccd1 vccd1 _21331_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__20813__RESET_B repeater212/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15211_ _15211_/A vssd1 vssd1 vccd1 vccd1 _15211_/Y sky130_fd_sc_hd__inv_2
XFILLER_185_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12423_ _12423_/A _12423_/B vssd1 vssd1 vccd1 vccd1 _12458_/A sky130_fd_sc_hd__or2_1
X_16191_ _19439_/Q _16187_/X _16147_/X _16188_/X vssd1 vssd1 vccd1 vccd1 _19439_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14762__B2 _20130_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12773__B1 _12673_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15142_ _15141_/Y _20059_/Q _20448_/Q _15073_/A vssd1 vssd1 vccd1 vccd1 _15142_/X
+ sky130_fd_sc_hd__o22a_1
X_12354_ _12325_/A _12325_/B _12350_/X _12352_/Y vssd1 vssd1 vccd1 vccd1 _20972_/D
+ sky130_fd_sc_hd__a211oi_2
X_11305_ _20902_/Q vssd1 vssd1 vccd1 vccd1 _11307_/B sky130_fd_sc_hd__inv_2
XANTENNA__19128__S1 _21017_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15073_ _15073_/A _15191_/A vssd1 vssd1 vccd1 vccd1 _15074_/B sky130_fd_sc_hd__or2_2
X_19950_ _20809_/CLK _19950_/D repeater189/X vssd1 vssd1 vccd1 vccd1 _19950_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_5_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12285_ _20921_/Q vssd1 vssd1 vccd1 vccd1 _12396_/A sky130_fd_sc_hd__inv_2
XFILLER_181_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18901_ _18900_/X _17176_/Y _18901_/S vssd1 vssd1 vccd1 vccd1 _18901_/X sky130_fd_sc_hd__mux2_1
X_14024_ _20298_/Q _14023_/Y _14015_/B _13965_/X vssd1 vssd1 vccd1 vccd1 _20298_/D
+ sky130_fd_sc_hd__o211a_1
X_11236_ _21196_/Q _11235_/A _11234_/Y _11235_/Y _19910_/Q vssd1 vssd1 vccd1 vccd1
+ _21196_/D sky130_fd_sc_hd__a221o_1
XFILLER_107_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19881_ _21185_/CLK _19881_/D repeater221/X vssd1 vssd1 vccd1 vccd1 _19881_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_150_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18832_ _18831_/X _10962_/Y _18928_/S vssd1 vssd1 vccd1 vccd1 _18832_/X sky130_fd_sc_hd__mux2_1
X_11167_ _16465_/A vssd1 vssd1 vccd1 vccd1 _15610_/A sky130_fd_sc_hd__buf_1
XFILLER_67_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10118_ _10157_/A _20793_/Q _10162_/C _20799_/Q _10117_/Y vssd1 vssd1 vccd1 vccd1
+ _10122_/C sky130_fd_sc_hd__o221a_1
XFILLER_121_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18763_ _18762_/X _17506_/Y _18927_/S vssd1 vssd1 vccd1 vccd1 _18763_/X sky130_fd_sc_hd__mux2_1
X_15975_ _16237_/A vssd1 vssd1 vccd1 vccd1 _15975_/X sky130_fd_sc_hd__buf_1
X_11098_ _11098_/A vssd1 vssd1 vccd1 vccd1 _11099_/B sky130_fd_sc_hd__inv_2
XFILLER_236_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17714_ _17712_/Y _17639_/X _17713_/Y _17142_/A vssd1 vssd1 vccd1 vccd1 _17714_/X
+ sky130_fd_sc_hd__o22a_1
X_14926_ _20572_/Q vssd1 vssd1 vccd1 vccd1 _14926_/Y sky130_fd_sc_hd__inv_2
X_10049_ _10049_/A vssd1 vssd1 vccd1 vccd1 _10205_/A sky130_fd_sc_hd__buf_1
XFILLER_63_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18694_ _18693_/X _14076_/A _18850_/S vssd1 vssd1 vccd1 vccd1 _18694_/X sky130_fd_sc_hd__mux2_1
XFILLER_209_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17645_ _17641_/Y _17290_/X _17642_/Y _17292_/X _17644_/X vssd1 vssd1 vccd1 vccd1
+ _17645_/X sky130_fd_sc_hd__o221a_1
X_14857_ _20076_/Q vssd1 vssd1 vccd1 vccd1 _14998_/A sky130_fd_sc_hd__inv_2
XANTENNA__12658__A input59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13808_ _20621_/Q vssd1 vssd1 vccd1 vccd1 _18004_/A sky130_fd_sc_hd__inv_2
XANTENNA__18716__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14788_ _14783_/A _14288_/X _14279_/A vssd1 vssd1 vccd1 vccd1 _14788_/X sky130_fd_sc_hd__o21a_1
X_17576_ _17576_/A vssd1 vssd1 vccd1 vccd1 _17908_/A sky130_fd_sc_hd__clkbuf_2
X_19315_ _20142_/CLK _19315_/D vssd1 vssd1 vccd1 vccd1 _19315_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_220_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13739_ _20607_/Q vssd1 vssd1 vccd1 vccd1 _17810_/A sky130_fd_sc_hd__inv_2
XANTENNA__15969__A _16231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16527_ _19984_/D _16527_/B vssd1 vssd1 vccd1 vccd1 _19983_/D sky130_fd_sc_hd__or2_1
XFILLER_189_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19246_ _19242_/X _19243_/X _19244_/X _19245_/X _21005_/Q _21006_/Q vssd1 vssd1 vccd1
+ vccd1 _19246_/X sky130_fd_sc_hd__mux4_2
XFILLER_32_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16458_ _19304_/Q _16452_/X _16332_/X _16454_/X vssd1 vssd1 vccd1 vccd1 _19304_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__20554__RESET_B repeater267/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13489__A input45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15409_ _19807_/Q _15405_/X _15352_/X _15406_/X vssd1 vssd1 vccd1 vccd1 _19807_/D
+ sky130_fd_sc_hd__a22o_1
X_16389_ _19342_/Q _16385_/X _16212_/X _16386_/X vssd1 vssd1 vccd1 vccd1 _19342_/D
+ sky130_fd_sc_hd__a22o_1
X_19177_ _19705_/Q _19569_/Q _19561_/Q _19553_/Q _19280_/S0 _20122_/Q vssd1 vssd1
+ vccd1 vccd1 _19177_/X sky130_fd_sc_hd__mux4_2
XANTENNA__15950__B1 _15949_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12764__B1 _12660_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18128_ _17079_/Y _12045_/Y _18908_/S vssd1 vssd1 vccd1 vccd1 _18128_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18059_ _18018_/X _18059_/B _18059_/C vssd1 vssd1 vccd1 vccd1 _18059_/Y sky130_fd_sc_hd__nand3b_4
XFILLER_172_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09901_ _09898_/X _09899_/X _20008_/Q _09900_/Y vssd1 vssd1 vccd1 vccd1 _17022_/A
+ sky130_fd_sc_hd__a31o_1
X_21070_ _21087_/CLK _21070_/D repeater228/X vssd1 vssd1 vccd1 vccd1 _21070_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_160_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20021_ _21419_/CLK _20021_/D repeater232/X vssd1 vssd1 vccd1 vccd1 _20021_/Q sky130_fd_sc_hd__dfrtp_1
X_09832_ _15876_/A vssd1 vssd1 vccd1 vccd1 _09832_/X sky130_fd_sc_hd__buf_1
XFILLER_140_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14269__B1 _13707_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_246_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__21342__RESET_B repeater211/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09763_ _21224_/Q vssd1 vssd1 vccd1 vccd1 _11113_/A sky130_fd_sc_hd__inv_2
XFILLER_246_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09694_ _15330_/A vssd1 vssd1 vccd1 vccd1 _09694_/X sky130_fd_sc_hd__buf_1
XFILLER_26_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20923_ _20930_/CLK _20923_/D repeater268/X vssd1 vssd1 vccd1 vccd1 _20923_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_54_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18954__S _18962_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12568__A _12580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_214_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_242_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20854_ _20857_/CLK _20854_/D repeater243/X vssd1 vssd1 vccd1 vccd1 _20854_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20785_ _21390_/CLK _20785_/D repeater239/X vssd1 vssd1 vccd1 vccd1 _20785_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20295__RESET_B repeater262/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20224__RESET_B repeater202/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21406_ _21406_/CLK _21406_/D repeater213/X vssd1 vssd1 vccd1 vccd1 _21406_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_108_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21337_ _21476_/CLK _21337_/D repeater204/X vssd1 vssd1 vccd1 vccd1 _21337_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_150_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12070_ _20953_/Q vssd1 vssd1 vccd1 vccd1 _12307_/A sky130_fd_sc_hd__inv_2
X_21268_ _21433_/CLK _21268_/D repeater236/X vssd1 vssd1 vccd1 vccd1 _21268_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_132_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11021_ _21241_/Q _11021_/B vssd1 vssd1 vccd1 vccd1 _11022_/B sky130_fd_sc_hd__nand2_1
X_20219_ _20220_/CLK _20219_/D repeater202/X vssd1 vssd1 vccd1 vccd1 _20219_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_238_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21199_ _21390_/CLK _21199_/D repeater240/X vssd1 vssd1 vccd1 vccd1 _21199_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_106_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19025__S _19026_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21012__RESET_B repeater238/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15760_ _15770_/A vssd1 vssd1 vccd1 vccd1 _15760_/X sky130_fd_sc_hd__buf_1
XFILLER_45_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12972_ _12966_/X _12970_/X _14686_/A _12969_/X vssd1 vssd1 vccd1 vccd1 _20701_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_66_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input11_A HADDR[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14711_ _14723_/A vssd1 vssd1 vccd1 vccd1 _14711_/X sky130_fd_sc_hd__buf_1
XFILLER_73_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11923_ _21222_/Q vssd1 vssd1 vccd1 vccd1 _16344_/A sky130_fd_sc_hd__buf_1
X_15691_ _19677_/Q _15688_/X _15657_/X _15690_/X vssd1 vssd1 vccd1 vccd1 _19677_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_45_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18864__S _18929_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14642_ _14642_/A vssd1 vssd1 vccd1 vccd1 _14642_/X sky130_fd_sc_hd__clkbuf_2
X_17430_ _19320_/Q vssd1 vssd1 vccd1 vccd1 _17430_/Y sky130_fd_sc_hd__inv_2
XPHY_4563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11854_ _11854_/A vssd1 vssd1 vccd1 vccd1 _21030_/D sky130_fd_sc_hd__inv_2
XPHY_4574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10805_ _21298_/Q _10804_/Y _10798_/X _10775_/B vssd1 vssd1 vccd1 vccd1 _21298_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_202_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14573_ _14573_/A _14641_/A vssd1 vssd1 vccd1 vccd1 _14574_/B sky130_fd_sc_hd__or2_2
X_17361_ _19351_/Q vssd1 vssd1 vccd1 vccd1 _17361_/Y sky130_fd_sc_hd__inv_2
X_11785_ _11357_/A _11784_/X _11376_/C vssd1 vssd1 vccd1 vccd1 _11786_/B sky130_fd_sc_hd__o21ai_1
XPHY_3873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19100_ _16670_/X _21078_/Q _19870_/D vssd1 vssd1 vccd1 vccd1 _19100_/X sky130_fd_sc_hd__mux2_1
XFILLER_41_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12994__B1 _12993_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16312_ _16319_/A vssd1 vssd1 vccd1 vccd1 _16312_/X sky130_fd_sc_hd__buf_1
X_13524_ _13528_/C _13524_/B vssd1 vssd1 vccd1 vccd1 _13524_/Y sky130_fd_sc_hd__nor2_1
X_17292_ _17292_/A vssd1 vssd1 vccd1 vccd1 _17292_/X sky130_fd_sc_hd__buf_1
X_10736_ _19923_/Q _16765_/A vssd1 vssd1 vccd1 vccd1 _16769_/A sky130_fd_sc_hd__or2_1
XFILLER_14_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16243_ _19416_/Q _16240_/X _16012_/X _16241_/X vssd1 vssd1 vccd1 vccd1 _19416_/D
+ sky130_fd_sc_hd__a22o_1
X_19031_ _16866_/X _20838_/Q _19046_/S vssd1 vssd1 vccd1 vccd1 _19945_/D sky130_fd_sc_hd__mux2_1
XFILLER_174_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13455_ _20465_/Q _13444_/X _13454_/X _13447_/X vssd1 vssd1 vccd1 vccd1 _20465_/D
+ sky130_fd_sc_hd__a22o_1
X_10667_ _21339_/Q _10666_/Y _10574_/C _10666_/A _10642_/X vssd1 vssd1 vccd1 vccd1
+ _21339_/D sky130_fd_sc_hd__o221a_1
XANTENNA_repeater150_A _18884_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15932__B1 _15795_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_repeater248_A repeater249/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12406_ _12418_/B _12406_/B _12406_/C vssd1 vssd1 vccd1 vccd1 _12436_/A sky130_fd_sc_hd__or3_1
X_16174_ _16174_/A vssd1 vssd1 vccd1 vccd1 _16174_/X sky130_fd_sc_hd__buf_1
XFILLER_127_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13386_ _13456_/B _17174_/B vssd1 vssd1 vccd1 vccd1 _13387_/S sky130_fd_sc_hd__or2_1
X_10598_ _21318_/Q _10596_/Y _10706_/A _20746_/Q _10597_/X vssd1 vssd1 vccd1 vccd1
+ _10605_/B sky130_fd_sc_hd__o221a_1
XFILLER_154_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15125_ _15122_/Y _20074_/Q _20463_/Q _15088_/A _15124_/X vssd1 vssd1 vccd1 vccd1
+ _15125_/X sky130_fd_sc_hd__o221a_1
XFILLER_217_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12337_ _12364_/A vssd1 vssd1 vccd1 vccd1 _12376_/A sky130_fd_sc_hd__clkbuf_4
Xoutput108 _17805_/Y vssd1 vssd1 vccd1 vccd1 HRDATA[7] sky130_fd_sc_hd__clkbuf_2
XFILLER_127_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput119 _18112_/Y vssd1 vssd1 vccd1 vccd1 IRQ[1] sky130_fd_sc_hd__clkbuf_2
XFILLER_142_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15056_ _20046_/Q vssd1 vssd1 vccd1 vccd1 _15061_/A sky130_fd_sc_hd__inv_2
X_19933_ _20159_/CLK _19933_/D repeater189/X vssd1 vssd1 vccd1 vccd1 _19933_/Q sky130_fd_sc_hd__dfrtp_1
X_12268_ _20524_/Q vssd1 vssd1 vccd1 vccd1 _12268_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14007_ _20304_/Q _14006_/Y _13988_/A _13881_/B vssd1 vssd1 vccd1 vccd1 _20304_/D
+ sky130_fd_sc_hd__o211a_1
X_11219_ _11225_/A vssd1 vssd1 vccd1 vccd1 _11219_/X sky130_fd_sc_hd__buf_1
X_19864_ _21164_/CLK _19864_/D repeater225/X vssd1 vssd1 vccd1 vccd1 _19864_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_150_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12199_ _20978_/Q _12198_/Y _12109_/X _20336_/Q vssd1 vssd1 vccd1 vccd1 _12199_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_233_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput90 _17329_/Y vssd1 vssd1 vccd1 vccd1 HRDATA[1] sky130_fd_sc_hd__clkbuf_2
XFILLER_228_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18815_ _18814_/X _13928_/Y _18849_/S vssd1 vssd1 vccd1 vccd1 _18815_/X sky130_fd_sc_hd__mux2_1
X_19795_ _19811_/CLK _19795_/D vssd1 vssd1 vccd1 vccd1 _19795_/Q sky130_fd_sc_hd__dfxtp_1
X_18746_ _18745_/X _21281_/Q _18880_/S vssd1 vssd1 vccd1 vccd1 _18746_/X sky130_fd_sc_hd__mux2_2
XANTENNA__13474__A1 _20456_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15958_ _19556_/Q _15954_/X _15891_/X _15956_/X vssd1 vssd1 vccd1 vccd1 _19556_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19285__S0 _19285_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_156_HCLK_A clkbuf_opt_1_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18059__B _18059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14909_ _20567_/Q vssd1 vssd1 vccd1 vccd1 _14909_/Y sky130_fd_sc_hd__inv_2
XFILLER_236_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18677_ _17755_/X _21204_/Q _18928_/S vssd1 vssd1 vccd1 vccd1 _18677_/X sky130_fd_sc_hd__mux2_1
XFILLER_224_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18774__S _18896_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15889_ _15897_/A vssd1 vssd1 vccd1 vccd1 _15889_/X sky130_fd_sc_hd__buf_1
X_17628_ _20174_/Q _17368_/A _14657_/X _17276_/Y _17627_/X vssd1 vssd1 vccd1 vccd1
+ _17628_/X sky130_fd_sc_hd__o221a_1
XFILLER_63_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17898__B _17898_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20735__RESET_B repeater210/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17559_ _16518_/Y _17550_/X _17551_/Y _17376_/X _17558_/X vssd1 vssd1 vccd1 vccd1
+ _17559_/X sky130_fd_sc_hd__o221a_2
XANTENNA__09697__A _15523_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20570_ _20590_/CLK _20570_/D repeater260/X vssd1 vssd1 vccd1 vccd1 _20570_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_220_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19229_ _17517_/Y _17518_/Y _17519_/Y _17520_/Y _20130_/Q _20131_/Q vssd1 vssd1 vccd1
+ vccd1 _19229_/X sky130_fd_sc_hd__mux4_1
XFILLER_192_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15923__B1 _15887_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13012__A _13012_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21122_ _21433_/CLK _21122_/D repeater236/X vssd1 vssd1 vccd1 vccd1 _21122_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18949__S _18962_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19989__RESET_B repeater218/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13162__B1 _12957_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21053_ _21164_/CLK _21053_/D repeater225/X vssd1 vssd1 vccd1 vccd1 _21053_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_99_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20004_ _20004_/CLK _20004_/D repeater225/X vssd1 vssd1 vccd1 vccd1 _20004_/Q sky130_fd_sc_hd__dfstp_1
X_09815_ _09829_/A vssd1 vssd1 vccd1 vccd1 _09815_/X sky130_fd_sc_hd__buf_1
XANTENNA_input3_A HADDR[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09746_ _20145_/Q vssd1 vssd1 vccd1 vccd1 _09746_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19276__S0 _21005_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09677_ _09677_/A vssd1 vssd1 vccd1 vccd1 _15330_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_43_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18684__S _18885_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_15_HCLK_A clkbuf_opt_2_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20906_ _20908_/CLK _20906_/D repeater217/X vssd1 vssd1 vccd1 vccd1 _20906_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_78_HCLK_A clkbuf_4_13_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_3_HCLK_A clkbuf_opt_2_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11228__B1 _10896_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20405__RESET_B repeater184/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20837_ _20930_/CLK _20837_/D repeater257/X vssd1 vssd1 vccd1 vccd1 _20837_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11570_ _15523_/A vssd1 vssd1 vccd1 vccd1 _13171_/A sky130_fd_sc_hd__buf_2
X_20768_ _21319_/CLK _20768_/D repeater191/X vssd1 vssd1 vccd1 vccd1 _20768_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10521_ _10755_/A _20667_/Q _21293_/Q _10517_/Y _10520_/X vssd1 vssd1 vccd1 vccd1
+ _10522_/D sky130_fd_sc_hd__o221a_1
XFILLER_11_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20699_ _21342_/CLK _20699_/D repeater210/X vssd1 vssd1 vccd1 vccd1 _20699_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_7_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13240_ _14258_/A vssd1 vssd1 vccd1 vccd1 _13240_/X sky130_fd_sc_hd__buf_2
XFILLER_182_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10452_ _21279_/Q _10447_/Y _10756_/A _20668_/Q _10451_/X vssd1 vssd1 vccd1 vccd1
+ _10452_/X sky130_fd_sc_hd__a221o_1
XANTENNA__19200__S0 _20130_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_182_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13171_ _13171_/A vssd1 vssd1 vccd1 vccd1 _13171_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_124_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10383_ _10397_/A vssd1 vssd1 vccd1 vccd1 _10383_/X sky130_fd_sc_hd__buf_2
XFILLER_108_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12122_ _20952_/Q vssd1 vssd1 vccd1 vccd1 _12306_/A sky130_fd_sc_hd__inv_2
XANTENNA_input59_A HWDATA[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13153__B1 _13151_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12053_ _20973_/Q _12048_/Y _12326_/A _20387_/Q _12052_/X vssd1 vssd1 vccd1 vccd1
+ _12060_/C sky130_fd_sc_hd__o221a_1
X_16930_ _16930_/A vssd1 vssd1 vccd1 vccd1 _16930_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11004_ _10988_/X _10992_/X _11896_/B vssd1 vssd1 vccd1 vccd1 _11004_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_120_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16861_ _19944_/Q _16861_/B vssd1 vssd1 vccd1 vccd1 _16862_/A sky130_fd_sc_hd__or2_1
XFILLER_238_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18600_ _18848_/A0 _14160_/Y _18902_/S vssd1 vssd1 vccd1 vccd1 _18600_/X sky130_fd_sc_hd__mux2_1
X_15812_ _16163_/A vssd1 vssd1 vccd1 vccd1 _15812_/X sky130_fd_sc_hd__clkbuf_2
X_19580_ _21040_/CLK _19580_/D vssd1 vssd1 vccd1 vccd1 _19580_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__19267__S0 _20130_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16792_ _16795_/B _16791_/Y _16779_/X vssd1 vssd1 vccd1 vccd1 _16792_/X sky130_fd_sc_hd__o21a_1
XFILLER_218_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18531_ _18530_/X _21361_/Q _18850_/S vssd1 vssd1 vccd1 vccd1 _18531_/X sky130_fd_sc_hd__mux2_1
XFILLER_246_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15743_ _15750_/A vssd1 vssd1 vccd1 vccd1 _15743_/X sky130_fd_sc_hd__buf_1
XFILLER_93_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12955_ _20709_/Q _12948_/X _12954_/X _12951_/X vssd1 vssd1 vccd1 vccd1 _20709_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18594__S _18884_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_233_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11906_ _11906_/A vssd1 vssd1 vccd1 vccd1 _11906_/Y sky130_fd_sc_hd__inv_2
X_18462_ _18461_/X _10584_/Y _18775_/S vssd1 vssd1 vccd1 vccd1 _18462_/X sky130_fd_sc_hd__mux2_1
XFILLER_73_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15674_ _15681_/A vssd1 vssd1 vccd1 vccd1 _15674_/X sky130_fd_sc_hd__buf_1
X_12886_ _13104_/B vssd1 vssd1 vccd1 vccd1 _17178_/A sky130_fd_sc_hd__clkbuf_2
XPHY_4360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17413_ _19393_/Q vssd1 vssd1 vccd1 vccd1 _17413_/Y sky130_fd_sc_hd__inv_2
XPHY_4393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14625_ _20193_/Q _14623_/Y _14624_/X _14583_/B vssd1 vssd1 vccd1 vccd1 _20193_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__20146__RESET_B repeater250/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11837_ _11837_/A vssd1 vssd1 vccd1 vccd1 _11838_/B sky130_fd_sc_hd__inv_2
XFILLER_33_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18393_ _18848_/A0 _14116_/Y _18902_/S vssd1 vssd1 vccd1 vccd1 _18393_/X sky130_fd_sc_hd__mux2_1
XPHY_3670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14556_ _20137_/Q vssd1 vssd1 vccd1 vccd1 _15799_/A sky130_fd_sc_hd__buf_1
X_17344_ _19294_/Q vssd1 vssd1 vccd1 vccd1 _17344_/Y sky130_fd_sc_hd__inv_2
X_11768_ _19085_/X _11764_/X _21049_/Q _11765_/X vssd1 vssd1 vccd1 vccd1 _21049_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_60_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10719_ _21315_/Q _10718_/Y _10704_/B _10712_/X vssd1 vssd1 vccd1 vccd1 _21315_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13507_ _13515_/A vssd1 vssd1 vccd1 vccd1 _13507_/X sky130_fd_sc_hd__buf_1
X_14487_ _20226_/Q _14486_/Y _14370_/B _14477_/X vssd1 vssd1 vccd1 vccd1 _20226_/D
+ sky130_fd_sc_hd__o211a_1
X_17275_ _20140_/Q vssd1 vssd1 vccd1 vccd1 _17275_/Y sky130_fd_sc_hd__inv_2
X_11699_ _11705_/A vssd1 vssd1 vccd1 vccd1 _11699_/X sky130_fd_sc_hd__buf_1
XFILLER_228_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19014_ _16935_/Y _20409_/Q _19019_/S vssd1 vssd1 vccd1 vccd1 _19962_/D sky130_fd_sc_hd__mux2_1
X_13438_ _20472_/Q _13436_/X _13240_/X _13437_/X vssd1 vssd1 vccd1 vccd1 _20472_/D
+ sky130_fd_sc_hd__a22o_1
X_16226_ _19424_/Q _16223_/X _16123_/X _16224_/X vssd1 vssd1 vccd1 vccd1 _19424_/D
+ sky130_fd_sc_hd__a22o_1
Xrebuffer1 _20027_/Q vssd1 vssd1 vccd1 vccd1 _15331_/A1 sky130_fd_sc_hd__dlygate4sd1_1
X_16157_ _19458_/Q _16151_/X _16139_/X _16153_/X vssd1 vssd1 vccd1 vccd1 _19458_/D
+ sky130_fd_sc_hd__a22o_1
X_13369_ _20507_/Q _13365_/X _13311_/X _13366_/X vssd1 vssd1 vccd1 vccd1 _20507_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_182_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15108_ _15103_/Y _20073_/Q _20440_/Q _15066_/A vssd1 vssd1 vccd1 vccd1 _15108_/X
+ sky130_fd_sc_hd__o22a_1
X_16088_ _16088_/A vssd1 vssd1 vccd1 vccd1 _16088_/X sky130_fd_sc_hd__buf_1
XANTENNA__16330__B1 _16235_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18769__S _18879_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19916_ _21196_/CLK _19916_/D repeater220/X vssd1 vssd1 vccd1 vccd1 _19916_/Q sky130_fd_sc_hd__dfrtp_1
X_15039_ _20063_/Q vssd1 vssd1 vccd1 vccd1 _15077_/A sky130_fd_sc_hd__inv_2
XFILLER_170_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19847_ _20042_/CLK _19847_/D repeater219/X vssd1 vssd1 vccd1 vccd1 _19847_/Q sky130_fd_sc_hd__dfrtp_1
X_09600_ _20888_/Q _09937_/B _10973_/C vssd1 vssd1 vccd1 vccd1 _14303_/C sky130_fd_sc_hd__or3_4
XFILLER_68_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20916__RESET_B repeater218/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19258__S0 _20130_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19778_ _21222_/CLK _19778_/D vssd1 vssd1 vccd1 vccd1 _19778_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_243_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11458__B1 _21071_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18729_ _18728_/X _12180_/Y _18787_/S vssd1 vssd1 vccd1 vccd1 _18729_/X sky130_fd_sc_hd__mux2_2
XFILLER_243_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_236_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13007__A _13013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16397__B1 _16237_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12958__B1 _12957_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20622_ _20622_/CLK _20622_/D repeater195/X vssd1 vssd1 vccd1 vccd1 _20622_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15222__A _20481_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16149__B1 _15916_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17140__C _17838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20553_ _20947_/CLK _20553_/D repeater266/X vssd1 vssd1 vccd1 vccd1 _20553_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_137_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20484_ _20944_/CLK _20484_/D repeater274/X vssd1 vssd1 vccd1 vccd1 _20484_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_164_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17149__A _17553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16321__B1 _16009_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18679__S _18835_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13135__B1 _12928_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21105_ _21424_/CLK _21105_/D repeater231/X vssd1 vssd1 vccd1 vccd1 _21105_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_78_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21036_ _21207_/CLK _21036_/D repeater242/X vssd1 vssd1 vccd1 vccd1 _21036_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_59_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19249__S0 _20130_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_228_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09729_ _09724_/Y _20159_/Q _21239_/Q _09725_/Y _09728_/X vssd1 vssd1 vccd1 vccd1
+ _09769_/B sky130_fd_sc_hd__o221a_1
XFILLER_28_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12740_ _14686_/A _12740_/B vssd1 vssd1 vccd1 vccd1 _14674_/A sky130_fd_sc_hd__or2_2
XFILLER_216_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17585__C1 _17584_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_231_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12671_ _20835_/Q _12662_/X _12670_/X _12664_/X vssd1 vssd1 vccd1 vccd1 _20835_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14410_ _20236_/Q vssd1 vssd1 vccd1 vccd1 _14410_/Y sky130_fd_sc_hd__inv_2
XPHY_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11622_ _14813_/B _11625_/B _11617_/X vssd1 vssd1 vccd1 vccd1 _21109_/D sky130_fd_sc_hd__a21o_1
XPHY_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15390_ _15390_/A vssd1 vssd1 vccd1 vccd1 _15390_/X sky130_fd_sc_hd__buf_1
XPHY_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14341_ _20224_/Q vssd1 vssd1 vccd1 vccd1 _14462_/A sky130_fd_sc_hd__inv_2
XPHY_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11553_ _11562_/A vssd1 vssd1 vccd1 vccd1 _11566_/A sky130_fd_sc_hd__inv_2
XPHY_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17888__B1 _18415_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10504_ _21286_/Q vssd1 vssd1 vccd1 vccd1 _10763_/B sky130_fd_sc_hd__inv_2
XPHY_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17060_ _17060_/A _17060_/B _17060_/C vssd1 vssd1 vccd1 vccd1 _18912_/S sky130_fd_sc_hd__and3_1
XPHY_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14272_ _20244_/Q _14267_/X _13714_/X _14268_/X vssd1 vssd1 vccd1 vccd1 _20244_/D
+ sky130_fd_sc_hd__a22o_1
X_11484_ _19105_/X _11480_/X _21153_/Q _11481_/X vssd1 vssd1 vccd1 vccd1 _21153_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_171_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16011_ _19529_/Q _16008_/X _16009_/X _16010_/X vssd1 vssd1 vccd1 vccd1 _19529_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_7_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13223_ input45/X vssd1 vssd1 vccd1 vccd1 _13223_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__13374__B1 _13243_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10435_ _20680_/Q vssd1 vssd1 vccd1 vccd1 _17900_/A sky130_fd_sc_hd__inv_2
XFILLER_109_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13154_ input39/X vssd1 vssd1 vccd1 vccd1 _13154_/X sky130_fd_sc_hd__buf_2
XFILLER_88_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10366_ _10366_/A vssd1 vssd1 vccd1 vccd1 _10397_/A sky130_fd_sc_hd__buf_1
XANTENNA__18589__S _18787_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12105_ _12323_/A vssd1 vssd1 vccd1 vccd1 _12105_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_69_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17962_ _18527_/X _17926_/X _18520_/X _17927_/X _17961_/X vssd1 vssd1 vccd1 vccd1
+ _17966_/B sky130_fd_sc_hd__o221a_2
XFILLER_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13085_ _20646_/Q _13079_/X _12857_/X _13081_/X vssd1 vssd1 vccd1 vccd1 _20646_/D
+ sky130_fd_sc_hd__a22o_1
X_10297_ _21363_/Q _10296_/Y _10273_/A _20717_/Q vssd1 vssd1 vccd1 vccd1 _10297_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_239_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19701_ _20432_/CLK _19701_/D vssd1 vssd1 vccd1 vccd1 _19701_/Q sky130_fd_sc_hd__dfxtp_1
X_16913_ _16913_/A vssd1 vssd1 vccd1 vccd1 _16913_/Y sky130_fd_sc_hd__inv_2
X_12036_ _12317_/A vssd1 vssd1 vccd1 vccd1 _12036_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_104_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17893_ _18079_/A vssd1 vssd1 vccd1 vccd1 _17974_/A sky130_fd_sc_hd__buf_1
XFILLER_120_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19632_ _19821_/CLK _19632_/D vssd1 vssd1 vccd1 vccd1 _19632_/Q sky130_fd_sc_hd__dfxtp_1
X_16844_ _16844_/A vssd1 vssd1 vccd1 vccd1 _16844_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20398__RESET_B repeater270/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_225_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19563_ _19812_/CLK _19563_/D vssd1 vssd1 vccd1 vccd1 _19563_/Q sky130_fd_sc_hd__dfxtp_1
X_16775_ _16778_/B _16774_/Y _16762_/X vssd1 vssd1 vccd1 vccd1 _16775_/X sky130_fd_sc_hd__o21a_1
XANTENNA__20327__RESET_B repeater235/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_225_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13987_ _13987_/A vssd1 vssd1 vccd1 vccd1 _13988_/A sky130_fd_sc_hd__buf_1
XFILLER_218_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_230_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18514_ _18513_/X _13935_/Y _18849_/S vssd1 vssd1 vccd1 vccd1 _18514_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15726_ _15736_/A vssd1 vssd1 vccd1 vccd1 _15737_/A sky130_fd_sc_hd__inv_2
X_19494_ _20326_/CLK _19494_/D vssd1 vssd1 vccd1 vccd1 _19494_/Q sky130_fd_sc_hd__dfxtp_1
X_12938_ _20718_/Q _12935_/X _12849_/X _12937_/X vssd1 vssd1 vccd1 vccd1 _20718_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_33_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_233_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18445_ _17902_/Y _16805_/Y _18875_/S vssd1 vssd1 vccd1 vccd1 _18445_/X sky130_fd_sc_hd__mux2_1
X_15657_ _15657_/A vssd1 vssd1 vccd1 vccd1 _15657_/X sky130_fd_sc_hd__buf_1
XPHY_4190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_61_HCLK_A clkbuf_4_14_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12869_ _20745_/Q _12867_/X _12544_/X _12868_/X vssd1 vssd1 vccd1 vccd1 _20745_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12666__A input56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11570__A _15523_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14608_ _14591_/A _14591_/B _14607_/X _14605_/Y vssd1 vssd1 vccd1 vccd1 _20202_/D
+ sky130_fd_sc_hd__a211oi_2
X_18376_ _18375_/X _20196_/Q _18748_/S vssd1 vssd1 vccd1 vccd1 _18376_/X sky130_fd_sc_hd__mux2_2
X_15588_ _15588_/A vssd1 vssd1 vccd1 vccd1 _15588_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__17328__C1 _17322_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_92_HCLK clkbuf_4_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _21375_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_193_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17327_ _18838_/X _17324_/X _18847_/X _17326_/X vssd1 vssd1 vccd1 vccd1 _17327_/X
+ sky130_fd_sc_hd__o22a_1
X_14539_ _15815_/A _15832_/B vssd1 vssd1 vccd1 vccd1 _15902_/B sky130_fd_sc_hd__or2_2
XFILLER_239_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20504__CLK _20930_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17258_ _19447_/Q vssd1 vssd1 vccd1 vccd1 _17258_/Y sky130_fd_sc_hd__inv_2
XFILLER_128_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21115__RESET_B repeater233/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16209_ _19433_/Q _16206_/X _16207_/X _16208_/X vssd1 vssd1 vccd1 vccd1 _19433_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19677__CLK _19813_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17189_ _21309_/Q vssd1 vssd1 vccd1 vccd1 _17189_/Y sky130_fd_sc_hd__inv_2
XFILLER_161_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15106__B2 _15099_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18499__S _18908_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13117__B1 _12989_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18056__B1 _18267_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17803__B1 _18141_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20750__RESET_B repeater210/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20068__RESET_B repeater276/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_225_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18962__S _18962_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20605_ _20622_/CLK _20605_/D repeater195/X vssd1 vssd1 vccd1 vccd1 _20605_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_rebuffer1_A _20027_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15887__A _16231_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14791__A _20119_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20536_ _20947_/CLK _20536_/D repeater267/X vssd1 vssd1 vccd1 vccd1 _20536_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_181_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20467_ _20937_/CLK _20467_/D repeater277/X vssd1 vssd1 vccd1 vccd1 _20467_/Q sky130_fd_sc_hd__dfrtp_1
X_10220_ _10220_/A vssd1 vssd1 vccd1 vccd1 _10221_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_3_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20398_ _21234_/CLK _20398_/D repeater270/X vssd1 vssd1 vccd1 vccd1 _20398_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10151_ _10151_/A _10151_/B vssd1 vssd1 vccd1 vccd1 _10193_/A sky130_fd_sc_hd__or2_1
XFILLER_134_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20838__RESET_B repeater257/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18202__S _18884_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18047__B1 _18264_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10082_ _20798_/Q vssd1 vssd1 vccd1 vccd1 _10082_/Y sky130_fd_sc_hd__inv_2
XFILLER_121_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21019_ _21021_/CLK _21019_/D repeater238/X vssd1 vssd1 vccd1 vccd1 _21019_/Q sky130_fd_sc_hd__dfrtp_2
X_13910_ _13907_/Y _20291_/Q _20634_/Q _14009_/A _13909_/X vssd1 vssd1 vccd1 vccd1
+ _13914_/C sky130_fd_sc_hd__o221a_1
XFILLER_247_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14890_ _14889_/Y _20102_/Q _20569_/Q _15000_/A vssd1 vssd1 vccd1 vccd1 _14894_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09770__D _14309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20420__RESET_B repeater187/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13841_ _20321_/Q vssd1 vssd1 vccd1 vccd1 _13897_/A sky130_fd_sc_hd__inv_2
XFILLER_235_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19033__S _19046_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16560_ _16564_/A vssd1 vssd1 vccd1 vccd1 _16744_/A sky130_fd_sc_hd__buf_1
X_13772_ _13770_/Y _20202_/Q _20610_/Q _14576_/A vssd1 vssd1 vccd1 vccd1 _13772_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_15_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10984_ _21245_/Q vssd1 vssd1 vccd1 vccd1 _10985_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_74_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15511_ _19764_/Q _15507_/X _15454_/X _15509_/X vssd1 vssd1 vccd1 vccd1 _19764_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_215_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12723_ _13535_/B _13106_/B vssd1 vssd1 vccd1 vccd1 _12724_/S sky130_fd_sc_hd__or2_1
XANTENNA__18872__S _18910_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16491_ _16526_/B vssd1 vssd1 vccd1 vccd1 _16491_/Y sky130_fd_sc_hd__inv_2
XFILLER_203_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18230_ _20854_/Q input3/X _18236_/S vssd1 vssd1 vccd1 vccd1 _18230_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15442_ _15442_/A vssd1 vssd1 vccd1 vccd1 _15442_/X sky130_fd_sc_hd__buf_1
X_12654_ _12680_/A vssd1 vssd1 vccd1 vccd1 _12654_/X sky130_fd_sc_hd__buf_1
XFILLER_231_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11605_ _11605_/A vssd1 vssd1 vccd1 vccd1 _11605_/X sky130_fd_sc_hd__buf_1
X_18161_ _18004_/Y _21485_/Q _18669_/S vssd1 vssd1 vccd1 vccd1 _18161_/X sky130_fd_sc_hd__mux2_1
XPHY_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15797__A _15832_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12585_ _20883_/Q _12581_/X _18235_/X _12583_/X vssd1 vssd1 vccd1 vccd1 _20883_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15373_ _15505_/C vssd1 vssd1 vccd1 vccd1 _16594_/B sky130_fd_sc_hd__buf_1
XFILLER_196_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17112_ _17773_/B vssd1 vssd1 vccd1 vccd1 _17369_/B sky130_fd_sc_hd__clkbuf_2
X_11536_ _21139_/Q _11534_/X _10894_/X _11535_/X vssd1 vssd1 vccd1 vccd1 _21139_/D
+ sky130_fd_sc_hd__a22o_1
X_14324_ _14324_/A _14324_/B _14324_/C _14324_/D vssd1 vssd1 vccd1 vccd1 _14324_/X
+ sky130_fd_sc_hd__or4_4
XPHY_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18092_ _20427_/Q vssd1 vssd1 vccd1 vccd1 _18092_/Y sky130_fd_sc_hd__inv_2
XFILLER_183_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13347__B1 _13287_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14255_ _20251_/Q vssd1 vssd1 vccd1 vccd1 _16720_/A sky130_fd_sc_hd__buf_2
XFILLER_116_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17043_ _21409_/Q vssd1 vssd1 vccd1 vccd1 _17043_/Y sky130_fd_sc_hd__inv_2
X_11467_ _19094_/X _11461_/X _21164_/Q _11463_/X vssd1 vssd1 vccd1 vccd1 _21164_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_109_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13110__A _13110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13206_ _13215_/A vssd1 vssd1 vccd1 vccd1 _13206_/X sky130_fd_sc_hd__buf_1
X_10418_ _10418_/A vssd1 vssd1 vccd1 vccd1 _10418_/Y sky130_fd_sc_hd__inv_2
X_14186_ _14095_/A _14095_/B _14185_/X _14182_/Y vssd1 vssd1 vccd1 vccd1 _20285_/D
+ sky130_fd_sc_hd__a211oi_2
X_11398_ _11342_/A _11395_/Y _11396_/X vssd1 vssd1 vccd1 vccd1 _11418_/A sky130_fd_sc_hd__o21ai_2
XFILLER_124_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13137_ _20615_/Q _13132_/X _12932_/X _13133_/X vssd1 vssd1 vccd1 vccd1 _20615_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_225_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10349_ _21345_/Q _10347_/Y _21371_/Q _10348_/Y vssd1 vssd1 vccd1 vccd1 _10349_/X
+ sky130_fd_sc_hd__o22a_1
X_18994_ _17027_/Y _11022_/B _20005_/Q vssd1 vssd1 vccd1 vccd1 _20005_/D sky130_fd_sc_hd__mux2_1
XFILLER_239_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17945_ _18085_/B vssd1 vssd1 vccd1 vccd1 _18007_/B sky130_fd_sc_hd__clkbuf_2
X_13068_ _20657_/Q _13066_/X _13006_/X _13067_/X vssd1 vssd1 vccd1 vccd1 _20657_/D
+ sky130_fd_sc_hd__a22o_1
Xrepeater205 repeater206/X vssd1 vssd1 vccd1 vccd1 repeater205/X sky130_fd_sc_hd__buf_6
XFILLER_239_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater216 repeater219/X vssd1 vssd1 vccd1 vccd1 repeater216/X sky130_fd_sc_hd__buf_8
X_12019_ _19071_/X _12017_/X _20994_/Q _12018_/X vssd1 vssd1 vccd1 vccd1 _20994_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11565__A _13166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater227 repeater228/X vssd1 vssd1 vccd1 vccd1 repeater227/X sky130_fd_sc_hd__buf_8
X_17876_ _20823_/Q vssd1 vssd1 vccd1 vccd1 _17876_/Y sky130_fd_sc_hd__inv_2
Xrepeater238 repeater241/X vssd1 vssd1 vccd1 vccd1 repeater238/X sky130_fd_sc_hd__buf_8
XFILLER_241_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater249 repeater250/X vssd1 vssd1 vccd1 vccd1 repeater249/X sky130_fd_sc_hd__buf_8
XFILLER_93_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19615_ _20137_/CLK _19615_/D vssd1 vssd1 vccd1 vccd1 _19615_/Q sky130_fd_sc_hd__dfxtp_1
X_16827_ _19937_/Q _16827_/B vssd1 vssd1 vccd1 vccd1 _16843_/B sky130_fd_sc_hd__or2_1
XFILLER_207_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19546_ _19789_/CLK _19546_/D vssd1 vssd1 vccd1 vccd1 _19546_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_opt_6_HCLK_A clkbuf_opt_7_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16758_ _16758_/A _16758_/B vssd1 vssd1 vccd1 vccd1 _16758_/Y sky130_fd_sc_hd__nor2_1
XFILLER_53_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18210__A0 _18209_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15709_ _15716_/A vssd1 vssd1 vccd1 vccd1 _15709_/X sky130_fd_sc_hd__clkbuf_2
X_19477_ _20432_/CLK _19477_/D vssd1 vssd1 vccd1 vccd1 _19477_/Q sky130_fd_sc_hd__dfxtp_1
X_16689_ _16689_/A _16689_/B _16689_/C vssd1 vssd1 vccd1 vccd1 _19881_/D sky130_fd_sc_hd__and3_1
XANTENNA__18782__S _18850_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18761__A1 _19231_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18428_ _18427_/X _16933_/Y _18680_/S vssd1 vssd1 vccd1 vccd1 _18428_/X sky130_fd_sc_hd__mux2_2
XANTENNA__21367__RESET_B repeater254/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21452__CLK _21452_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18359_ _18358_/X _16999_/A _18875_/S vssd1 vssd1 vccd1 vccd1 _18359_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15327__A1 _20029_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21370_ _21374_/CLK _21370_/D repeater255/X vssd1 vssd1 vccd1 vccd1 _21370_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_190_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13338__B1 _13274_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20321_ _20665_/CLK _20321_/D repeater261/X vssd1 vssd1 vccd1 vccd1 _20321_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_147_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11459__B _19870_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20252_ _21055_/CLK _20252_/D repeater221/X vssd1 vssd1 vccd1 vccd1 _20252_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_115_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20183_ _21480_/CLK _20183_/D repeater206/X vssd1 vssd1 vccd1 vccd1 _20183_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_170_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09994_ _20023_/Q vssd1 vssd1 vccd1 vccd1 _09994_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18957__S _18962_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13510__B1 _13509_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_229_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20003__D _20003_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18692__S _18902_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19842__CLK _21134_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13577__B1 _13422_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21037__RESET_B repeater242/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12370_ _20963_/Q _12369_/Y _12359_/X _12317_/B vssd1 vssd1 vccd1 vccd1 _20963_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_165_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11321_ _16587_/A vssd1 vssd1 vccd1 vccd1 _16564_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_181_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20519_ _20943_/CLK _20519_/D repeater275/X vssd1 vssd1 vccd1 vccd1 _20519_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_176_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14040_ _20288_/Q vssd1 vssd1 vccd1 vccd1 _14098_/A sky130_fd_sc_hd__inv_2
X_11252_ _19063_/X _11250_/X _21189_/Q _11251_/X vssd1 vssd1 vccd1 vccd1 _21189_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_4_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10203_ _10203_/A _10203_/B vssd1 vssd1 vccd1 vccd1 _10213_/A sky130_fd_sc_hd__or2_1
XFILLER_69_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19028__S _19058_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11183_ _15884_/A vssd1 vssd1 vccd1 vccd1 _15847_/A sky130_fd_sc_hd__buf_1
XFILLER_192_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input41_A HWDATA[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10134_ _21399_/Q _10133_/Y _10160_/A _20796_/Q vssd1 vssd1 vccd1 vccd1 _10134_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15991_ _19539_/Q _15986_/X _15975_/X _15988_/X vssd1 vssd1 vccd1 vccd1 _19539_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_192_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18867__S _18927_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13501__B1 _13429_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17730_ _18706_/X _17216_/A _18680_/X _17223_/A vssd1 vssd1 vccd1 vccd1 _17730_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_48_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14942_ _20570_/Q vssd1 vssd1 vccd1 vccd1 _14942_/Y sky130_fd_sc_hd__inv_2
X_10065_ _21395_/Q vssd1 vssd1 vccd1 vccd1 _10156_/A sky130_fd_sc_hd__inv_2
XFILLER_48_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17661_ _18724_/X _17839_/A _18727_/X _17319_/X _17660_/X vssd1 vssd1 vccd1 vccd1
+ _17661_/X sky130_fd_sc_hd__o221a_2
X_14873_ _14961_/C _14984_/A vssd1 vssd1 vccd1 vccd1 _14874_/B sky130_fd_sc_hd__or2_2
XFILLER_91_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output128_A _21120_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19400_ _19812_/CLK _19400_/D vssd1 vssd1 vccd1 vccd1 _19400_/Q sky130_fd_sc_hd__dfxtp_1
X_16612_ _16537_/Y _16611_/X _16610_/Y _16604_/X _16564_/X vssd1 vssd1 vccd1 vccd1
+ _19987_/D sky130_fd_sc_hd__o221ai_1
X_13824_ _20605_/Q vssd1 vssd1 vccd1 vccd1 _13824_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12607__A2 _12600_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17592_ _19363_/Q vssd1 vssd1 vccd1 vccd1 _17592_/Y sky130_fd_sc_hd__inv_2
XFILLER_141_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19331_ _19834_/CLK _19331_/D vssd1 vssd1 vccd1 vccd1 _19331_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_216_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16543_ _16740_/A _16535_/X _16737_/A _16542_/Y vssd1 vssd1 vccd1 vccd1 _19993_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_189_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13755_ _20606_/Q vssd1 vssd1 vccd1 vccd1 _13755_/Y sky130_fd_sc_hd__inv_2
X_10967_ _10965_/Y _10966_/Y _21212_/Q _21039_/Q vssd1 vssd1 vccd1 vccd1 _10967_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_231_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18743__A1 _20777_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12706_ _20815_/Q _12701_/X _11733_/X _12702_/X vssd1 vssd1 vccd1 vccd1 _20815_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__21460__RESET_B repeater245/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19262_ _17236_/Y _17237_/Y _17238_/Y _17239_/Y _19275_/S0 _21004_/Q vssd1 vssd1
+ vccd1 vccd1 _19262_/X sky130_fd_sc_hd__mux4_2
XFILLER_31_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16474_ _16474_/A vssd1 vssd1 vccd1 vccd1 _16474_/X sky130_fd_sc_hd__buf_1
XANTENNA__16754__B1 _16835_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13686_ _13706_/A vssd1 vssd1 vccd1 vccd1 _13686_/X sky130_fd_sc_hd__buf_1
X_10898_ _10898_/A vssd1 vssd1 vccd1 vccd1 _10898_/X sky130_fd_sc_hd__buf_2
XFILLER_70_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18213_ _18212_/X _14586_/A _18748_/S vssd1 vssd1 vccd1 vccd1 _18213_/X sky130_fd_sc_hd__mux2_1
X_15425_ _15425_/A vssd1 vssd1 vccd1 vccd1 _15425_/X sky130_fd_sc_hd__buf_1
X_19193_ _19548_/Q _19540_/Q _19532_/Q _19516_/Q _19280_/S0 _20122_/Q vssd1 vssd1
+ vccd1 vccd1 _19193_/X sky130_fd_sc_hd__mux4_2
X_12637_ _12637_/A vssd1 vssd1 vccd1 vccd1 _12637_/X sky130_fd_sc_hd__buf_1
XPHY_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18144_ _18143_/X _13832_/Y _18748_/S vssd1 vssd1 vccd1 vccd1 _18144_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12568_ _12580_/A vssd1 vssd1 vccd1 vccd1 _12582_/A sky130_fd_sc_hd__inv_2
X_15356_ _19830_/Q _15345_/X _15355_/X _15347_/X vssd1 vssd1 vccd1 vccd1 _19830_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_8_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11519_ _21145_/Q vssd1 vssd1 vccd1 vccd1 _17064_/A sky130_fd_sc_hd__inv_2
XFILLER_145_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14307_ _21442_/Q _14307_/B _14307_/C vssd1 vssd1 vccd1 vccd1 _14308_/A sky130_fd_sc_hd__and3_1
XFILLER_7_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18075_ _18130_/X _17219_/X _18660_/X _18064_/X _18074_/X vssd1 vssd1 vccd1 vccd1
+ _18076_/C sky130_fd_sc_hd__o221a_1
X_12499_ _16587_/A vssd1 vssd1 vccd1 vccd1 _16609_/A sky130_fd_sc_hd__buf_1
X_15287_ _19852_/Q _19853_/Q vssd1 vssd1 vccd1 vccd1 _15288_/B sky130_fd_sc_hd__or2_1
XFILLER_236_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18259__A0 _17079_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17026_ _17026_/A _17026_/B vssd1 vssd1 vccd1 vccd1 _20012_/D sky130_fd_sc_hd__nor2_1
X_14238_ _19898_/Q _14238_/B vssd1 vssd1 vccd1 vccd1 _14239_/B sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_122_HCLK clkbuf_opt_3_HCLK/A vssd1 vssd1 vccd1 vccd1 _20971_/CLK sky130_fd_sc_hd__clkbuf_16
X_14169_ _14167_/Y _20260_/Q _20546_/Q _14085_/A _14168_/X vssd1 vssd1 vccd1 vccd1
+ _14170_/D sky130_fd_sc_hd__o221a_1
XFILLER_124_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19715__CLK _21009_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17482__A1 _17060_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18977_ _21429_/Q _21102_/Q _18983_/S vssd1 vssd1 vccd1 vccd1 _18977_/X sky130_fd_sc_hd__mux2_1
XANTENNA__18777__S _18896_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17928_ _17928_/A vssd1 vssd1 vccd1 vccd1 _17928_/X sky130_fd_sc_hd__buf_1
XFILLER_239_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17859_ _18596_/X _17857_/X _18587_/X _17858_/X vssd1 vssd1 vccd1 vccd1 _17859_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_242_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20870_ _21431_/CLK _20870_/D repeater238/X vssd1 vssd1 vccd1 vccd1 _20870_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_242_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19529_ _19784_/CLK _19529_/D vssd1 vssd1 vccd1 vccd1 _19529_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_207_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21422_ _21424_/CLK _21422_/D repeater231/X vssd1 vssd1 vccd1 vccd1 _21422_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18498__A0 _18497_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21353_ _21368_/CLK _21353_/D repeater255/X vssd1 vssd1 vccd1 vccd1 _21353_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_162_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20304_ _20693_/CLK _20304_/D repeater196/X vssd1 vssd1 vccd1 vccd1 _20304_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__11189__B _11549_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21284_ _21306_/CLK _21284_/D repeater207/X vssd1 vssd1 vccd1 vccd1 _21284_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__15884__B _17153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20235_ _21477_/CLK _20235_/D repeater203/X vssd1 vssd1 vccd1 vccd1 _20235_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17157__A _17169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20166_ _21011_/CLK _20166_/D repeater237/X vssd1 vssd1 vccd1 vccd1 _20166_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18687__S _18775_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09977_ _21417_/Q _09975_/X _09682_/X _09976_/X vssd1 vssd1 vccd1 vccd1 _21417_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_103_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20097_ _20101_/CLK _20097_/D repeater259/X vssd1 vssd1 vccd1 vccd1 _20097_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_29_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11870_ _11180_/X _10964_/X _11822_/B _11869_/X vssd1 vssd1 vccd1 vccd1 _21026_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_169_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13798__B1 _20602_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10821_ _10821_/A vssd1 vssd1 vccd1 vccd1 _10824_/B sky130_fd_sc_hd__inv_2
XFILLER_232_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__21218__RESET_B repeater242/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20999_ _21223_/CLK _20999_/D repeater241/X vssd1 vssd1 vccd1 vccd1 _20999_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_41_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13540_ _13574_/A vssd1 vssd1 vccd1 vccd1 _13567_/A sky130_fd_sc_hd__clkbuf_2
X_10752_ _19289_/Q _10752_/B vssd1 vssd1 vccd1 vccd1 _10752_/X sky130_fd_sc_hd__and2_1
XFILLER_186_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13471_ _20457_/Q _13466_/X _13284_/X _13467_/X vssd1 vssd1 vccd1 vccd1 _20457_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10683_ _10683_/A vssd1 vssd1 vccd1 vccd1 _10683_/Y sky130_fd_sc_hd__inv_2
XFILLER_197_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15210_ _15128_/X _15063_/B _15208_/Y _15179_/A vssd1 vssd1 vccd1 vccd1 _20048_/D
+ sky130_fd_sc_hd__a211oi_2
X_12422_ _12422_/A _12461_/A vssd1 vssd1 vccd1 vccd1 _12423_/B sky130_fd_sc_hd__or2_2
XANTENNA__18489__A0 _18488_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16190_ _19440_/Q _16187_/X _16145_/X _16188_/X vssd1 vssd1 vccd1 vccd1 _19440_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_127_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_145_HCLK clkbuf_opt_1_HCLK/A vssd1 vssd1 vccd1 vccd1 _20172_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_127_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12353_ _20973_/Q _12352_/Y _12344_/X _12327_/B vssd1 vssd1 vccd1 vccd1 _20973_/D
+ sky130_fd_sc_hd__o211a_1
X_15141_ _20448_/Q vssd1 vssd1 vccd1 vccd1 _15141_/Y sky130_fd_sc_hd__inv_2
XFILLER_139_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20853__RESET_B repeater243/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11304_ _11315_/C _11315_/A _20915_/Q _11304_/D vssd1 vssd1 vccd1 vccd1 _12502_/B
+ sky130_fd_sc_hd__and4b_1
XFILLER_153_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15072_ _15099_/A _15072_/B vssd1 vssd1 vccd1 vccd1 _15191_/A sky130_fd_sc_hd__or2_1
XANTENNA__19738__CLK _19765_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12284_ _20516_/Q vssd1 vssd1 vccd1 vccd1 _12284_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18900_ _18899_/X _14824_/Y _18910_/S vssd1 vssd1 vccd1 vccd1 _18900_/X sky130_fd_sc_hd__mux2_1
X_14023_ _14023_/A vssd1 vssd1 vccd1 vccd1 _14023_/Y sky130_fd_sc_hd__inv_2
X_11235_ _11235_/A vssd1 vssd1 vccd1 vccd1 _11235_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13595__A _13595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19880_ _21147_/CLK _19880_/D repeater212/X vssd1 vssd1 vccd1 vccd1 _19880_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_96_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18831_ _18830_/X _17346_/Y _18927_/S vssd1 vssd1 vccd1 vccd1 _18831_/X sky130_fd_sc_hd__mux2_1
XFILLER_122_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11166_ _11123_/Y _11151_/X _11138_/Y _11165_/X vssd1 vssd1 vccd1 vccd1 _21223_/D
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__18597__S _18884_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10117_ _10059_/A _20793_/Q _10071_/A _20795_/Q vssd1 vssd1 vccd1 vccd1 _10117_/Y
+ sky130_fd_sc_hd__a22oi_1
X_18762_ _17508_/Y _17507_/Y _18926_/S vssd1 vssd1 vccd1 vccd1 _18762_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12004__A _21185_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15974_ _19548_/Q _15968_/X _15973_/X _15971_/X vssd1 vssd1 vccd1 vccd1 _19548_/D
+ sky130_fd_sc_hd__a22o_1
X_11097_ _11093_/B _11066_/B _11096_/X _11050_/A _11096_/A vssd1 vssd1 vccd1 vccd1
+ _21231_/D sky130_fd_sc_hd__a32o_1
XFILLER_95_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17713_ _19845_/Q vssd1 vssd1 vccd1 vccd1 _17713_/Y sky130_fd_sc_hd__inv_2
X_14925_ _14897_/Y _20077_/Q _14922_/Y _20099_/Q _14924_/X vssd1 vssd1 vccd1 vccd1
+ _14933_/B sky130_fd_sc_hd__o221a_1
X_10048_ _21384_/Q vssd1 vssd1 vccd1 vccd1 _10049_/A sky130_fd_sc_hd__inv_2
X_18693_ _18692_/X _13939_/Y _18849_/S vssd1 vssd1 vccd1 vccd1 _18693_/X sky130_fd_sc_hd__mux2_1
XFILLER_236_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17644_ _16512_/Y _17550_/A _17643_/Y _17295_/X vssd1 vssd1 vccd1 vccd1 _17644_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_75_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14856_ _20081_/Q vssd1 vssd1 vccd1 vccd1 _15001_/A sky130_fd_sc_hd__inv_2
XFILLER_224_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13807_ _20198_/Q vssd1 vssd1 vccd1 vccd1 _14587_/A sky130_fd_sc_hd__inv_2
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17575_ _17575_/A vssd1 vssd1 vccd1 vccd1 _17576_/A sky130_fd_sc_hd__inv_2
X_14787_ _14787_/A _14787_/B vssd1 vssd1 vccd1 vccd1 _20123_/D sky130_fd_sc_hd__nor2_1
X_11999_ _20993_/Q _11999_/B vssd1 vssd1 vccd1 vccd1 _12000_/B sky130_fd_sc_hd__or2_1
XFILLER_16_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19314_ _20142_/CLK _19314_/D vssd1 vssd1 vccd1 vccd1 _19314_/Q sky130_fd_sc_hd__dfxtp_1
X_16526_ _16526_/A _16526_/B vssd1 vssd1 vccd1 vccd1 _16526_/Y sky130_fd_sc_hd__nor2_1
XFILLER_232_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13738_ _14575_/B vssd1 vssd1 vccd1 vccd1 _13738_/X sky130_fd_sc_hd__buf_1
XFILLER_220_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19245_ _17419_/Y _17420_/Y _17421_/Y _17422_/Y _19275_/S0 _21004_/Q vssd1 vssd1
+ vccd1 vccd1 _19245_/X sky130_fd_sc_hd__mux4_2
XFILLER_176_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16457_ _19305_/Q _16452_/X _11504_/X _16454_/X vssd1 vssd1 vccd1 vccd1 _19305_/D
+ sky130_fd_sc_hd__a22o_1
X_13669_ _20359_/Q _13667_/X _13550_/X _13668_/X vssd1 vssd1 vccd1 vccd1 _20359_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15408_ _19808_/Q _15405_/X _15350_/X _15406_/X vssd1 vssd1 vccd1 vccd1 _19808_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_176_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19176_ _19172_/X _19173_/X _19174_/X _19175_/X _20123_/Q _20124_/Q vssd1 vssd1 vccd1
+ vccd1 _19176_/X sky130_fd_sc_hd__mux4_2
XFILLER_191_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16388_ _19343_/Q _16385_/X _16210_/X _16386_/X vssd1 vssd1 vccd1 vccd1 _19343_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_129_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_116_HCLK_A clkbuf_opt_3_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18127_ _18126_/X _14096_/A _18850_/S vssd1 vssd1 vccd1 vccd1 _18127_/X sky130_fd_sc_hd__mux2_1
X_15339_ _15347_/A vssd1 vssd1 vccd1 vccd1 _15339_/X sky130_fd_sc_hd__buf_1
XFILLER_247_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18058_ _18321_/X _18024_/X _18359_/X _17995_/X _18057_/X vssd1 vssd1 vccd1 vccd1
+ _18059_/C sky130_fd_sc_hd__o221a_1
XANTENNA__18080__B _18083_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13713__B1 _13712_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17009_ _19978_/Q _17004_/A _19979_/Q vssd1 vssd1 vccd1 vccd1 _17009_/X sky130_fd_sc_hd__o21a_1
X_09900_ _09898_/X _20007_/Q _20008_/Q vssd1 vssd1 vccd1 vccd1 _09900_/Y sky130_fd_sc_hd__a21oi_1
X_20020_ _21419_/CLK _20020_/D repeater232/X vssd1 vssd1 vccd1 vccd1 _20020_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18652__A0 _17281_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09831_ _21448_/Q vssd1 vssd1 vccd1 vccd1 _15879_/A sky130_fd_sc_hd__buf_1
XFILLER_101_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09762_ _20152_/Q vssd1 vssd1 vccd1 vccd1 _09762_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18300__S _18680_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17207__A1 _18898_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17207__B2 _17157_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_26_HCLK clkbuf_opt_4_HCLK/A vssd1 vssd1 vccd1 vccd1 _21433_/CLK sky130_fd_sc_hd__clkbuf_16
X_09693_ _11739_/A vssd1 vssd1 vccd1 vccd1 _09693_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_39_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18955__A1 _21081_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12849__A _12849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20922_ _20930_/CLK _20922_/D repeater268/X vssd1 vssd1 vccd1 vccd1 _20922_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_4019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_214_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20853_ _20857_/CLK _20853_/D repeater243/X vssd1 vssd1 vccd1 vccd1 _20853_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20784_ _21406_/CLK _20784_/D repeater213/X vssd1 vssd1 vccd1 vccd1 _20784_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_23_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_168_HCLK clkbuf_opt_0_HCLK/A vssd1 vssd1 vccd1 vccd1 _21457_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_195_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21405_ _21405_/CLK _21405_/D repeater252/X vssd1 vssd1 vccd1 vccd1 _21405_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_163_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21336_ _21341_/CLK _21336_/D repeater204/X vssd1 vssd1 vccd1 vccd1 _21336_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_151_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_38_HCLK_A _20004_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21267_ _21417_/CLK _21267_/D repeater231/X vssd1 vssd1 vccd1 vccd1 _21267_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__14304__A _14304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18643__A0 _18848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11020_ _18992_/S vssd1 vssd1 vccd1 vccd1 _11596_/A sky130_fd_sc_hd__inv_2
X_20218_ _20220_/CLK _20218_/D repeater202/X vssd1 vssd1 vccd1 vccd1 _20218_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_2_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21198_ _21255_/CLK _21198_/D repeater241/X vssd1 vssd1 vccd1 vccd1 _21198_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__15457__B1 _15456_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_238_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20149_ _21239_/CLK _20149_/D repeater250/X vssd1 vssd1 vccd1 vccd1 _20149_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_106_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18210__S _18910_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_246_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12971_ _12966_/X _12970_/X _12751_/A _12969_/X vssd1 vssd1 vccd1 vccd1 _20702_/D
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__20118__CLK _21452_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14710_ _20156_/Q _14704_/X _12857_/A _14706_/X vssd1 vssd1 vccd1 vccd1 _20156_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_246_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11922_ _11142_/X _11921_/X _11142_/X _11921_/X vssd1 vssd1 vccd1 vccd1 _11926_/C
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_17_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12691__B1 _09649_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15690_ _15698_/A vssd1 vssd1 vccd1 vccd1 _15690_/X sky130_fd_sc_hd__buf_1
XPHY_4520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21052__RESET_B repeater225/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14641_ _14641_/A vssd1 vssd1 vccd1 vccd1 _14641_/Y sky130_fd_sc_hd__inv_2
XPHY_4553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11853_ _11848_/B _11851_/Y _11822_/B _11852_/X _11807_/A vssd1 vssd1 vccd1 vccd1
+ _11854_/A sky130_fd_sc_hd__o32a_1
XFILLER_122_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14432__A1 _21485_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19041__S _19046_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_214_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10804_ _10804_/A vssd1 vssd1 vccd1 vccd1 _10804_/Y sky130_fd_sc_hd__inv_2
X_17360_ _19616_/Q vssd1 vssd1 vccd1 vccd1 _17360_/Y sky130_fd_sc_hd__inv_2
XPHY_4597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11784_ _11784_/A vssd1 vssd1 vccd1 vccd1 _11784_/X sky130_fd_sc_hd__clkbuf_1
X_14572_ _14572_/A _14572_/B vssd1 vssd1 vccd1 vccd1 _14641_/A sky130_fd_sc_hd__or2_1
XPHY_3863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16311_ _16311_/A _16311_/B _16311_/C vssd1 vssd1 vccd1 vccd1 _16319_/A sky130_fd_sc_hd__or3_4
XPHY_3896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13523_ _13528_/A _13527_/A _13181_/C _13175_/A _13182_/B vssd1 vssd1 vccd1 vccd1
+ _13524_/B sky130_fd_sc_hd__o32a_1
XFILLER_198_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17291_ _21065_/Q vssd1 vssd1 vccd1 vccd1 _17291_/Y sky130_fd_sc_hd__inv_2
X_10735_ _19922_/Q _16760_/A vssd1 vssd1 vccd1 vccd1 _16765_/A sky130_fd_sc_hd__or2_1
XFILLER_41_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18880__S _18880_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19030_ _16870_/Y _20839_/Q _19046_/S vssd1 vssd1 vccd1 vccd1 _19946_/D sky130_fd_sc_hd__mux2_1
X_16242_ _19417_/Q _16240_/X _16009_/X _16241_/X vssd1 vssd1 vccd1 vccd1 _19417_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_13_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10666_ _10666_/A vssd1 vssd1 vccd1 vccd1 _10666_/Y sky130_fd_sc_hd__inv_2
X_13454_ _13714_/A vssd1 vssd1 vccd1 vccd1 _13454_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__19560__CLK _19706_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12405_ _12430_/A _12429_/A _12432_/A _12431_/A vssd1 vssd1 vccd1 vccd1 _12406_/C
+ sky130_fd_sc_hd__or4_4
X_16173_ _16173_/A vssd1 vssd1 vccd1 vccd1 _16173_/X sky130_fd_sc_hd__buf_1
X_13385_ _13601_/B vssd1 vssd1 vccd1 vccd1 _17174_/B sky130_fd_sc_hd__buf_6
XFILLER_182_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10597_ _21334_/Q _20762_/Q _21334_/Q _20762_/Q vssd1 vssd1 vccd1 vccd1 _10597_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_15124_ _15123_/Y _20070_/Q _20444_/Q _15069_/A vssd1 vssd1 vccd1 vccd1 _15124_/X
+ sky130_fd_sc_hd__o22a_1
X_12336_ _12373_/A vssd1 vssd1 vccd1 vccd1 _12364_/A sky130_fd_sc_hd__inv_2
Xoutput109 _17828_/Y vssd1 vssd1 vccd1 vccd1 HRDATA[8] sky130_fd_sc_hd__clkbuf_2
XFILLER_217_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15055_ _20047_/Q vssd1 vssd1 vccd1 vccd1 _15062_/A sky130_fd_sc_hd__inv_2
X_12267_ _20934_/Q _12263_/Y _20928_/Q _12264_/Y _12266_/X vssd1 vssd1 vccd1 vccd1
+ _12278_/B sky130_fd_sc_hd__o221a_1
X_19932_ _21242_/CLK _19932_/D repeater189/X vssd1 vssd1 vccd1 vccd1 _19932_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18634__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11218_ _21205_/Q _11213_/X _09666_/X _11214_/X vssd1 vssd1 vccd1 vccd1 _21205_/D
+ sky130_fd_sc_hd__a22o_1
X_14006_ _14006_/A vssd1 vssd1 vccd1 vccd1 _14006_/Y sky130_fd_sc_hd__inv_2
X_19863_ _21164_/CLK _19863_/D repeater225/X vssd1 vssd1 vccd1 vccd1 _19863_/Q sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_49_HCLK clkbuf_4_9_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _21087_/CLK sky130_fd_sc_hd__clkbuf_16
X_12198_ _20360_/Q vssd1 vssd1 vccd1 vccd1 _12198_/Y sky130_fd_sc_hd__inv_2
Xoutput80 _17865_/Y vssd1 vssd1 vccd1 vccd1 HRDATA[10] sky130_fd_sc_hd__clkbuf_2
XFILLER_96_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput91 _17989_/X vssd1 vssd1 vccd1 vccd1 HRDATA[20] sky130_fd_sc_hd__clkbuf_2
XFILLER_150_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18814_ _18848_/A0 _14121_/Y _18902_/S vssd1 vssd1 vccd1 vccd1 _18814_/X sky130_fd_sc_hd__mux2_1
X_11149_ _15609_/A _15609_/B _15594_/A vssd1 vssd1 vccd1 vccd1 _11149_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_122_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19794_ _19811_/CLK _19794_/D vssd1 vssd1 vccd1 vccd1 _19794_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18745_ _17544_/Y _20742_/Q _18775_/S vssd1 vssd1 vccd1 vccd1 _18745_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15957_ _19557_/Q _15954_/X _15887_/X _15956_/X vssd1 vssd1 vccd1 vccd1 _19557_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18937__A1 _21139_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19285__S1 _21017_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14908_ _20573_/Q _15004_/A _14906_/Y _20084_/Q _14907_/X vssd1 vssd1 vccd1 vccd1
+ _14918_/B sky130_fd_sc_hd__o221a_1
XANTENNA__12682__B1 _09633_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18676_ _17756_/Y _19206_/X _18930_/S vssd1 vssd1 vccd1 vccd1 _18676_/X sky130_fd_sc_hd__mux2_1
X_15888_ _15896_/A vssd1 vssd1 vccd1 vccd1 _15897_/A sky130_fd_sc_hd__inv_2
XFILLER_64_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17627_ _14657_/X _17276_/Y _20172_/Q _17131_/Y vssd1 vssd1 vccd1 vccd1 _17627_/X
+ sky130_fd_sc_hd__a22o_1
X_14839_ _20095_/Q vssd1 vssd1 vccd1 vccd1 _14961_/C sky130_fd_sc_hd__inv_2
XANTENNA__14423__B2 _20029_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_224_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17558_ _17552_/Y _17553_/X _17554_/Y _17387_/X _17557_/X vssd1 vssd1 vccd1 vccd1
+ _17558_/X sky130_fd_sc_hd__o221a_1
XFILLER_211_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16509_ _16681_/B _20000_/Q _16509_/C vssd1 vssd1 vccd1 vccd1 _16510_/A sky130_fd_sc_hd__and3_1
XFILLER_177_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17489_ _19426_/Q vssd1 vssd1 vccd1 vccd1 _17489_/Y sky130_fd_sc_hd__inv_2
XFILLER_176_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19228_ _17513_/Y _17514_/Y _17515_/Y _17516_/Y _20130_/Q _20131_/Q vssd1 vssd1 vccd1
+ vccd1 _19228_/X sky130_fd_sc_hd__mux4_2
XFILLER_177_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20704__RESET_B repeater210/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19114__A1 _10985_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19159_ _19692_/Q _19380_/Q _19676_/Q _19668_/Q _19285_/S0 _21017_/Q vssd1 vssd1
+ vccd1 vccd1 _19159_/X sky130_fd_sc_hd__mux4_2
XFILLER_11_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21121_ _21121_/CLK _21121_/D repeater237/X vssd1 vssd1 vccd1 vccd1 _21121_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_160_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21052_ _21164_/CLK _21052_/D repeater225/X vssd1 vssd1 vccd1 vccd1 _21052_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20003_ _20331_/CLK _20003_/D repeater190/X vssd1 vssd1 vccd1 vccd1 _20003_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_143_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09814_ _09827_/A vssd1 vssd1 vccd1 vccd1 _09829_/A sky130_fd_sc_hd__inv_2
XFILLER_101_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09745_ _20144_/Q vssd1 vssd1 vccd1 vccd1 _09745_/Y sky130_fd_sc_hd__inv_2
XFILLER_100_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19276__S1 _21006_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19958__RESET_B repeater184/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09676_ _12548_/A vssd1 vssd1 vccd1 vccd1 _09676_/X sky130_fd_sc_hd__buf_4
X_20905_ _20908_/CLK _20905_/D repeater217/X vssd1 vssd1 vccd1 vccd1 _20905_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20836_ _20930_/CLK _20836_/D repeater257/X vssd1 vssd1 vccd1 vccd1 _20836_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20767_ _21342_/CLK _20767_/D repeater191/X vssd1 vssd1 vccd1 vccd1 _20767_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10520_ _21308_/Q _10518_/Y _21301_/Q _18034_/A vssd1 vssd1 vccd1 vccd1 _10520_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20560__CLK _20592_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20698_ _21481_/CLK _20698_/D repeater205/X vssd1 vssd1 vccd1 vccd1 _20698_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_155_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10451_ _21290_/Q _20679_/Q _10766_/A _10450_/Y vssd1 vssd1 vccd1 vccd1 _10451_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_164_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18205__S _18908_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19200__S1 _20131_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13170_ _20601_/Q _13165_/X _13169_/X _13167_/X vssd1 vssd1 vccd1 vccd1 _20601_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_201_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10382_ _21367_/Q _10380_/Y _10283_/B _10381_/X vssd1 vssd1 vccd1 vccd1 _21367_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA_clkbuf_leaf_162_HCLK_A clkbuf_opt_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12121_ _20388_/Q vssd1 vssd1 vccd1 vccd1 _18029_/A sky130_fd_sc_hd__inv_2
XFILLER_108_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21319_ _21319_/CLK _21319_/D repeater191/X vssd1 vssd1 vccd1 vccd1 _21319_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_190_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12052_ _12322_/A _20383_/Q _20969_/Q _12051_/Y vssd1 vssd1 vccd1 vccd1 _12052_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_78_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11003_ _21014_/Q vssd1 vssd1 vccd1 vccd1 _11003_/X sky130_fd_sc_hd__buf_1
XANTENNA__19036__S _19046_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16860_ _19944_/Q vssd1 vssd1 vccd1 vccd1 _16863_/A sky130_fd_sc_hd__inv_2
XANTENNA__21066__CLK _21134_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_237_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15811_ _19623_/Q _15807_/X _09838_/X _15808_/X vssd1 vssd1 vccd1 vccd1 _19623_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17064__B _17064_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__21233__RESET_B repeater270/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16791_ _16791_/A _16791_/B vssd1 vssd1 vccd1 vccd1 _16791_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__19267__S1 _20131_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18875__S _18875_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18530_ _17943_/Y _20790_/Q _18644_/S vssd1 vssd1 vccd1 vccd1 _18530_/X sky130_fd_sc_hd__mux2_1
XFILLER_93_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15742_ _16311_/A _15778_/B _16311_/C vssd1 vssd1 vccd1 vccd1 _15750_/A sky130_fd_sc_hd__or3_4
X_12954_ _14262_/A vssd1 vssd1 vccd1 vccd1 _12954_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__17999__B _17999_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18461_ _18845_/A0 _10499_/Y _18884_/S vssd1 vssd1 vccd1 vccd1 _18461_/X sky130_fd_sc_hd__mux2_1
X_11905_ _11913_/A _15374_/B vssd1 vssd1 vccd1 vccd1 _11906_/A sky130_fd_sc_hd__or2_1
XFILLER_233_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output110_A _17847_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15673_ _15673_/A _16311_/B _15722_/C vssd1 vssd1 vccd1 vccd1 _15681_/A sky130_fd_sc_hd__or3_4
XPHY_4350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12885_ _20738_/Q _12874_/X _12884_/X _12876_/X vssd1 vssd1 vccd1 vccd1 _20738_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17412_ _19425_/Q vssd1 vssd1 vccd1 vccd1 _17412_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17080__A _17080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14624_ _14624_/A vssd1 vssd1 vccd1 vccd1 _14624_/X sky130_fd_sc_hd__clkbuf_2
XPHY_4383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18392_ _18391_/X _14926_/Y _18907_/S vssd1 vssd1 vccd1 vccd1 _18392_/X sky130_fd_sc_hd__mux2_2
X_11836_ _11836_/A vssd1 vssd1 vccd1 vccd1 _21035_/D sky130_fd_sc_hd__inv_2
XPHY_4394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17343_ _19776_/Q vssd1 vssd1 vccd1 vccd1 _17343_/Y sky130_fd_sc_hd__inv_2
XPHY_3682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14555_ _14535_/Y _14544_/X _14769_/A vssd1 vssd1 vccd1 vccd1 _14555_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA_repeater260_A repeater267/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11767_ _19084_/X _11764_/X _21050_/Q _11765_/X vssd1 vssd1 vccd1 vccd1 _21050_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13506_ _14258_/A vssd1 vssd1 vccd1 vccd1 _13506_/X sky130_fd_sc_hd__clkbuf_2
X_17274_ _11424_/Y _16575_/Y _17273_/X vssd1 vssd1 vccd1 vccd1 _19914_/D sky130_fd_sc_hd__o21ai_1
X_10718_ _10718_/A vssd1 vssd1 vccd1 vccd1 _10718_/Y sky130_fd_sc_hd__inv_2
XPHY_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14486_ _14486_/A vssd1 vssd1 vccd1 vccd1 _14486_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20186__RESET_B repeater193/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11698_ _11704_/A vssd1 vssd1 vccd1 vccd1 _11705_/A sky130_fd_sc_hd__inv_2
X_19013_ _16940_/X _20410_/Q _19019_/S vssd1 vssd1 vccd1 vccd1 _19963_/D sky130_fd_sc_hd__mux2_1
X_16225_ _19425_/Q _16223_/X _16120_/X _16224_/X vssd1 vssd1 vccd1 vccd1 _19425_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_228_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13437_ _13447_/A vssd1 vssd1 vccd1 vccd1 _13437_/X sky130_fd_sc_hd__buf_1
X_10649_ _10649_/A _10729_/C _10649_/C vssd1 vssd1 vccd1 vccd1 _21340_/D sky130_fd_sc_hd__nor3_2
XFILLER_174_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrebuffer2 _20027_/Q vssd1 vssd1 vccd1 vccd1 _18052_/A sky130_fd_sc_hd__dlygate4sd1_1
X_16156_ _19459_/Q _16151_/X _16137_/X _16153_/X vssd1 vssd1 vccd1 vccd1 _19459_/D
+ sky130_fd_sc_hd__a22o_1
X_13368_ _20508_/Q _13365_/X _13154_/X _13366_/X vssd1 vssd1 vccd1 vccd1 _20508_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_170_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15669__B1 _15588_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15107_ _20440_/Q vssd1 vssd1 vccd1 vccd1 _15107_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16866__C1 _16779_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12319_ _12319_/A _12319_/B vssd1 vssd1 vccd1 vccd1 _12362_/A sky130_fd_sc_hd__or2_1
X_16087_ _16087_/A vssd1 vssd1 vccd1 vccd1 _16087_/X sky130_fd_sc_hd__buf_1
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13299_ _13299_/A vssd1 vssd1 vccd1 vccd1 _13321_/A sky130_fd_sc_hd__buf_1
XFILLER_244_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_21_HCLK_A clkbuf_4_3_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19915_ _21167_/CLK _19915_/D repeater225/X vssd1 vssd1 vccd1 vccd1 _19915_/Q sky130_fd_sc_hd__dfrtp_1
X_15038_ _20064_/Q vssd1 vssd1 vccd1 vccd1 _15112_/A sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_84_HCLK_A clkbuf_4_12_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19846_ _20042_/CLK _19846_/D repeater219/X vssd1 vssd1 vccd1 vccd1 _19846_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_69_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16989_ _19974_/Q _16989_/B vssd1 vssd1 vccd1 vccd1 _16989_/X sky130_fd_sc_hd__and2_1
X_19777_ _19777_/CLK _19777_/D vssd1 vssd1 vccd1 vccd1 _19777_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__18785__S _18907_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19258__S1 _20131_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18728_ _17079_/Y _12125_/Y _18908_/S vssd1 vssd1 vccd1 vccd1 _18728_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12655__B1 _12651_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18659_ _17281_/X _18071_/Y _18874_/S vssd1 vssd1 vccd1 vccd1 _18659_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20956__RESET_B repeater187/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20621_ _20622_/CLK _20621_/D repeater195/X vssd1 vssd1 vccd1 vccd1 _20621_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20552_ _20947_/CLK _20552_/D repeater266/X vssd1 vssd1 vccd1 vccd1 _20552_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_137_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20483_ _20944_/CLK _20483_/D repeater273/X vssd1 vssd1 vccd1 vccd1 _20483_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__19194__S0 _19280_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21104_ _21417_/CLK _21104_/D repeater231/X vssd1 vssd1 vccd1 vccd1 _21104_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_133_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21035_ _21207_/CLK _21035_/D repeater242/X vssd1 vssd1 vccd1 vccd1 _21035_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_247_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18695__S _18908_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19249__S1 _20131_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09728_ _11063_/A _20158_/Q _21238_/Q _09727_/Y vssd1 vssd1 vccd1 vccd1 _09728_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_228_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09659_ _12863_/A vssd1 vssd1 vccd1 vccd1 _09659_/X sky130_fd_sc_hd__buf_4
XANTENNA__20697__RESET_B repeater193/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10121__B2 _20774_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12670_ input54/X vssd1 vssd1 vccd1 vccd1 _12670_/X sky130_fd_sc_hd__clkbuf_4
XPHY_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20626__RESET_B repeater193/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11621_ _11621_/A _11621_/B vssd1 vssd1 vccd1 vccd1 _11625_/B sky130_fd_sc_hd__or2_1
XPHY_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20819_ _21374_/CLK _20819_/D repeater256/X vssd1 vssd1 vccd1 vccd1 _20819_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13071__B1 _12922_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_211_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14340_ _20225_/Q vssd1 vssd1 vccd1 vccd1 _14461_/D sky130_fd_sc_hd__inv_2
XPHY_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11552_ _11562_/A vssd1 vssd1 vccd1 vccd1 _11552_/X sky130_fd_sc_hd__buf_1
XPHY_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15899__B1 _15791_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10503_ _21298_/Q vssd1 vssd1 vccd1 vccd1 _10774_/A sky130_fd_sc_hd__inv_2
XPHY_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11483_ _19104_/X _11480_/X _21154_/Q _11481_/X vssd1 vssd1 vccd1 vccd1 _21154_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_10_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14271_ _20245_/Q _14267_/X _13712_/X _14268_/X vssd1 vssd1 vccd1 vccd1 _20245_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16010_ _16010_/A vssd1 vssd1 vccd1 vccd1 _16010_/X sky130_fd_sc_hd__buf_1
XANTENNA__12177__A2 _20361_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19185__S0 _19280_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13374__A1 _20504_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input71_A MSI_S2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10434_ _21304_/Q vssd1 vssd1 vccd1 vccd1 _10780_/A sky130_fd_sc_hd__inv_2
XANTENNA__18837__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13222_ _20582_/Q _13215_/X _13221_/X _13217_/X vssd1 vssd1 vccd1 vccd1 _20582_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_164_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21485__RESET_B repeater200/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10365_ _21375_/Q _10290_/Y _10291_/Y _10290_/A _10364_/X vssd1 vssd1 vccd1 vccd1
+ _21375_/D sky130_fd_sc_hd__o221a_1
X_13153_ _20610_/Q _13150_/X _13151_/X _13152_/X vssd1 vssd1 vccd1 vccd1 _20610_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_152_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14323__B1 _20124_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12104_ _20970_/Q vssd1 vssd1 vccd1 vccd1 _12323_/A sky130_fd_sc_hd__inv_2
X_17961_ _18178_/X _17928_/X _18188_/X _17960_/X vssd1 vssd1 vccd1 vccd1 _17961_/X
+ sky130_fd_sc_hd__o22a_2
X_13084_ _20647_/Q _13079_/X _12855_/X _13081_/X vssd1 vssd1 vccd1 vccd1 _20647_/D
+ sky130_fd_sc_hd__a22o_1
X_10296_ _20722_/Q vssd1 vssd1 vccd1 vccd1 _10296_/Y sky130_fd_sc_hd__inv_2
XFILLER_239_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16912_ _19957_/Q vssd1 vssd1 vccd1 vccd1 _16914_/A sky130_fd_sc_hd__inv_2
X_12035_ _20964_/Q vssd1 vssd1 vccd1 vccd1 _12317_/A sky130_fd_sc_hd__inv_2
X_19700_ _20432_/CLK _19700_/D vssd1 vssd1 vccd1 vccd1 _19700_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11688__A1 _21084_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12885__B1 _12884_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17892_ _14702_/A _17886_/X _17888_/X _17891_/X vssd1 vssd1 vccd1 vccd1 _17892_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_77_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16843_ _16843_/A _16843_/B vssd1 vssd1 vccd1 vccd1 _16844_/A sky130_fd_sc_hd__or2_1
X_19631_ _21021_/CLK _19631_/D vssd1 vssd1 vccd1 vccd1 _19631_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19562_ _19812_/CLK _19562_/D vssd1 vssd1 vccd1 vccd1 _19562_/Q sky130_fd_sc_hd__dfxtp_1
X_16774_ _16774_/A _16774_/B vssd1 vssd1 vccd1 vccd1 _16774_/Y sky130_fd_sc_hd__nor2_1
XFILLER_46_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13986_ _13986_/A vssd1 vssd1 vccd1 vccd1 _13986_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18513_ _18848_/A0 _14130_/Y _18902_/S vssd1 vssd1 vccd1 vccd1 _18513_/X sky130_fd_sc_hd__mux2_1
XFILLER_218_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15725_ _16231_/A vssd1 vssd1 vccd1 vccd1 _15725_/X sky130_fd_sc_hd__buf_1
X_19493_ _21040_/CLK _19493_/D vssd1 vssd1 vccd1 vccd1 _19493_/Q sky130_fd_sc_hd__dfxtp_1
X_12937_ _12961_/A vssd1 vssd1 vccd1 vccd1 _12937_/X sky130_fd_sc_hd__buf_1
XFILLER_233_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18444_ _18443_/X _12263_/Y _18910_/S vssd1 vssd1 vccd1 vccd1 _18444_/X sky130_fd_sc_hd__mux2_1
XANTENNA__15323__A _15329_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15656_ _15666_/A vssd1 vssd1 vccd1 vccd1 _15656_/X sky130_fd_sc_hd__buf_1
XPHY_4180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12868_ _12876_/A vssd1 vssd1 vccd1 vccd1 _12868_/X sky130_fd_sc_hd__buf_1
XFILLER_233_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14607_ _14639_/A vssd1 vssd1 vccd1 vccd1 _14607_/X sky130_fd_sc_hd__buf_2
XFILLER_21_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18375_ _17978_/Y _21483_/Q _18669_/S vssd1 vssd1 vccd1 vccd1 _18375_/X sky130_fd_sc_hd__mux2_1
X_11819_ _21039_/Q _11803_/X _11815_/X _10966_/Y _11818_/Y vssd1 vssd1 vccd1 vccd1
+ _11820_/A sky130_fd_sc_hd__o32a_1
XFILLER_21_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15587_ _19729_/Q _15584_/X _15585_/X _15586_/X vssd1 vssd1 vccd1 vccd1 _19729_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13062__B1 _12996_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12799_ _20780_/Q _12797_/X _12544_/X _12798_/X vssd1 vssd1 vccd1 vccd1 _20780_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_239_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17326_ _17928_/A vssd1 vssd1 vccd1 vccd1 _17326_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_175_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14538_ _20134_/Q vssd1 vssd1 vccd1 vccd1 _15832_/B sky130_fd_sc_hd__inv_2
Xclkbuf_2_2_0_HCLK clkbuf_2_3_0_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_187_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17257_ _19479_/Q vssd1 vssd1 vccd1 vccd1 _17257_/Y sky130_fd_sc_hd__inv_2
X_14469_ _14488_/A vssd1 vssd1 vccd1 vccd1 _14469_/X sky130_fd_sc_hd__buf_2
X_16208_ _16208_/A vssd1 vssd1 vccd1 vccd1 _16208_/X sky130_fd_sc_hd__buf_1
XANTENNA__19176__S0 _20123_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17188_ _20811_/Q vssd1 vssd1 vccd1 vccd1 _17188_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16139_ _21450_/Q vssd1 vssd1 vccd1 vccd1 _16139_/X sky130_fd_sc_hd__buf_1
XFILLER_115_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19829_ _19835_/CLK _19829_/D vssd1 vssd1 vccd1 vccd1 _19829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12857__A _12857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20790__RESET_B repeater255/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_240_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20604_ _21302_/CLK _20604_/D repeater209/X vssd1 vssd1 vccd1 vccd1 _20604_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__12800__B1 _12548_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20535_ _20929_/CLK _20535_/D repeater265/X vssd1 vssd1 vccd1 vccd1 _20535_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__19621__CLK _21452_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_229_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19167__S0 _19280_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18819__A0 _18818_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20466_ _20937_/CLK _20466_/D repeater277/X vssd1 vssd1 vccd1 vccd1 _20466_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_181_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20397_ _20809_/CLK _20397_/D repeater270/X vssd1 vssd1 vccd1 vccd1 _20397_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_106_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09980__B1 _09693_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10150_ _10150_/A _10196_/A vssd1 vssd1 vccd1 vccd1 _10151_/B sky130_fd_sc_hd__or2_2
XANTENNA__10590__B2 _20750_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19973__RESET_B repeater184/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10081_ _20779_/Q vssd1 vssd1 vccd1 vccd1 _10081_/Y sky130_fd_sc_hd__inv_2
XFILLER_102_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21018_ _21431_/CLK _21018_/D repeater238/X vssd1 vssd1 vccd1 vccd1 _21018_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_87_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20878__RESET_B repeater243/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13840_ _20323_/Q _14636_/A _13735_/Y vssd1 vssd1 vccd1 vccd1 _20323_/D sky130_fd_sc_hd__o21a_1
XFILLER_74_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13771_ _20187_/Q vssd1 vssd1 vccd1 vccd1 _14576_/A sky130_fd_sc_hd__inv_2
XFILLER_74_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10983_ _10983_/A vssd1 vssd1 vccd1 vccd1 _19115_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_28_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15510_ _19765_/Q _15507_/X _15450_/X _15509_/X vssd1 vssd1 vccd1 vccd1 _19765_/D
+ sky130_fd_sc_hd__a22o_1
X_12722_ _17177_/A _17378_/A vssd1 vssd1 vccd1 vccd1 _13106_/B sky130_fd_sc_hd__or2_4
X_16490_ _16526_/A _16490_/B vssd1 vssd1 vccd1 vccd1 _16490_/X sky130_fd_sc_hd__or2_1
XFILLER_215_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20460__RESET_B repeater276/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15441_ _15441_/A vssd1 vssd1 vccd1 vccd1 _15441_/X sky130_fd_sc_hd__buf_1
XANTENNA__13044__B1 _12881_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12653_ _12687_/A vssd1 vssd1 vccd1 vccd1 _12680_/A sky130_fd_sc_hd__buf_1
XPHY_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11604_ _18989_/X _11598_/X _21117_/Q _11600_/X vssd1 vssd1 vccd1 vccd1 _21117_/D
+ sky130_fd_sc_hd__a22o_1
X_18160_ _18159_/X _16839_/Y _18667_/S vssd1 vssd1 vccd1 vccd1 _18160_/X sky130_fd_sc_hd__mux2_1
XPHY_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15372_ _15559_/A vssd1 vssd1 vccd1 vccd1 _15542_/B sky130_fd_sc_hd__buf_1
XPHY_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12584_ _20884_/Q _12581_/X _18236_/X _12583_/X vssd1 vssd1 vccd1 vccd1 _20884_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17111_ _17254_/A vssd1 vssd1 vccd1 vccd1 _17773_/B sky130_fd_sc_hd__buf_1
XPHY_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14323_ _20124_/Q _14322_/X _20124_/Q _14322_/X vssd1 vssd1 vccd1 vccd1 _14324_/D
+ sky130_fd_sc_hd__a2bb2o_1
XPHY_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11535_ _11535_/A vssd1 vssd1 vccd1 vccd1 _11535_/X sky130_fd_sc_hd__buf_1
XFILLER_11_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18091_ _20841_/Q vssd1 vssd1 vccd1 vccd1 _18091_/Y sky130_fd_sc_hd__inv_2
XPHY_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17730__B1 _18680_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19158__S0 _19285_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17042_ _21247_/Q vssd1 vssd1 vccd1 vccd1 _17042_/Y sky130_fd_sc_hd__inv_2
X_14254_ _19989_/Q _12498_/Y _20252_/Q _16689_/A vssd1 vssd1 vccd1 vccd1 _20252_/D
+ sky130_fd_sc_hd__o22a_1
X_11466_ _19093_/X _11461_/X _21165_/Q _11463_/X vssd1 vssd1 vccd1 vccd1 _21165_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_143_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13205_ _20589_/Q _13200_/X _13003_/X _13201_/X vssd1 vssd1 vccd1 vccd1 _20589_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18286__A1 _10602_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13110__B _13261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10417_ _10262_/A _10262_/B _10415_/Y _10375_/X vssd1 vssd1 vccd1 vccd1 _21346_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_136_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11397_ _15310_/A _11327_/X _11412_/C _11357_/A _11396_/X vssd1 vssd1 vccd1 vccd1
+ _21184_/D sky130_fd_sc_hd__a32o_1
X_14185_ _14207_/A vssd1 vssd1 vccd1 vccd1 _14185_/X sky130_fd_sc_hd__buf_2
XANTENNA__16702__A _16720_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13136_ _20616_/Q _13132_/X _12930_/X _13133_/X vssd1 vssd1 vccd1 vccd1 _20616_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09971__B1 _09663_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10348_ _20730_/Q vssd1 vssd1 vccd1 vccd1 _10348_/Y sky130_fd_sc_hd__inv_2
XFILLER_225_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18993_ _21250_/Q _17028_/Y _18993_/S vssd1 vssd1 vccd1 vccd1 _18993_/X sky130_fd_sc_hd__mux2_1
XFILLER_151_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12858__B1 _12857_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17944_ _20828_/Q _17944_/B vssd1 vssd1 vccd1 vccd1 _17944_/Y sky130_fd_sc_hd__nand2_1
X_10279_ _10279_/A _10279_/B vssd1 vssd1 vccd1 vccd1 _10385_/A sky130_fd_sc_hd__or2_1
X_13067_ _13073_/A vssd1 vssd1 vccd1 vccd1 _13067_/X sky130_fd_sc_hd__buf_1
XFILLER_239_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater206 repeater207/X vssd1 vssd1 vccd1 vccd1 repeater206/X sky130_fd_sc_hd__buf_8
Xrepeater217 repeater218/X vssd1 vssd1 vccd1 vccd1 repeater217/X sky130_fd_sc_hd__buf_8
X_12018_ _12030_/A vssd1 vssd1 vccd1 vccd1 _12018_/X sky130_fd_sc_hd__buf_1
XFILLER_38_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_239_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater228 repeater229/X vssd1 vssd1 vccd1 vccd1 repeater228/X sky130_fd_sc_hd__buf_6
X_17875_ _20344_/Q vssd1 vssd1 vccd1 vccd1 _17875_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11530__B1 _10884_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater239 repeater240/X vssd1 vssd1 vccd1 vccd1 repeater239/X sky130_fd_sc_hd__buf_6
XFILLER_120_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19614_ _20137_/CLK _19614_/D vssd1 vssd1 vccd1 vccd1 _19614_/Q sky130_fd_sc_hd__dfxtp_1
X_16826_ _19937_/Q vssd1 vssd1 vccd1 vccd1 _16830_/A sky130_fd_sc_hd__inv_2
XFILLER_93_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_242_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16757_ _19920_/Q _16756_/A _16755_/Y _16756_/Y vssd1 vssd1 vccd1 vccd1 _16758_/B
+ sky130_fd_sc_hd__o22a_1
X_19545_ _19784_/CLK _19545_/D vssd1 vssd1 vccd1 vccd1 _19545_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13283__B1 _13282_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13969_ _13987_/A vssd1 vssd1 vccd1 vccd1 _13969_/X sky130_fd_sc_hd__buf_1
XFILLER_222_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15708_ _15722_/A _16311_/B _15708_/C vssd1 vssd1 vccd1 vccd1 _15716_/A sky130_fd_sc_hd__or3_4
XANTENNA__10636__A2 _10635_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16688_ _16688_/A _16688_/B vssd1 vssd1 vccd1 vccd1 _19875_/D sky130_fd_sc_hd__nor2_1
X_19476_ _20432_/CLK _19476_/D vssd1 vssd1 vccd1 vccd1 _19476_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18427_ _17281_/X _17877_/Y _18835_/S vssd1 vssd1 vccd1 vccd1 _18427_/X sky130_fd_sc_hd__mux2_1
X_15639_ _15756_/A _15756_/B _16465_/C vssd1 vssd1 vccd1 vccd1 _15647_/A sky130_fd_sc_hd__or3_4
XANTENNA__20130__RESET_B repeater249/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18358_ _17281_/X _18054_/Y _18909_/S vssd1 vssd1 vccd1 vccd1 _18358_/X sky130_fd_sc_hd__mux2_1
XANTENNA__18083__B _18083_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17309_ _17299_/Y _17175_/B _17302_/X _17308_/X vssd1 vssd1 vccd1 vccd1 _17309_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_30_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18289_ _17816_/Y _16917_/Y _18680_/S vssd1 vssd1 vccd1 vccd1 _18289_/X sky130_fd_sc_hd__mux2_2
XANTENNA__19149__S0 _19285_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20320_ _20322_/CLK _20320_/D repeater262/X vssd1 vssd1 vccd1 vccd1 _20320_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__21336__RESET_B repeater204/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20251_ _21147_/CLK _20251_/D repeater215/X vssd1 vssd1 vccd1 vccd1 _20251_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_134_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17708__A _20744_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18303__S _18908_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09962__B1 _09702_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20182_ _21483_/CLK _20182_/D repeater193/X vssd1 vssd1 vccd1 vccd1 _20182_/Q sky130_fd_sc_hd__dfrtp_1
X_09993_ _09991_/Y _17037_/A _09991_/Y _17037_/A vssd1 vssd1 vccd1 vccd1 _10017_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_130_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21127__CLK _21134_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_215_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20971__RESET_B repeater187/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20218__RESET_B repeater202/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11491__A _20889_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_231_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09796__A3 input74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13211__A input51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11320_ _12515_/A vssd1 vssd1 vccd1 vccd1 _16587_/A sky130_fd_sc_hd__buf_1
XFILLER_193_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20518_ _20944_/CLK _20518_/D repeater275/X vssd1 vssd1 vccd1 vccd1 _20518_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_180_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11251_ _11251_/A vssd1 vssd1 vccd1 vccd1 _11251_/X sky130_fd_sc_hd__buf_1
XANTENNA__18268__A1 _20795_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20449_ _20476_/CLK _20449_/D repeater183/X vssd1 vssd1 vccd1 vccd1 _20449_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21006__RESET_B repeater235/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18213__S _18748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09953__B1 _09670_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10202_ _10202_/A _10216_/A vssd1 vssd1 vccd1 vccd1 _10203_/B sky130_fd_sc_hd__or2_1
X_11182_ _11182_/A vssd1 vssd1 vccd1 vccd1 _17290_/A sky130_fd_sc_hd__buf_2
XFILLER_133_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11666__A _21071_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10133_ _20796_/Q vssd1 vssd1 vccd1 vccd1 _10133_/Y sky130_fd_sc_hd__inv_2
XFILLER_192_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15990_ _19540_/Q _15986_/X _15973_/X _15988_/X vssd1 vssd1 vccd1 vccd1 _19540_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input34_A HRESETn vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14941_ _14937_/Y _20101_/Q _20583_/Q _14961_/A _14940_/X vssd1 vssd1 vccd1 vccd1
+ _14948_/B sky130_fd_sc_hd__o221a_1
X_10064_ _21393_/Q vssd1 vssd1 vccd1 vccd1 _10154_/A sky130_fd_sc_hd__inv_2
XFILLER_248_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_82_HCLK clkbuf_4_13_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _21302_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_236_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19044__S _19046_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18440__A1 _20346_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17660_ _18730_/X _17401_/X _18735_/X _17320_/X vssd1 vssd1 vccd1 vccd1 _17660_/X
+ sky130_fd_sc_hd__o22a_1
X_14872_ _14961_/A _14872_/B vssd1 vssd1 vccd1 vccd1 _14984_/A sky130_fd_sc_hd__or2_1
XFILLER_208_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16611_ _16609_/A _16546_/A _16610_/Y _16541_/X vssd1 vssd1 vccd1 vccd1 _16611_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_91_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13823_ _13818_/Y _20197_/Q _13819_/Y _20185_/Q _13822_/X vssd1 vssd1 vccd1 vccd1
+ _13836_/B sky130_fd_sc_hd__o221a_1
X_17591_ _19475_/Q vssd1 vssd1 vccd1 vccd1 _17591_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19667__CLK _19813_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18883__S _18901_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16542_ _16537_/Y _16539_/X _16541_/X vssd1 vssd1 vccd1 vccd1 _16542_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_141_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19330_ _19834_/CLK _19330_/D vssd1 vssd1 vccd1 vccd1 _19330_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13754_ _13749_/Y _20203_/Q _20613_/Q _14579_/A _13753_/X vssd1 vssd1 vccd1 vccd1
+ _13761_/C sky130_fd_sc_hd__o221a_1
XFILLER_232_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10966_ _21039_/Q vssd1 vssd1 vccd1 vccd1 _10966_/Y sky130_fd_sc_hd__inv_2
XFILLER_189_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12705_ _20816_/Q _12701_/X _12550_/X _12702_/X vssd1 vssd1 vccd1 vccd1 _20816_/D
+ sky130_fd_sc_hd__a22o_1
X_19261_ _19257_/X _19258_/X _19259_/X _19260_/X _20132_/Q _20133_/Q vssd1 vssd1 vccd1
+ vccd1 _19261_/X sky130_fd_sc_hd__mux4_2
XANTENNA__17400__C1 _17399_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_231_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13017__B1 _12932_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16473_ _16473_/A vssd1 vssd1 vccd1 vccd1 _16473_/X sky130_fd_sc_hd__buf_1
XANTENNA_repeater173_A _18879_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13685_ _13685_/A vssd1 vssd1 vccd1 vccd1 _13706_/A sky130_fd_sc_hd__clkbuf_2
X_10897_ _21252_/Q _10888_/X _10896_/X _10890_/X vssd1 vssd1 vccd1 vccd1 _21252_/D
+ sky130_fd_sc_hd__a22o_1
X_18212_ _18211_/X _14411_/Y _18669_/S vssd1 vssd1 vccd1 vccd1 _18212_/X sky130_fd_sc_hd__mux2_1
X_15424_ _15424_/A vssd1 vssd1 vccd1 vccd1 _15424_/X sky130_fd_sc_hd__clkbuf_2
XPHY_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12636_ input28/X _12631_/X _20848_/Q _12632_/X vssd1 vssd1 vccd1 vccd1 _20848_/D
+ sky130_fd_sc_hd__o22a_1
X_19192_ _19708_/Q _19572_/Q _19564_/Q _19556_/Q _19280_/S0 _20122_/Q vssd1 vssd1
+ vccd1 vccd1 _19192_/X sky130_fd_sc_hd__mux4_2
XPHY_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18143_ _18142_/X _14416_/Y _18669_/S vssd1 vssd1 vccd1 vccd1 _18143_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15355_ _15592_/A vssd1 vssd1 vccd1 vccd1 _15355_/X sky130_fd_sc_hd__clkbuf_2
X_12567_ _20891_/Q vssd1 vssd1 vccd1 vccd1 _17169_/A sky130_fd_sc_hd__clkbuf_4
XPHY_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14306_ _15574_/C vssd1 vssd1 vccd1 vccd1 _14792_/A sky130_fd_sc_hd__inv_2
XFILLER_8_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11518_ _11518_/A vssd1 vssd1 vccd1 vccd1 _21146_/D sky130_fd_sc_hd__inv_2
X_18074_ _18667_/X _18048_/X _18624_/X _18065_/X vssd1 vssd1 vccd1 vccd1 _18074_/X
+ sky130_fd_sc_hd__o22a_1
X_15286_ _15232_/X _15250_/X _15285_/X _20043_/Q _15160_/X vssd1 vssd1 vccd1 vccd1
+ _20043_/D sky130_fd_sc_hd__a32o_1
X_12498_ _16689_/A vssd1 vssd1 vccd1 vccd1 _12498_/Y sky130_fd_sc_hd__inv_2
XFILLER_144_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17025_ _17025_/A _17026_/B vssd1 vssd1 vccd1 vccd1 _20011_/D sky130_fd_sc_hd__nor2_1
XFILLER_236_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14237_ _19897_/Q _14237_/B vssd1 vssd1 vccd1 vccd1 _14238_/B sky130_fd_sc_hd__or2_1
X_11449_ _21161_/Q _11449_/B vssd1 vssd1 vccd1 vccd1 _11450_/B sky130_fd_sc_hd__or2_1
XFILLER_172_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14168_ _20561_/Q _14101_/Y _20554_/Q _14093_/A vssd1 vssd1 vccd1 vccd1 _14168_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_124_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13119_ _20627_/Q _13112_/X _12993_/X _13115_/X vssd1 vssd1 vccd1 vccd1 _20627_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_3_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18976_ _10843_/X _18281_/S _18976_/S vssd1 vssd1 vccd1 vccd1 _18976_/X sky130_fd_sc_hd__mux2_1
X_14099_ _14099_/A _14099_/B vssd1 vssd1 vccd1 vccd1 _14100_/A sky130_fd_sc_hd__or2_1
XFILLER_67_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20729__RESET_B repeater257/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17927_ _18020_/A vssd1 vssd1 vccd1 vccd1 _17927_/X sky130_fd_sc_hd__buf_1
XFILLER_38_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17858_ _17869_/A vssd1 vssd1 vccd1 vccd1 _17858_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__15245__A1 _20481_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18078__B _18078_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16809_ _16813_/B vssd1 vssd1 vccd1 vccd1 _16815_/B sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_139_HCLK_A clkbuf_4_3_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13256__A0 _13254_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18793__S _18928_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17789_ _21134_/Q vssd1 vssd1 vccd1 vccd1 _17789_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19528_ _19784_/CLK _19528_/D vssd1 vssd1 vccd1 vccd1 _19528_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__18195__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13008__B1 _13006_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19459_ _20136_/CLK _19459_/D vssd1 vssd1 vccd1 vccd1 _19459_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21421_ _21421_/CLK _21421_/D repeater214/X vssd1 vssd1 vccd1 vccd1 _21421_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_147_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21352_ _21407_/CLK _21352_/D repeater252/X vssd1 vssd1 vccd1 vccd1 _21352_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__21170__RESET_B repeater216/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20303_ _20693_/CLK _20303_/D repeater196/X vssd1 vssd1 vccd1 vccd1 _20303_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_190_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21283_ _21342_/CLK _21283_/D repeater211/X vssd1 vssd1 vccd1 vccd1 _21283_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_146_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16342__A _16342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20234_ _21484_/CLK _20234_/D repeater203/X vssd1 vssd1 vccd1 vccd1 _20234_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_150_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17157__B _17169_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11742__B1 _11741_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20165_ _21011_/CLK _20165_/D repeater237/X vssd1 vssd1 vccd1 vccd1 _20165_/Q sky130_fd_sc_hd__dfrtp_1
X_09976_ _09976_/A vssd1 vssd1 vccd1 vccd1 _09976_/X sky130_fd_sc_hd__buf_1
XFILLER_104_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20014__D input71/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20096_ _20101_/CLK _20096_/D repeater259/X vssd1 vssd1 vccd1 vccd1 _20096_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__13495__B1 _13418_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20052__RESET_B repeater281/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13247__B1 _13163_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10820_ _10765_/A _10765_/B _10809_/X _10818_/Y vssd1 vssd1 vccd1 vccd1 _21289_/D
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__18186__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_214_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20998_ _21185_/CLK _20998_/D repeater221/X vssd1 vssd1 vccd1 vccd1 _20998_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_198_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10751_ _16749_/B vssd1 vssd1 vccd1 vccd1 _10752_/B sky130_fd_sc_hd__inv_2
XFILLER_40_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18208__S _18908_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15421__A _15421_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_240_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13470_ _20458_/Q _13466_/X _13282_/X _13467_/X vssd1 vssd1 vccd1 vccd1 _20458_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_231_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10682_ _10661_/A _10661_/B _10677_/X _10679_/Y vssd1 vssd1 vccd1 vccd1 _21332_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_40_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12421_ _12421_/A _12421_/B vssd1 vssd1 vccd1 vccd1 _12461_/A sky130_fd_sc_hd__or2_1
XANTENNA__20253__SET_B repeater217/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15140_ _20459_/Q _15084_/A _15136_/Y _20044_/Q _15139_/X vssd1 vssd1 vccd1 vccd1
+ _15144_/C sky130_fd_sc_hd__o221a_1
X_12352_ _12352_/A vssd1 vssd1 vccd1 vccd1 _12352_/Y sky130_fd_sc_hd__inv_2
XFILLER_181_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11303_ _20916_/Q vssd1 vssd1 vccd1 vccd1 _11315_/A sky130_fd_sc_hd__inv_2
X_15071_ _15071_/A _15195_/A vssd1 vssd1 vccd1 vccd1 _15072_/B sky130_fd_sc_hd__or2_2
XANTENNA__19039__S _19046_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12283_ _20943_/Q vssd1 vssd1 vccd1 vccd1 _12432_/A sky130_fd_sc_hd__inv_2
XFILLER_153_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14022_ _14015_/A _14015_/B _14020_/Y _14004_/X vssd1 vssd1 vccd1 vccd1 _20299_/D
+ sky130_fd_sc_hd__a211oi_2
X_11234_ _21196_/Q vssd1 vssd1 vccd1 vccd1 _11234_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18878__S _18901_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18661__A1 _20361_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18830_ _17349_/Y _17348_/X _18926_/S vssd1 vssd1 vccd1 vccd1 _18830_/X sky130_fd_sc_hd__mux2_1
X_11165_ _11929_/A vssd1 vssd1 vccd1 vccd1 _11165_/X sky130_fd_sc_hd__buf_1
XFILLER_121_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10116_ _10207_/A _20783_/Q _10159_/A _20795_/Q _10115_/X vssd1 vssd1 vccd1 vccd1
+ _10122_/B sky130_fd_sc_hd__o221a_1
XANTENNA_output140_A _21043_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15973_ _16235_/A vssd1 vssd1 vccd1 vccd1 _15973_/X sky130_fd_sc_hd__buf_1
X_18761_ _18760_/X _19231_/X _18930_/S vssd1 vssd1 vccd1 vccd1 _18761_/X sky130_fd_sc_hd__mux2_2
X_11096_ _11096_/A _11096_/B vssd1 vssd1 vccd1 vccd1 _11096_/X sky130_fd_sc_hd__or2_1
XFILLER_209_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17712_ _21078_/Q vssd1 vssd1 vccd1 vccd1 _17712_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17083__A _17083_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14924_ _14923_/Y _20082_/Q _14889_/Y _20102_/Q vssd1 vssd1 vccd1 vccd1 _14924_/X
+ sky130_fd_sc_hd__o22a_1
X_10047_ _21385_/Q vssd1 vssd1 vccd1 vccd1 _10206_/A sky130_fd_sc_hd__inv_2
XFILLER_208_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18692_ _18848_/A0 _14163_/Y _18902_/S vssd1 vssd1 vccd1 vccd1 _18692_/X sky130_fd_sc_hd__mux2_1
XFILLER_236_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17643_ _21049_/Q vssd1 vssd1 vccd1 vccd1 _17643_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13238__B1 _13032_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14855_ _20082_/Q vssd1 vssd1 vccd1 vccd1 _15002_/A sky130_fd_sc_hd__inv_2
XFILLER_17_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13806_ _20603_/Q vssd1 vssd1 vccd1 vccd1 _17542_/A sky130_fd_sc_hd__inv_2
XFILLER_91_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17574_ _17574_/A vssd1 vssd1 vccd1 vccd1 _17907_/A sky130_fd_sc_hd__clkbuf_2
X_14786_ _19126_/X _14280_/X _14293_/X vssd1 vssd1 vccd1 vccd1 _14787_/B sky130_fd_sc_hd__a21oi_1
X_11998_ _20992_/Q _11998_/B vssd1 vssd1 vccd1 vccd1 _11999_/B sky130_fd_sc_hd__or2_1
XFILLER_232_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19313_ _20142_/CLK _19313_/D vssd1 vssd1 vccd1 vccd1 _19313_/Q sky130_fd_sc_hd__dfxtp_1
X_16525_ _16525_/A _16525_/B _16525_/C vssd1 vssd1 vccd1 vccd1 _16525_/X sky130_fd_sc_hd__and3_1
X_13737_ _20185_/Q vssd1 vssd1 vccd1 vccd1 _14575_/B sky130_fd_sc_hd__inv_2
XFILLER_43_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10949_ _10947_/Y _21034_/Q _10948_/Y _21027_/Q vssd1 vssd1 vccd1 vccd1 _10949_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_232_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16456_ _19306_/Q _16452_/X _11502_/X _16454_/X vssd1 vssd1 vccd1 vccd1 _19306_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14738__B1 _13714_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19244_ _17415_/Y _17416_/Y _17417_/Y _17418_/Y _19275_/S0 _21004_/Q vssd1 vssd1
+ vccd1 vccd1 _19244_/X sky130_fd_sc_hd__mux4_2
Xclkbuf_opt_7_HCLK clkbuf_opt_7_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_opt_7_HCLK/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_177_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13668_ _13680_/A vssd1 vssd1 vccd1 vccd1 _13668_/X sky130_fd_sc_hd__buf_1
X_15407_ _19809_/Q _15405_/X _15346_/X _15406_/X vssd1 vssd1 vccd1 vccd1 _19809_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12619_ _12619_/A vssd1 vssd1 vccd1 vccd1 _12619_/X sky130_fd_sc_hd__buf_1
X_19175_ _19302_/Q _19824_/Q _19832_/Q _19416_/Q _19280_/S0 _20122_/Q vssd1 vssd1
+ vccd1 vccd1 _19175_/X sky130_fd_sc_hd__mux4_2
XFILLER_192_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16387_ _19344_/Q _16385_/X _16207_/X _16386_/X vssd1 vssd1 vccd1 vccd1 _19344_/D
+ sky130_fd_sc_hd__a22o_1
X_13599_ _20397_/Q _13594_/X _13454_/X _13595_/X vssd1 vssd1 vccd1 vccd1 _20397_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_118_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18126_ _18125_/X _13908_/Y _18849_/S vssd1 vssd1 vccd1 vccd1 _18126_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15338_ _15345_/A vssd1 vssd1 vccd1 vccd1 _15347_/A sky130_fd_sc_hd__inv_2
XFILLER_145_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18057_ _18298_/X _18048_/X _18361_/X _17996_/X vssd1 vssd1 vccd1 vccd1 _18057_/X
+ sky130_fd_sc_hd__o22a_1
X_15269_ _20480_/Q vssd1 vssd1 vccd1 vccd1 _15269_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20038__SET_B repeater216/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17008_ _17008_/A vssd1 vssd1 vccd1 vccd1 _17008_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18788__S _18910_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09830_ _15876_/A _09827_/X _09828_/X _09829_/X vssd1 vssd1 vccd1 vccd1 _21449_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_113_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09761_ _21236_/Q _09756_/Y _11061_/A _20156_/Q _09760_/X vssd1 vssd1 vccd1 vccd1
+ _09768_/C sky130_fd_sc_hd__o221a_1
X_18959_ _16640_/X _21077_/Q _18962_/S vssd1 vssd1 vccd1 vccd1 _18959_/X sky130_fd_sc_hd__mux2_1
XANTENNA__18404__A1 _20441_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17207__A2 _17205_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09692_ _16338_/A vssd1 vssd1 vccd1 vccd1 _11739_/A sky130_fd_sc_hd__buf_1
XFILLER_55_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20921_ _20930_/CLK _20921_/D repeater266/X vssd1 vssd1 vccd1 vccd1 _20921_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__13229__B1 _13140_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13026__A _13040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20852_ _20857_/CLK _20852_/D repeater243/X vssd1 vssd1 vccd1 vccd1 _20852_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_214_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14441__A2 _20026_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20783_ _21406_/CLK _20783_/D repeater213/X vssd1 vssd1 vccd1 vccd1 _20783_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21351__RESET_B repeater252/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13401__B1 _13280_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21404_ _21405_/CLK _21404_/D repeater252/X vssd1 vssd1 vccd1 vccd1 _21404_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_109_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21335_ _21476_/CLK _21335_/D repeater203/X vssd1 vssd1 vccd1 vccd1 _21335_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_237_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21266_ _21417_/CLK _21266_/D repeater231/X vssd1 vssd1 vccd1 vccd1 _21266_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18698__S _18908_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14304__B _17320_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20217_ _20220_/CLK _20217_/D repeater202/X vssd1 vssd1 vccd1 vccd1 _20217_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_89_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21197_ _21401_/CLK _21197_/D repeater241/X vssd1 vssd1 vccd1 vccd1 _21197_/Q sky130_fd_sc_hd__dfrtp_1
X_20148_ _21239_/CLK _20148_/D repeater250/X vssd1 vssd1 vccd1 vccd1 _20148_/Q sky130_fd_sc_hd__dfrtp_1
X_09959_ _21425_/Q _09957_/X _09688_/X _09958_/X vssd1 vssd1 vccd1 vccd1 _21425_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13468__B1 _13277_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20233__RESET_B repeater203/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20079_ _20107_/CLK _20079_/D repeater259/X vssd1 vssd1 vccd1 vccd1 _20079_/Q sky130_fd_sc_hd__dfrtp_1
X_12970_ _12751_/A _12968_/X _12969_/X vssd1 vssd1 vccd1 vccd1 _12970_/X sky130_fd_sc_hd__o21ba_1
XFILLER_181_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11921_ _16215_/B _15594_/A _11173_/B vssd1 vssd1 vccd1 vccd1 _11921_/X sky130_fd_sc_hd__a21bo_1
XPHY_4510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14640_ _14574_/A _14574_/B _14639_/X _14637_/Y vssd1 vssd1 vccd1 vccd1 _20184_/D
+ sky130_fd_sc_hd__a211oi_2
XPHY_4543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18159__A0 _18848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11852_ _21218_/Q vssd1 vssd1 vccd1 vccd1 _11852_/X sky130_fd_sc_hd__buf_1
XPHY_4554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21439__RESET_B repeater245/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_122_HCLK_A clkbuf_opt_3_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_112_HCLK clkbuf_opt_3_HCLK/A vssd1 vssd1 vccd1 vccd1 _20066_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_4576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10803_ _10775_/A _10775_/B _10795_/X _10801_/Y vssd1 vssd1 vccd1 vccd1 _21299_/D
+ sky130_fd_sc_hd__a211oi_2
XPHY_4587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14571_ _14571_/A _14645_/A vssd1 vssd1 vccd1 vccd1 _14572_/B sky130_fd_sc_hd__or2_2
XPHY_4598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11783_ _21181_/Q _11783_/B _11783_/C _11783_/D vssd1 vssd1 vccd1 vccd1 _11784_/A
+ sky130_fd_sc_hd__or4_4
XPHY_3853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17906__B1 _18434_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16310_ _19382_/Q _16305_/X _16295_/X _16306_/X vssd1 vssd1 vccd1 vccd1 _19382_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_198_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13522_ _13528_/C vssd1 vssd1 vccd1 vccd1 _13530_/B sky130_fd_sc_hd__buf_1
XPHY_3886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21092__RESET_B repeater226/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17290_ _17290_/A vssd1 vssd1 vccd1 vccd1 _17290_/X sky130_fd_sc_hd__clkbuf_2
X_10734_ _19920_/Q _16750_/A _19921_/Q vssd1 vssd1 vccd1 vccd1 _16760_/A sky130_fd_sc_hd__or3_1
XPHY_3897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16241_ _16241_/A vssd1 vssd1 vccd1 vccd1 _16241_/X sky130_fd_sc_hd__buf_1
X_13453_ _20466_/Q _13444_/X _13452_/X _13447_/X vssd1 vssd1 vccd1 vccd1 _20466_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__15393__B1 _15352_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21021__RESET_B repeater238/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10665_ _10665_/A _10672_/A vssd1 vssd1 vccd1 vccd1 _10666_/A sky130_fd_sc_hd__or2_2
X_12404_ _20942_/Q vssd1 vssd1 vccd1 vccd1 _12431_/A sky130_fd_sc_hd__inv_2
X_16172_ _19450_/Q _16166_/X _16139_/X _16168_/X vssd1 vssd1 vccd1 vccd1 _19450_/D
+ sky130_fd_sc_hd__a22o_1
X_13384_ _17177_/A _17169_/C _13384_/C _20872_/Q vssd1 vssd1 vccd1 vccd1 _13601_/B
+ sky130_fd_sc_hd__or4b_4
X_10596_ _20746_/Q vssd1 vssd1 vccd1 vccd1 _10596_/Y sky130_fd_sc_hd__inv_2
XFILLER_166_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15123_ _20459_/Q vssd1 vssd1 vccd1 vccd1 _15123_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12335_ _20981_/Q _12334_/Y _12064_/Y _12334_/A _12206_/X vssd1 vssd1 vccd1 vccd1
+ _20981_/D sky130_fd_sc_hd__o221a_1
XFILLER_5_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15054_ _20048_/Q vssd1 vssd1 vccd1 vccd1 _15128_/A sky130_fd_sc_hd__inv_2
X_19931_ _21238_/CLK _19931_/D repeater251/X vssd1 vssd1 vccd1 vccd1 _19931_/Q sky130_fd_sc_hd__dfrtp_1
X_12266_ _12228_/A _20520_/Q _20919_/Q _12265_/Y vssd1 vssd1 vccd1 vccd1 _12266_/X
+ sky130_fd_sc_hd__o22a_1
X_14005_ _13971_/C _13881_/B _14002_/Y _14004_/X vssd1 vssd1 vccd1 vccd1 _20305_/D
+ sky130_fd_sc_hd__a211oi_2
X_11217_ _21206_/Q _11213_/X _09663_/X _11214_/X vssd1 vssd1 vccd1 vccd1 _21206_/D
+ sky130_fd_sc_hd__a22o_1
X_19862_ _21164_/CLK _19862_/D repeater226/X vssd1 vssd1 vccd1 vccd1 _19862_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17806__A _17806_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12197_ _20976_/Q _12191_/Y _20981_/Q _12194_/Y _12196_/X vssd1 vssd1 vccd1 vccd1
+ _12204_/B sky130_fd_sc_hd__o221a_1
XANTENNA__18401__S _18841_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput81 _17874_/Y vssd1 vssd1 vccd1 vccd1 HRDATA[11] sky130_fd_sc_hd__clkbuf_2
X_18813_ _18812_/X _14568_/A _18898_/S vssd1 vssd1 vccd1 vccd1 _18813_/X sky130_fd_sc_hd__mux2_2
Xoutput92 _17999_/Y vssd1 vssd1 vccd1 vccd1 HRDATA[21] sky130_fd_sc_hd__clkbuf_2
XFILLER_68_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11148_ _11172_/B vssd1 vssd1 vccd1 vccd1 _15594_/A sky130_fd_sc_hd__buf_1
XFILLER_122_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19793_ _19820_/CLK _19793_/D vssd1 vssd1 vccd1 vccd1 _19793_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_233_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18744_ _18743_/X _21348_/Q _18841_/S vssd1 vssd1 vccd1 vccd1 _18744_/X sky130_fd_sc_hd__mux2_2
X_11079_ _11100_/A vssd1 vssd1 vccd1 vccd1 _11079_/X sky130_fd_sc_hd__buf_1
X_15956_ _15962_/A vssd1 vssd1 vccd1 vccd1 _15956_/X sky130_fd_sc_hd__buf_1
XFILLER_64_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14907_ _20589_/Q _20100_/Q _20589_/Q _20100_/Q vssd1 vssd1 vccd1 vccd1 _14907_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_15887_ _16231_/A vssd1 vssd1 vccd1 vccd1 _15887_/X sky130_fd_sc_hd__clkbuf_2
X_18675_ _17773_/X _19340_/Q _18926_/S vssd1 vssd1 vccd1 vccd1 _18675_/X sky130_fd_sc_hd__mux2_1
X_17626_ _19467_/Q vssd1 vssd1 vccd1 vccd1 _17626_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14838_ _14838_/A vssd1 vssd1 vccd1 vccd1 _14960_/B sky130_fd_sc_hd__buf_1
XFILLER_51_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17557_ _17555_/Y _17639_/A _17556_/Y _17381_/X vssd1 vssd1 vccd1 vccd1 _17557_/X
+ sky130_fd_sc_hd__o22a_1
X_14769_ _14769_/A _14769_/B _14769_/C _14769_/D vssd1 vssd1 vccd1 vccd1 _14769_/Y
+ sky130_fd_sc_hd__nor4_2
XFILLER_44_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16508_ _16508_/A vssd1 vssd1 vccd1 vccd1 _16688_/A sky130_fd_sc_hd__buf_1
XFILLER_204_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_44_HCLK_A clkbuf_4_11_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17488_ _19362_/Q vssd1 vssd1 vccd1 vccd1 _17488_/Y sky130_fd_sc_hd__inv_2
XFILLER_176_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19227_ _17509_/Y _17510_/Y _17511_/Y _17512_/Y _20130_/Q _20131_/Q vssd1 vssd1 vccd1
+ vccd1 _19227_/X sky130_fd_sc_hd__mux4_1
X_16439_ _19314_/Q _16434_/X _11504_/X _16436_/X vssd1 vssd1 vccd1 vccd1 _19314_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_176_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18322__A0 _17281_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19158_ _19764_/Q _19756_/Q _19748_/Q _19740_/Q _19285_/S0 _21017_/Q vssd1 vssd1
+ vccd1 vccd1 _19158_/X sky130_fd_sc_hd__mux4_2
XFILLER_9_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18109_ _18109_/A _18109_/B vssd1 vssd1 vccd1 vccd1 _18109_/Y sky130_fd_sc_hd__nor2_8
X_19089_ _21044_/Q _21057_/Q _19872_/Q vssd1 vssd1 vccd1 vccd1 _19089_/X sky130_fd_sc_hd__mux2_1
X_21120_ _21120_/CLK _21120_/D repeater231/X vssd1 vssd1 vccd1 vccd1 _21120_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__13698__B1 _13586_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21051_ _21164_/CLK _21051_/D repeater226/X vssd1 vssd1 vccd1 vccd1 _21051_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__18311__S _18748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20002_ _21055_/CLK _20002_/D repeater220/X vssd1 vssd1 vccd1 vccd1 _20002_/Q sky130_fd_sc_hd__dfrtp_1
X_09813_ _09827_/A vssd1 vssd1 vccd1 vccd1 _09813_/X sky130_fd_sc_hd__buf_1
XFILLER_247_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09744_ _21224_/Q vssd1 vssd1 vccd1 vccd1 _09744_/X sky130_fd_sc_hd__buf_1
XFILLER_74_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18389__A0 _18388_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_135_HCLK clkbuf_4_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20159_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_36_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09675_ _15382_/A vssd1 vssd1 vccd1 vccd1 _12548_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_228_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20904_ _20908_/CLK _20904_/D repeater217/X vssd1 vssd1 vccd1 vccd1 _20904_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_243_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20835_ _20930_/CLK _20835_/D repeater257/X vssd1 vssd1 vccd1 vccd1 _20835_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20766_ _21342_/CLK _20766_/D repeater191/X vssd1 vssd1 vccd1 vccd1 _20766_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20697_ _20697_/CLK _20697_/D repeater193/X vssd1 vssd1 vccd1 vccd1 _20697_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10450_ _20679_/Q vssd1 vssd1 vccd1 vccd1 _10450_/Y sky130_fd_sc_hd__inv_2
XFILLER_164_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18864__A1 _14275_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10381_ _10381_/A vssd1 vssd1 vccd1 vccd1 _10381_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_164_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12120_ _20976_/Q vssd1 vssd1 vccd1 vccd1 _12329_/A sky130_fd_sc_hd__inv_2
X_21318_ _21319_/CLK _21318_/D repeater191/X vssd1 vssd1 vccd1 vccd1 _21318_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_136_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20414__RESET_B repeater186/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13689__B1 _12849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18616__A1 _20767_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12051_ _20383_/Q vssd1 vssd1 vccd1 vccd1 _12051_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21249_ _21431_/CLK _21249_/D repeater237/X vssd1 vssd1 vccd1 vccd1 _21249_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18221__S _18236_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11002_ _11983_/B _19108_/X vssd1 vssd1 vccd1 vccd1 _11012_/B sky130_fd_sc_hd__or2b_1
XFILLER_78_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15810_ _19624_/Q _15807_/X _09835_/X _15808_/X vssd1 vssd1 vccd1 vccd1 _19624_/D
+ sky130_fd_sc_hd__a22o_1
X_16790_ _16790_/A vssd1 vssd1 vccd1 vccd1 _16795_/B sky130_fd_sc_hd__inv_2
XFILLER_19_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14653__A2 _14469_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15741_ _19654_/Q _15736_/X _15706_/X _15737_/X vssd1 vssd1 vccd1 vccd1 _19654_/D
+ sky130_fd_sc_hd__a22o_1
X_12953_ _15382_/A vssd1 vssd1 vccd1 vccd1 _14262_/A sky130_fd_sc_hd__buf_2
XANTENNA__19052__S _19058_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11904_ _19115_/X vssd1 vssd1 vccd1 vccd1 _11913_/A sky130_fd_sc_hd__inv_2
X_18460_ _18459_/X _14580_/A _18898_/S vssd1 vssd1 vccd1 vccd1 _18460_/X sky130_fd_sc_hd__mux2_2
XANTENNA__21273__RESET_B repeater245/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15672_ _21014_/Q vssd1 vssd1 vccd1 vccd1 _16311_/B sky130_fd_sc_hd__buf_1
X_12884_ _13714_/A vssd1 vssd1 vccd1 vccd1 _12884_/X sky130_fd_sc_hd__buf_2
XPHY_4340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14623_ _14623_/A vssd1 vssd1 vccd1 vccd1 _14623_/Y sky130_fd_sc_hd__inv_2
X_17411_ _19361_/Q vssd1 vssd1 vccd1 vccd1 _17411_/Y sky130_fd_sc_hd__inv_2
XPHY_4373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18391_ _18390_/X _15107_/Y _18784_/S vssd1 vssd1 vccd1 vccd1 _18391_/X sky130_fd_sc_hd__mux2_2
X_11835_ _11829_/B _11827_/X _11833_/Y _11834_/X _11812_/A vssd1 vssd1 vccd1 vccd1
+ _11836_/A sky130_fd_sc_hd__o32a_1
XPHY_4384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18891__S _18891_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output103_A _18105_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17342_ _19712_/Q vssd1 vssd1 vccd1 vccd1 _17342_/Y sky130_fd_sc_hd__inv_2
XFILLER_214_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14554_ _20131_/Q _14553_/A _14751_/A _14553_/Y vssd1 vssd1 vccd1 vccd1 _14769_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_198_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11766_ _19083_/X _11764_/X _21051_/Q _11765_/X vssd1 vssd1 vccd1 vccd1 _21051_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13505_ _13514_/A vssd1 vssd1 vccd1 vccd1 _13505_/X sky130_fd_sc_hd__buf_1
X_17273_ _16511_/Y _16688_/A _16501_/X _16505_/X vssd1 vssd1 vccd1 vccd1 _17273_/X
+ sky130_fd_sc_hd__o31a_1
X_10717_ _10704_/A _10704_/B _10715_/Y _10677_/X vssd1 vssd1 vccd1 vccd1 _21316_/D
+ sky130_fd_sc_hd__a211oi_2
XPHY_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14485_ _14461_/A _14370_/B _14483_/Y _14474_/X vssd1 vssd1 vccd1 vccd1 _20227_/D
+ sky130_fd_sc_hd__a211oi_2
XPHY_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11697_ _11704_/A vssd1 vssd1 vccd1 vccd1 _11697_/X sky130_fd_sc_hd__buf_1
XFILLER_158_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_repeater253_A repeater255/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19012_ _16943_/Y _20411_/Q _19019_/S vssd1 vssd1 vccd1 vccd1 _19964_/D sky130_fd_sc_hd__mux2_1
X_16224_ _16224_/A vssd1 vssd1 vccd1 vccd1 _16224_/X sky130_fd_sc_hd__buf_1
XFILLER_201_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13436_ _13444_/A vssd1 vssd1 vccd1 vccd1 _13436_/X sky130_fd_sc_hd__buf_1
X_10648_ _10575_/C _10668_/B _10575_/A vssd1 vssd1 vccd1 vccd1 _10649_/C sky130_fd_sc_hd__o21a_1
XFILLER_167_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_16_HCLK clkbuf_4_3_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19820_/CLK sky130_fd_sc_hd__clkbuf_16
Xrebuffer3 _20027_/Q vssd1 vssd1 vccd1 vccd1 _14425_/B2 sky130_fd_sc_hd__dlygate4sd1_1
XANTENNA_clkbuf_1_0_0_HCLK_A clkbuf_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16155_ _19460_/Q _16151_/X _16135_/X _16153_/X vssd1 vssd1 vccd1 vccd1 _19460_/D
+ sky130_fd_sc_hd__a22o_1
X_13367_ _20509_/Q _13365_/X _13151_/X _13366_/X vssd1 vssd1 vccd1 vccd1 _20509_/D
+ sky130_fd_sc_hd__a22o_1
X_10579_ _10702_/A _20742_/Q _10656_/A _20755_/Q vssd1 vssd1 vccd1 vccd1 _10579_/Y
+ sky130_fd_sc_hd__a22oi_1
X_15106_ _15102_/Y _20071_/Q _20447_/Q _15099_/X _15105_/Y vssd1 vssd1 vccd1 vccd1
+ _15106_/X sky130_fd_sc_hd__o221a_1
XFILLER_127_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12318_ _12318_/A _12366_/A vssd1 vssd1 vccd1 vccd1 _12319_/B sky130_fd_sc_hd__or2_2
X_16086_ _19490_/Q _16080_/X _15873_/X _16082_/X vssd1 vssd1 vccd1 vccd1 _19490_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_5_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13298_ _20546_/Q _13293_/X _13223_/X _13294_/X vssd1 vssd1 vccd1 vccd1 _20546_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_244_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19914_ _21167_/CLK _19914_/D repeater219/X vssd1 vssd1 vccd1 vccd1 _19914_/Q sky130_fd_sc_hd__dfrtp_1
X_15037_ _20065_/Q vssd1 vssd1 vccd1 vccd1 _15079_/A sky130_fd_sc_hd__inv_2
X_12249_ _20918_/Q vssd1 vssd1 vccd1 vccd1 _12468_/A sky130_fd_sc_hd__inv_2
XANTENNA__18131__S _18896_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_158_HCLK clkbuf_opt_1_HCLK/A vssd1 vssd1 vccd1 vccd1 _19834_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_68_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19845_ _21184_/CLK _19845_/D repeater219/X vssd1 vssd1 vccd1 vccd1 _19845_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_150_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19776_ _19776_/CLK _19776_/D vssd1 vssd1 vccd1 vccd1 _19776_/Q sky130_fd_sc_hd__dfxtp_1
X_16988_ _16992_/B vssd1 vssd1 vccd1 vccd1 _16994_/B sky130_fd_sc_hd__inv_2
XFILLER_96_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18727_ _18726_/X _14942_/Y _18907_/S vssd1 vssd1 vccd1 vccd1 _18727_/X sky130_fd_sc_hd__mux2_1
XFILLER_83_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15939_ _19564_/Q _15935_/X _15891_/X _15937_/X vssd1 vssd1 vccd1 vccd1 _19564_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_225_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18658_ _18657_/X _20205_/Q _18748_/S vssd1 vssd1 vccd1 vccd1 _18658_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17609_ _17774_/B vssd1 vssd1 vccd1 vccd1 _17703_/B sky130_fd_sc_hd__buf_1
XFILLER_91_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18589_ _18588_/X _12186_/Y _18787_/S vssd1 vssd1 vccd1 vccd1 _18589_/X sky130_fd_sc_hd__mux2_2
XFILLER_40_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20620_ _20622_/CLK _20620_/D repeater195/X vssd1 vssd1 vccd1 vccd1 _20620_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_20_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20551_ _20947_/CLK _20551_/D repeater258/X vssd1 vssd1 vccd1 vccd1 _20551_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_177_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18306__S _18884_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20482_ _20944_/CLK _20482_/D repeater274/X vssd1 vssd1 vccd1 vccd1 _20482_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__19194__S1 _20122_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14135__A _20550_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21103_ _21429_/CLK _21103_/D repeater229/X vssd1 vssd1 vccd1 vccd1 _21103_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_154_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21034_ _21207_/CLK _21034_/D repeater242/X vssd1 vssd1 vccd1 vccd1 _21034_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_99_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19550__CLK _19706_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09727_ _20158_/Q vssd1 vssd1 vccd1 vccd1 _09727_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09658_ input39/X vssd1 vssd1 vccd1 vccd1 _12863_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_27_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17585__A1 _12605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_243_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11620_ _21109_/Q vssd1 vssd1 vccd1 vccd1 _14813_/B sky130_fd_sc_hd__clkbuf_2
XPHY_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20818_ _21379_/CLK _20818_/D repeater211/X vssd1 vssd1 vccd1 vccd1 _20818_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_39_HCLK _20004_/CLK vssd1 vssd1 vccd1 vccd1 _21184_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_144_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11551_ _17301_/A _14273_/D vssd1 vssd1 vccd1 vccd1 _11562_/A sky130_fd_sc_hd__or2_2
XANTENNA__15348__B1 _15346_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20749_ _21306_/CLK _20749_/D repeater207/X vssd1 vssd1 vccd1 vccd1 _20749_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17888__A2 _17200_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20666__RESET_B repeater207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18216__S _18904_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10502_ _21281_/Q _17544_/A _10757_/A _20669_/Q _10501_/X vssd1 vssd1 vccd1 vccd1
+ _10522_/A sky130_fd_sc_hd__o221a_1
XPHY_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_90_HCLK_A clkbuf_4_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14270_ _20246_/Q _14267_/X _13710_/X _14268_/X vssd1 vssd1 vccd1 vccd1 _20246_/D
+ sky130_fd_sc_hd__a22o_1
X_11482_ _19103_/X _11480_/X _21155_/Q _11481_/X vssd1 vssd1 vccd1 vccd1 _21155_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13221_ input46/X vssd1 vssd1 vccd1 vccd1 _13221_/X sky130_fd_sc_hd__clkbuf_2
X_10433_ _21295_/Q _10428_/Y _10776_/A _20689_/Q _10432_/X vssd1 vssd1 vccd1 vccd1
+ _10446_/B sky130_fd_sc_hd__o221a_1
XANTENNA__19185__S1 _20122_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input64_A HWDATA[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13152_ _13167_/A vssd1 vssd1 vccd1 vccd1 _13152_/X sky130_fd_sc_hd__buf_1
X_10364_ _10381_/A vssd1 vssd1 vccd1 vccd1 _10364_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_98_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12103_ _12103_/A _12103_/B _12103_/C _12102_/X vssd1 vssd1 vccd1 vccd1 _12103_/X
+ sky130_fd_sc_hd__or4b_4
XANTENNA__19047__S _19058_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17960_ _18045_/A vssd1 vssd1 vccd1 vccd1 _17960_/X sky130_fd_sc_hd__buf_1
X_13083_ _20648_/Q _13079_/X _12853_/X _13081_/X vssd1 vssd1 vccd1 vccd1 _20648_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_78_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10295_ _20721_/Q vssd1 vssd1 vccd1 vccd1 _10295_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12034_ _19082_/X _12029_/X _20983_/Q _12030_/X vssd1 vssd1 vccd1 vccd1 _20983_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_151_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16911_ _16914_/B _16910_/Y _16898_/X vssd1 vssd1 vccd1 vccd1 _16911_/X sky130_fd_sc_hd__o21a_1
XFILLER_239_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17891_ _18454_/X _17861_/X _18437_/X _17862_/X _17890_/X vssd1 vssd1 vccd1 vccd1
+ _17891_/X sky130_fd_sc_hd__o221a_4
XANTENNA__18886__S _18886_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19630_ _19821_/CLK _19630_/D vssd1 vssd1 vccd1 vccd1 _19630_/Q sky130_fd_sc_hd__dfxtp_1
X_16842_ _19940_/Q vssd1 vssd1 vccd1 vccd1 _16842_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__21454__RESET_B repeater245/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13108__B _13108_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19561_ _19828_/CLK _19561_/D vssd1 vssd1 vccd1 vccd1 _19561_/Q sky130_fd_sc_hd__dfxtp_1
X_16773_ _16773_/A vssd1 vssd1 vccd1 vccd1 _16778_/B sky130_fd_sc_hd__inv_2
X_13985_ _13891_/A _13891_/B _13983_/Y _14037_/C vssd1 vssd1 vccd1 vccd1 _20315_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_207_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18512_ _18511_/X _17001_/Y _18875_/S vssd1 vssd1 vccd1 vccd1 _18512_/X sky130_fd_sc_hd__mux2_1
XFILLER_207_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15724_ input67/X vssd1 vssd1 vccd1 vccd1 _16231_/A sky130_fd_sc_hd__buf_2
X_12936_ _12936_/A vssd1 vssd1 vccd1 vccd1 _12961_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_34_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19492_ _21040_/CLK _19492_/D vssd1 vssd1 vccd1 vccd1 _19492_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09602__A _20891_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18443_ _18442_/X _17920_/Y _18787_/S vssd1 vssd1 vccd1 vccd1 _18443_/X sky130_fd_sc_hd__mux2_2
XFILLER_233_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12867_ _12874_/A vssd1 vssd1 vccd1 vccd1 _12867_/X sky130_fd_sc_hd__buf_1
XANTENNA__15587__B1 _15585_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15655_ _15722_/A _15655_/B _15722_/C vssd1 vssd1 vccd1 vccd1 _15666_/A sky130_fd_sc_hd__or3_4
XPHY_4170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14606_ _20203_/Q _14605_/Y _14599_/X _14593_/B vssd1 vssd1 vccd1 vccd1 _20203_/D
+ sky130_fd_sc_hd__o211a_1
X_11818_ _11815_/X _11816_/Y _11817_/X vssd1 vssd1 vccd1 vccd1 _11818_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__18525__A0 _17079_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15586_ _15586_/A vssd1 vssd1 vccd1 vccd1 _15586_/X sky130_fd_sc_hd__buf_1
X_18374_ _18373_/X _20520_/Q _18910_/S vssd1 vssd1 vccd1 vccd1 _18374_/X sky130_fd_sc_hd__mux2_1
X_12798_ _12804_/A vssd1 vssd1 vccd1 vccd1 _12798_/X sky130_fd_sc_hd__buf_1
XPHY_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14537_ _20135_/Q vssd1 vssd1 vccd1 vccd1 _15815_/A sky130_fd_sc_hd__inv_2
X_17325_ _18021_/A vssd1 vssd1 vccd1 vccd1 _17928_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_239_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11749_ _11749_/A vssd1 vssd1 vccd1 vccd1 _11749_/Y sky130_fd_sc_hd__inv_2
XFILLER_175_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18126__S _18849_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14468_ _20236_/Q _14380_/C _14410_/Y _14379_/A _14458_/X vssd1 vssd1 vccd1 vccd1
+ _20236_/D sky130_fd_sc_hd__o221a_1
X_17256_ _19599_/Q _17533_/B vssd1 vssd1 vccd1 vccd1 _17256_/Y sky130_fd_sc_hd__nand2_1
XFILLER_174_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16207_ _21449_/Q vssd1 vssd1 vccd1 vccd1 _16207_/X sky130_fd_sc_hd__buf_1
XANTENNA__19176__S1 _20124_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13419_ _13419_/A vssd1 vssd1 vccd1 vccd1 _13447_/A sky130_fd_sc_hd__clkbuf_2
X_17187_ _20737_/Q _17187_/B vssd1 vssd1 vccd1 vccd1 _17187_/Y sky130_fd_sc_hd__nor2_1
X_14399_ _14395_/Y _20225_/Q _14396_/Y _20219_/Q _14398_/X vssd1 vssd1 vccd1 vccd1
+ _14401_/C sky130_fd_sc_hd__a221o_1
XFILLER_127_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12573__B1 _18241_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16138_ _19467_/Q _16130_/X _16137_/X _16133_/X vssd1 vssd1 vccd1 vccd1 _19467_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_170_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15511__B1 _15454_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16069_ _19499_/Q _16064_/X _15764_/X _16066_/X vssd1 vssd1 vccd1 vccd1 _19499_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18796__S _18926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19828_ _19828_/CLK _19828_/D vssd1 vssd1 vccd1 vccd1 _19828_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10887__B1 _10886_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21195__RESET_B repeater220/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17803__A2 _17856_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19759_ _19765_/CLK _19759_/D vssd1 vssd1 vccd1 vccd1 _19759_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__21124__RESET_B repeater190/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17016__B1 _16984_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_240_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13034__A _13040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14250__B1 _19907_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20603_ _20622_/CLK _20603_/D repeater195/X vssd1 vssd1 vccd1 vccd1 _20603_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_149_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20534_ _20947_/CLK _20534_/D repeater265/X vssd1 vssd1 vccd1 vccd1 _20534_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_137_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20077__RESET_B repeater259/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11489__A _13383_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19167__S1 _20122_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_229_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20465_ _20937_/CLK _20465_/D repeater277/X vssd1 vssd1 vccd1 vccd1 _20465_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_193_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20396_ _20930_/CLK _20396_/D repeater268/X vssd1 vssd1 vccd1 vccd1 _20396_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_106_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10590__A2 _20755_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10080_ _20800_/Q vssd1 vssd1 vccd1 vccd1 _10080_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13209__A input52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21017_ _21431_/CLK _21017_/D repeater238/X vssd1 vssd1 vccd1 vccd1 _21017_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_181_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_247_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15424__A _15424_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19942__RESET_B repeater251/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13770_ _20625_/Q vssd1 vssd1 vccd1 vccd1 _13770_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13292__A1 _20550_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10982_ _11883_/A vssd1 vssd1 vccd1 vccd1 _10983_/A sky130_fd_sc_hd__inv_2
XFILLER_55_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12721_ _17549_/A vssd1 vssd1 vccd1 vccd1 _17378_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15440_ _19794_/Q _15434_/X _15421_/X _15436_/X vssd1 vssd1 vccd1 vccd1 _19794_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12652_ _12685_/A vssd1 vssd1 vccd1 vccd1 _12687_/A sky130_fd_sc_hd__inv_2
XPHY_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11603_ _18988_/X _11598_/X _21118_/Q _11600_/X vssd1 vssd1 vccd1 vccd1 _21118_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15371_ _19822_/Q _15366_/X _15355_/X _15367_/X vssd1 vssd1 vccd1 vccd1 _19822_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12583_ _12601_/A vssd1 vssd1 vccd1 vccd1 _12583_/X sky130_fd_sc_hd__buf_1
XPHY_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14322_ _16034_/A _14318_/X _16034_/A _14318_/A vssd1 vssd1 vccd1 vccd1 _14322_/X
+ sky130_fd_sc_hd__o2bb2a_1
XPHY_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17110_ _19582_/Q vssd1 vssd1 vccd1 vccd1 _17110_/Y sky130_fd_sc_hd__inv_2
XPHY_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11534_ _11534_/A vssd1 vssd1 vccd1 vccd1 _11534_/X sky130_fd_sc_hd__buf_1
XPHY_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18090_ _18090_/A _18090_/B _18090_/C _18090_/D vssd1 vssd1 vccd1 vccd1 _18090_/X
+ sky130_fd_sc_hd__or4_4
XPHY_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17041_ _21413_/Q _11617_/X _17040_/Y _14813_/B _11621_/A vssd1 vssd1 vccd1 vccd1
+ _18984_/S sky130_fd_sc_hd__a221oi_2
XPHY_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14253_ _20253_/Q _14246_/A _19905_/Q _14249_/X vssd1 vssd1 vccd1 vccd1 _20253_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19158__S1 _21017_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11465_ _19092_/X _11461_/X _21166_/Q _11463_/X vssd1 vssd1 vccd1 vccd1 _21166_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_139_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12555__B1 _11736_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13204_ _20590_/Q _13200_/X _13001_/X _13201_/X vssd1 vssd1 vccd1 vccd1 _20590_/D
+ sky130_fd_sc_hd__a22o_1
X_10416_ _21347_/Q _10415_/Y _10381_/A _10264_/B vssd1 vssd1 vccd1 vccd1 _21347_/D
+ sky130_fd_sc_hd__o211a_1
X_14184_ _20286_/Q _14182_/Y _14183_/X _14097_/B vssd1 vssd1 vccd1 vccd1 _20286_/D
+ sky130_fd_sc_hd__o211a_1
X_11396_ _16632_/C _11782_/B _11376_/X _11393_/Y _11395_/Y vssd1 vssd1 vccd1 vccd1
+ _11396_/X sky130_fd_sc_hd__a41o_1
XFILLER_180_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13135_ _20617_/Q _13132_/X _12928_/X _13133_/X vssd1 vssd1 vccd1 vccd1 _20617_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_140_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10347_ _20704_/Q vssd1 vssd1 vccd1 vccd1 _10347_/Y sky130_fd_sc_hd__inv_2
XFILLER_151_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18992_ _21261_/Q _21113_/Q _18992_/S vssd1 vssd1 vccd1 vccd1 _18992_/X sky130_fd_sc_hd__mux2_1
XFILLER_155_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17943_ _17943_/A _17943_/B vssd1 vssd1 vccd1 vccd1 _17943_/Y sky130_fd_sc_hd__nor2_1
X_13066_ _13072_/A vssd1 vssd1 vccd1 vccd1 _13066_/X sky130_fd_sc_hd__buf_1
XANTENNA__12858__A1 _20750_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10278_ _10278_/A _10388_/A vssd1 vssd1 vccd1 vccd1 _10279_/B sky130_fd_sc_hd__or2_1
X_12017_ _12029_/A vssd1 vssd1 vccd1 vccd1 _12017_/X sky130_fd_sc_hd__buf_1
Xrepeater207 repeater208/X vssd1 vssd1 vccd1 vccd1 repeater207/X sky130_fd_sc_hd__buf_8
XANTENNA__10869__B1 _09682_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater218 repeater220/X vssd1 vssd1 vccd1 vccd1 repeater218/X sky130_fd_sc_hd__buf_6
XFILLER_39_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17874_ _17852_/X _17868_/X _17871_/X _17873_/X vssd1 vssd1 vccd1 vccd1 _17874_/Y
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__11530__A1 _21143_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater229 repeater230/X vssd1 vssd1 vccd1 vccd1 repeater229/X sky130_fd_sc_hd__clkbuf_8
XFILLER_66_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19613_ _21040_/CLK _19613_/D vssd1 vssd1 vccd1 vccd1 _19613_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16825_ _16830_/B _16824_/X _16803_/X vssd1 vssd1 vccd1 vccd1 _16825_/X sky130_fd_sc_hd__o21a_1
XFILLER_120_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15334__A _15574_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19544_ _19784_/CLK _19544_/D vssd1 vssd1 vccd1 vccd1 _19544_/Q sky130_fd_sc_hd__dfxtp_1
X_16756_ _16756_/A vssd1 vssd1 vccd1 vccd1 _16756_/Y sky130_fd_sc_hd__inv_2
X_13968_ _13897_/A _13897_/B _13898_/Y _14037_/C vssd1 vssd1 vccd1 vccd1 _20321_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_207_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15707_ _19670_/Q _15696_/X _15706_/X _15698_/X vssd1 vssd1 vccd1 vccd1 _19670_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_222_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12919_ _20725_/Q _12915_/X _12918_/X _12916_/X vssd1 vssd1 vccd1 vccd1 _20725_/D
+ sky130_fd_sc_hd__a22o_1
X_19475_ _20432_/CLK _19475_/D vssd1 vssd1 vccd1 vccd1 _19475_/Q sky130_fd_sc_hd__dfxtp_1
X_16687_ _16498_/Y _16686_/Y _16684_/A vssd1 vssd1 vccd1 vccd1 _19872_/D sky130_fd_sc_hd__o21a_1
X_13899_ _20322_/Q vssd1 vssd1 vccd1 vccd1 _13899_/Y sky130_fd_sc_hd__inv_2
X_18426_ _17830_/X _10965_/Y _18928_/S vssd1 vssd1 vccd1 vccd1 _18426_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15638_ _15638_/A _21219_/Q _15638_/C vssd1 vssd1 vccd1 vccd1 _16465_/C sky130_fd_sc_hd__or3_4
XFILLER_210_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13789__A _20614_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18357_ _18356_/X _14092_/A _18850_/S vssd1 vssd1 vccd1 vccd1 _18357_/X sky130_fd_sc_hd__mux2_1
XFILLER_203_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12693__A _12707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15569_ _15569_/A vssd1 vssd1 vccd1 vccd1 _15569_/X sky130_fd_sc_hd__buf_1
XFILLER_187_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12794__B1 _09659_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17308_ _17303_/Y _17376_/A _17304_/Y _17150_/X _17307_/X vssd1 vssd1 vccd1 vccd1
+ _17308_/X sky130_fd_sc_hd__o221a_1
XFILLER_159_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19939__CLK _20930_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18288_ _17813_/Y _16781_/Y _18667_/S vssd1 vssd1 vccd1 vccd1 _18288_/X sky130_fd_sc_hd__mux2_1
XANTENNA__20170__RESET_B repeater233/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19149__S1 _21017_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17239_ _19471_/Q vssd1 vssd1 vccd1 vccd1 _17239_/Y sky130_fd_sc_hd__inv_2
XFILLER_162_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20250_ _21421_/CLK _20250_/D repeater214/X vssd1 vssd1 vccd1 vccd1 _20250_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_127_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20181_ _21483_/CLK _20181_/D repeater200/X vssd1 vssd1 vccd1 vccd1 _20181_/Q sky130_fd_sc_hd__dfrtp_1
X_09992_ _20021_/Q _09986_/B _09987_/A vssd1 vssd1 vccd1 vccd1 _17037_/A sky130_fd_sc_hd__o21ai_1
XFILLER_143_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17724__A _21142_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17788__A1 _16495_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_2_3_0_HCLK_A clkbuf_2_3_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12482__C1 _12445_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_231_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09650__B1 _09649_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20517_ _20944_/CLK _20517_/D repeater277/X vssd1 vssd1 vccd1 vccd1 _20517_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_165_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11250_ _11250_/A vssd1 vssd1 vccd1 vccd1 _11250_/X sky130_fd_sc_hd__buf_1
XFILLER_165_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20448_ _20480_/CLK _20448_/D repeater183/X vssd1 vssd1 vccd1 vccd1 _20448_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_162_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10201_ _10201_/A _10218_/A vssd1 vssd1 vccd1 vccd1 _10216_/A sky130_fd_sc_hd__or2_1
XANTENNA__17476__B1 _18768_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11181_ _11190_/A vssd1 vssd1 vccd1 vccd1 _15885_/A sky130_fd_sc_hd__buf_1
X_20379_ _20957_/CLK _20379_/D repeater186/X vssd1 vssd1 vccd1 vccd1 _20379_/Q sky130_fd_sc_hd__dfrtp_4
X_10132_ _20786_/Q vssd1 vssd1 vccd1 vccd1 _10132_/Y sky130_fd_sc_hd__inv_2
XFILLER_133_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__21046__RESET_B repeater226/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_9_HCLK_A clkbuf_opt_2_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14940_ _14938_/Y _20079_/Q _14939_/Y _20094_/Q vssd1 vssd1 vccd1 vccd1 _14940_/X
+ sky130_fd_sc_hd__o22a_1
X_10063_ _21394_/Q vssd1 vssd1 vccd1 vccd1 _10155_/A sky130_fd_sc_hd__inv_2
XFILLER_248_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_248_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_236_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input27_A HADDR[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14871_ _14961_/B _14987_/A vssd1 vssd1 vccd1 vccd1 _14872_/B sky130_fd_sc_hd__or2_2
X_16610_ _19987_/Q vssd1 vssd1 vccd1 vccd1 _16610_/Y sky130_fd_sc_hd__inv_2
X_13822_ _20600_/Q _14567_/A _20626_/Q _14592_/A vssd1 vssd1 vccd1 vccd1 _13822_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__18728__A0 _17079_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17590_ _19699_/Q vssd1 vssd1 vccd1 vccd1 _17590_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16541_ _16541_/A _16556_/A _16561_/A vssd1 vssd1 vccd1 vccd1 _16541_/X sky130_fd_sc_hd__or3_4
XFILLER_204_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13753_ _20628_/Q _14594_/A _18032_/A _20200_/Q vssd1 vssd1 vccd1 vccd1 _13753_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_28_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10965_ _21212_/Q vssd1 vssd1 vccd1 vccd1 _10965_/Y sky130_fd_sc_hd__inv_2
XFILLER_141_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19060__S _19910_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12704_ _20817_/Q _12701_/X _12548_/X _12702_/X vssd1 vssd1 vccd1 vccd1 _20817_/D
+ sky130_fd_sc_hd__a22o_1
X_19260_ _17269_/Y _17270_/Y _17271_/Y _17272_/Y _20130_/Q _20131_/Q vssd1 vssd1 vccd1
+ vccd1 _19260_/X sky130_fd_sc_hd__mux4_2
X_13684_ _20348_/Q _13679_/X _13489_/X _13680_/X vssd1 vssd1 vccd1 vccd1 _20348_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_44_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16472_ _19296_/Q _16466_/X _16285_/X _16468_/X vssd1 vssd1 vccd1 vccd1 _19296_/D
+ sky130_fd_sc_hd__a22o_1
X_10896_ _11739_/A vssd1 vssd1 vccd1 vccd1 _10896_/X sky130_fd_sc_hd__buf_2
XFILLER_204_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18211_ _18845_/A0 _13818_/Y _18896_/S vssd1 vssd1 vccd1 vccd1 _18211_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12635_ input29/X _12631_/X _20849_/Q _12632_/X vssd1 vssd1 vccd1 vccd1 _20849_/D
+ sky130_fd_sc_hd__o22a_1
XANTENNA__14765__A1 _20132_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15423_ _15423_/A vssd1 vssd1 vccd1 vccd1 _15423_/X sky130_fd_sc_hd__buf_1
X_19191_ _19187_/X _19188_/X _19189_/X _19190_/X _20123_/Q _20124_/Q vssd1 vssd1 vccd1
+ vccd1 _19191_/X sky130_fd_sc_hd__mux4_2
XFILLER_31_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_repeater166_A _18906_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12776__B1 _09628_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18142_ _18845_/A0 _13736_/Y _18896_/S vssd1 vssd1 vccd1 vccd1 _18142_/X sky130_fd_sc_hd__mux2_1
XPHY_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15354_ _15354_/A vssd1 vssd1 vccd1 vccd1 _15592_/A sky130_fd_sc_hd__clkbuf_2
X_12566_ _12574_/A vssd1 vssd1 vccd1 vccd1 _12566_/X sky130_fd_sc_hd__clkbuf_2
XPHY_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11517_ _16711_/A _11497_/A _11514_/Y _11516_/Y _11523_/S vssd1 vssd1 vccd1 vccd1
+ _11518_/A sky130_fd_sc_hd__o32a_1
XPHY_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14305_ _20241_/Q _14730_/B _16479_/A vssd1 vssd1 vccd1 vccd1 _15574_/C sky130_fd_sc_hd__or3_4
XFILLER_172_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15285_ _15259_/X _15285_/B _15285_/C _15285_/D vssd1 vssd1 vccd1 vccd1 _15285_/X
+ sky130_fd_sc_hd__and4b_1
X_18073_ _18408_/X _17858_/X _18515_/X _17211_/X _18072_/X vssd1 vssd1 vccd1 vccd1
+ _18076_/B sky130_fd_sc_hd__o221a_2
XFILLER_157_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18404__S _18906_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12497_ _12490_/A _12490_/B _20918_/Q _12415_/A _12438_/X vssd1 vssd1 vccd1 vccd1
+ _20918_/D sky130_fd_sc_hd__o221a_1
XFILLER_144_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14236_ _19896_/Q _14236_/B vssd1 vssd1 vccd1 vccd1 _14237_/B sky130_fd_sc_hd__or2_1
XANTENNA_output95_A _18042_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17024_ _17024_/A _17026_/B vssd1 vssd1 vccd1 vccd1 _20010_/D sky130_fd_sc_hd__nor2_1
X_11448_ _21160_/Q _11448_/B vssd1 vssd1 vccd1 vccd1 _11449_/B sky130_fd_sc_hd__or2_1
XFILLER_109_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14167_ _20531_/Q vssd1 vssd1 vccd1 vccd1 _14167_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15329__A _15329_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11379_ _11387_/A _11379_/B _11379_/C vssd1 vssd1 vccd1 vccd1 _11385_/D sky130_fd_sc_hd__or3_1
XFILLER_140_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13118_ _20628_/Q _13112_/X _12991_/X _13115_/X vssd1 vssd1 vccd1 vccd1 _20628_/D
+ sky130_fd_sc_hd__a22o_1
X_14098_ _14098_/A _14179_/A vssd1 vssd1 vccd1 vccd1 _14099_/B sky130_fd_sc_hd__or2_1
X_18975_ _16490_/X _16490_/B _18975_/S vssd1 vssd1 vccd1 vccd1 _18975_/X sky130_fd_sc_hd__mux2_1
XANTENNA__19864__RESET_B repeater225/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17926_ _18019_/A vssd1 vssd1 vccd1 vccd1 _17926_/X sky130_fd_sc_hd__buf_1
X_13049_ _13262_/B vssd1 vssd1 vccd1 vccd1 _13259_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11503__A1 _11502_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12700__B1 _12699_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17857_ _17857_/A vssd1 vssd1 vccd1 vccd1 _17857_/X sky130_fd_sc_hd__buf_1
XANTENNA__12688__A _12708_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19611__CLK _21452_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16808_ _19933_/Q vssd1 vssd1 vccd1 vccd1 _16808_/Y sky130_fd_sc_hd__inv_2
XFILLER_226_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18719__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17788_ _16495_/Y _17550_/X _17782_/X _17787_/X vssd1 vssd1 vccd1 vccd1 _17788_/X
+ sky130_fd_sc_hd__o211a_2
X_19527_ _21273_/CLK _19527_/D vssd1 vssd1 vccd1 vccd1 _19527_/Q sky130_fd_sc_hd__dfxtp_1
X_16739_ _19995_/Q _18932_/X _16737_/A _16738_/X vssd1 vssd1 vccd1 vccd1 _16739_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_179_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19458_ _20136_/CLK _19458_/D vssd1 vssd1 vccd1 vccd1 _19458_/Q sky130_fd_sc_hd__dfxtp_1
X_18409_ _17898_/Y _21477_/Q _18669_/S vssd1 vssd1 vccd1 vccd1 _18409_/X sky130_fd_sc_hd__mux2_1
XANTENNA__14756__A1 _20133_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19389_ _20432_/CLK _19389_/D vssd1 vssd1 vccd1 vccd1 _19389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_210_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12767__B1 _12663_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21420_ _21421_/CLK _21420_/D repeater214/X vssd1 vssd1 vccd1 vccd1 _21420_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_194_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21351_ _21407_/CLK _21351_/D repeater252/X vssd1 vssd1 vccd1 vccd1 _21351_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18314__S _18898_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20302_ _20316_/CLK _20302_/D repeater197/X vssd1 vssd1 vccd1 vccd1 _20302_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_135_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21282_ _21342_/CLK _21282_/D repeater207/X vssd1 vssd1 vccd1 vccd1 _21282_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_144_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20233_ _21484_/CLK _20233_/D repeater203/X vssd1 vssd1 vccd1 vccd1 _20233_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_115_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11742__A1 _21057_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09975_ _09975_/A vssd1 vssd1 vccd1 vccd1 _09975_/X sky130_fd_sc_hd__buf_1
X_20164_ _21121_/CLK _20164_/D repeater237/X vssd1 vssd1 vccd1 vccd1 _20164_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17454__A _21083_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09699__B1 _09698_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20095_ _20101_/CLK _20095_/D repeater273/X vssd1 vssd1 vccd1 vccd1 _20095_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_57_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17173__B _17174_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17901__B _17938_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20997_ _21185_/CLK _20997_/D repeater221/X vssd1 vssd1 vccd1 vccd1 _20997_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_53_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10750_ _19949_/Q _19948_/Q _16872_/A vssd1 vssd1 vccd1 vccd1 _16749_/B sky130_fd_sc_hd__or3_4
XFILLER_213_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09700__A input38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10681_ _21333_/Q _10679_/Y _10680_/X _10663_/B vssd1 vssd1 vccd1 vccd1 _21333_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_40_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12420_ _12420_/A _12465_/A vssd1 vssd1 vccd1 vccd1 _12421_/B sky130_fd_sc_hd__or2_2
XANTENNA__19230__S0 _20130_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_224_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12351_ _12119_/X _12327_/B _12350_/X _12347_/Y vssd1 vssd1 vccd1 vccd1 _20974_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_154_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18224__S _18236_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11302_ _11302_/A _12505_/B vssd1 vssd1 vccd1 vccd1 _11315_/C sky130_fd_sc_hd__or2_1
XFILLER_193_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15070_ _15070_/A _15070_/B vssd1 vssd1 vccd1 vccd1 _15195_/A sky130_fd_sc_hd__or2_1
XFILLER_154_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12282_ _12468_/A _20498_/Q _20932_/Q _12274_/Y _12281_/X vssd1 vssd1 vccd1 vccd1
+ _12282_/X sky130_fd_sc_hd__a221o_1
XFILLER_142_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__21227__RESET_B repeater249/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14021_ _20300_/Q _14020_/Y _14017_/B _13988_/X vssd1 vssd1 vccd1 vccd1 _20300_/D
+ sky130_fd_sc_hd__o211a_1
X_11233_ _21195_/Q _11241_/A _11233_/C vssd1 vssd1 vccd1 vccd1 _11235_/A sky130_fd_sc_hd__or3_1
XFILLER_106_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_145_HCLK_A clkbuf_opt_1_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11164_ _16616_/A _16593_/B vssd1 vssd1 vccd1 vccd1 _11929_/A sky130_fd_sc_hd__nand2_1
XFILLER_136_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19055__S _19058_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10115_ _10201_/A _20777_/Q _10034_/A _20801_/Q vssd1 vssd1 vccd1 vccd1 _10115_/X
+ sky130_fd_sc_hd__o22a_1
X_18760_ _18759_/X _17530_/X _18929_/S vssd1 vssd1 vccd1 vccd1 _18760_/X sky130_fd_sc_hd__mux2_1
X_15972_ _19549_/Q _15968_/X _15969_/X _15971_/X vssd1 vssd1 vccd1 vccd1 _19549_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13486__A1 _20451_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11095_ _11095_/A vssd1 vssd1 vccd1 vccd1 _21232_/D sky130_fd_sc_hd__inv_2
XFILLER_103_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17711_ _21062_/Q vssd1 vssd1 vccd1 vccd1 _17711_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14923_ _20571_/Q vssd1 vssd1 vccd1 vccd1 _14923_/Y sky130_fd_sc_hd__inv_2
X_10046_ _10204_/A _10203_/A _10202_/A _10199_/A vssd1 vssd1 vccd1 vccd1 _10053_/C
+ sky130_fd_sc_hd__or4_4
X_18691_ _18690_/X _14572_/A _18898_/S vssd1 vssd1 vccd1 vccd1 _18691_/X sky130_fd_sc_hd__mux2_2
XANTENNA_output133_A _21410_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18894__S _18910_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17642_ _21069_/Q vssd1 vssd1 vccd1 vccd1 _17642_/Y sky130_fd_sc_hd__inv_2
XFILLER_236_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14854_ _20083_/Q vssd1 vssd1 vccd1 vccd1 _15003_/A sky130_fd_sc_hd__inv_2
XFILLER_17_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13805_ _20186_/Q vssd1 vssd1 vccd1 vccd1 _14575_/A sky130_fd_sc_hd__inv_2
XANTENNA__17811__B _17812_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17573_ _17573_/A vssd1 vssd1 vccd1 vccd1 _17574_/A sky130_fd_sc_hd__inv_2
X_11997_ _20991_/Q _11997_/B vssd1 vssd1 vccd1 vccd1 _11998_/B sky130_fd_sc_hd__or2_1
X_14785_ _20124_/Q _14787_/A _14276_/Y _14784_/A vssd1 vssd1 vccd1 vccd1 _20124_/D
+ sky130_fd_sc_hd__o22a_1
X_19312_ _20241_/CLK _19312_/D vssd1 vssd1 vccd1 vccd1 _19312_/Q sky130_fd_sc_hd__dfxtp_1
X_16524_ _16524_/A vssd1 vssd1 vccd1 vccd1 _16524_/Y sky130_fd_sc_hd__inv_2
X_13736_ _20630_/Q vssd1 vssd1 vccd1 vccd1 _13736_/Y sky130_fd_sc_hd__inv_2
X_10948_ _21200_/Q vssd1 vssd1 vccd1 vccd1 _10948_/Y sky130_fd_sc_hd__inv_2
XFILLER_232_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19243_ _17411_/Y _17412_/Y _17413_/Y _17414_/Y _19275_/S0 _21004_/Q vssd1 vssd1
+ vccd1 vccd1 _19243_/X sky130_fd_sc_hd__mux4_1
XANTENNA__09610__A _20872_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16455_ _19307_/Q _16452_/X _11486_/X _16454_/X vssd1 vssd1 vccd1 vccd1 _19307_/D
+ sky130_fd_sc_hd__a22o_1
X_13667_ _13679_/A vssd1 vssd1 vccd1 vccd1 _13667_/X sky130_fd_sc_hd__buf_1
X_10879_ _10888_/A vssd1 vssd1 vccd1 vccd1 _10879_/X sky130_fd_sc_hd__buf_1
XPHY_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15406_ _15406_/A vssd1 vssd1 vccd1 vccd1 _15406_/X sky130_fd_sc_hd__clkbuf_2
X_12618_ input9/X _12613_/X _20860_/Q _12614_/X vssd1 vssd1 vccd1 vccd1 _20860_/D
+ sky130_fd_sc_hd__o22a_1
X_19174_ _19728_/Q _19368_/Q _19784_/Q _19768_/Q _19280_/S0 _20122_/Q vssd1 vssd1
+ vccd1 vccd1 _19174_/X sky130_fd_sc_hd__mux4_1
XPHY_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16386_ _16386_/A vssd1 vssd1 vccd1 vccd1 _16386_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__19221__S0 _20132_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13598_ _20398_/Q _13594_/X _13452_/X _13595_/X vssd1 vssd1 vccd1 vccd1 _20398_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_118_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18125_ _18848_/A0 _14112_/Y _18902_/S vssd1 vssd1 vccd1 vccd1 _18125_/X sky130_fd_sc_hd__mux2_1
XFILLER_247_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12549_ _20899_/Q _12543_/X _12548_/X _12546_/X vssd1 vssd1 vccd1 vccd1 _20899_/D
+ sky130_fd_sc_hd__a22o_1
X_15337_ _15345_/A vssd1 vssd1 vccd1 vccd1 _15337_/X sky130_fd_sc_hd__buf_1
XANTENNA__18134__S _18666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18056_ _18389_/X _18019_/X _18267_/X _18020_/X _18055_/X vssd1 vssd1 vccd1 vccd1
+ _18059_/B sky130_fd_sc_hd__o221a_2
X_15268_ _15265_/Y _20070_/Q _20494_/Q _15087_/A _15267_/X vssd1 vssd1 vccd1 vccd1
+ _15285_/C sky130_fd_sc_hd__o221a_1
XFILLER_126_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13174__B1 _13173_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17007_ _19979_/Q vssd1 vssd1 vccd1 vccd1 _17007_/Y sky130_fd_sc_hd__inv_2
X_14219_ _14219_/A vssd1 vssd1 vccd1 vccd1 _14219_/Y sky130_fd_sc_hd__inv_2
X_15199_ _20055_/Q _15201_/A _15185_/X _15070_/B vssd1 vssd1 vccd1 vccd1 _20055_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__18101__B2 _17861_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12921__B1 _12920_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09760_ _11053_/A _20148_/Q _21228_/Q _09759_/Y vssd1 vssd1 vccd1 vccd1 _09760_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__17860__B1 _18564_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_67_HCLK_A clkbuf_4_11_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18958_ _16642_/X _21078_/Q _18962_/S vssd1 vssd1 vccd1 vccd1 _18958_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17909_ _18420_/X _17954_/A _18410_/X _17572_/B vssd1 vssd1 vccd1 vccd1 _17909_/X
+ sky130_fd_sc_hd__a22o_1
X_09691_ input60/X vssd1 vssd1 vccd1 vccd1 _16338_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_239_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18889_ _18888_/X _17184_/Y _18901_/S vssd1 vssd1 vccd1 vccd1 _18889_/X sky130_fd_sc_hd__mux2_1
XFILLER_227_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20920_ _20930_/CLK _20920_/D repeater268/X vssd1 vssd1 vccd1 vccd1 _20920_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_55_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20851_ _20857_/CLK _20851_/D repeater243/X vssd1 vssd1 vccd1 vccd1 _20851_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18309__S _18896_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12988__B1 _12984_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20782_ _21379_/CLK _20782_/D repeater213/X vssd1 vssd1 vccd1 vccd1 _20782_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_211_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15926__B1 _15785_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19212__S0 _19275_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_72_HCLK clkbuf_opt_7_HCLK/A vssd1 vssd1 vccd1 vccd1 _21485_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_194_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21403_ _21405_/CLK _21403_/D repeater255/X vssd1 vssd1 vccd1 vccd1 _21403_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_157_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12881__A _13171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18340__A1 _20025_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21334_ _21334_/CLK _21334_/D repeater203/X vssd1 vssd1 vccd1 vccd1 _21334_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__21320__RESET_B repeater205/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11497__A _11497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_237_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21265_ _21417_/CLK _21265_/D repeater234/X vssd1 vssd1 vccd1 vccd1 _21265_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_104_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12912__B1 _12666_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20216_ _20220_/CLK _20216_/D repeater202/X vssd1 vssd1 vccd1 vccd1 _20216_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_103_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21196_ _21196_/CLK _21196_/D repeater218/X vssd1 vssd1 vccd1 vccd1 _21196_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_104_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20147_ _21239_/CLK _20147_/D repeater242/X vssd1 vssd1 vccd1 vccd1 _20147_/Q sky130_fd_sc_hd__dfrtp_4
X_09958_ _09958_/A vssd1 vssd1 vccd1 vccd1 _09958_/X sky130_fd_sc_hd__buf_1
XANTENNA__19279__S0 _19280_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20078_ _20107_/CLK _20078_/D repeater259/X vssd1 vssd1 vccd1 vccd1 _20078_/Q sky130_fd_sc_hd__dfrtp_1
X_09889_ _21259_/Q _17026_/A _21259_/Q _17026_/A vssd1 vssd1 vccd1 vccd1 _09916_/A
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__13217__A _13217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11920_ _16465_/B vssd1 vssd1 vccd1 vccd1 _16215_/B sky130_fd_sc_hd__buf_1
XFILLER_246_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20273__RESET_B repeater263/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11851_ _21030_/Q _11851_/B vssd1 vssd1 vccd1 vccd1 _11851_/Y sky130_fd_sc_hd__nor2_1
XPHY_4544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18219__S _18242_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10802_ _21300_/Q _10801_/Y _10798_/X _10777_/B vssd1 vssd1 vccd1 vccd1 _21300_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_32_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14570_ _14570_/A _14570_/B vssd1 vssd1 vccd1 vccd1 _14645_/A sky130_fd_sc_hd__or2_1
X_11782_ _18967_/X _11782_/B vssd1 vssd1 vccd1 vccd1 _16596_/D sky130_fd_sc_hd__nand2_1
XFILLER_214_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_0_0_HCLK clkbuf_4_1_0_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_opt_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XPHY_3865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10733_ _19919_/Q _19918_/Q vssd1 vssd1 vccd1 vccd1 _16750_/A sky130_fd_sc_hd__or2_1
X_13521_ _13521_/A _13520_/Y vssd1 vssd1 vccd1 vccd1 _13528_/C sky130_fd_sc_hd__or2b_1
XPHY_3887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15917__B1 _15916_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16240_ _16240_/A vssd1 vssd1 vccd1 vccd1 _16240_/X sky130_fd_sc_hd__buf_1
X_13452_ _15429_/A vssd1 vssd1 vccd1 vccd1 _13452_/X sky130_fd_sc_hd__buf_2
X_10664_ _10664_/A _10675_/A _10664_/C vssd1 vssd1 vccd1 vccd1 _10672_/A sky130_fd_sc_hd__or3_4
XFILLER_13_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15393__A1 _19815_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19203__S0 _19275_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12403_ _12422_/A _12421_/A _12403_/C _12403_/D vssd1 vssd1 vccd1 vccd1 _12406_/B
+ sky130_fd_sc_hd__or4_4
X_16171_ _19451_/Q _16166_/X _16137_/X _16168_/X vssd1 vssd1 vccd1 vccd1 _19451_/D
+ sky130_fd_sc_hd__a22o_1
X_13383_ _13383_/A vssd1 vssd1 vccd1 vccd1 _17169_/C sky130_fd_sc_hd__buf_1
X_10595_ _10652_/A _20751_/Q _21323_/Q _10592_/Y _10594_/X vssd1 vssd1 vccd1 vccd1
+ _10605_/A sky130_fd_sc_hd__o221a_1
X_12334_ _12334_/A vssd1 vssd1 vccd1 vccd1 _12334_/Y sky130_fd_sc_hd__inv_2
X_15122_ _20463_/Q vssd1 vssd1 vccd1 vccd1 _15122_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18889__S _18901_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13156__B1 _13030_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15053_ _20049_/Q vssd1 vssd1 vccd1 vccd1 _15064_/A sky130_fd_sc_hd__inv_2
X_19930_ _20841_/CLK _19930_/D repeater251/X vssd1 vssd1 vccd1 vccd1 _19930_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_182_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12265_ _20499_/Q vssd1 vssd1 vccd1 vccd1 _12265_/Y sky130_fd_sc_hd__inv_2
XFILLER_126_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14004_ _14004_/A vssd1 vssd1 vccd1 vccd1 _14004_/X sky130_fd_sc_hd__clkbuf_2
X_11216_ _21207_/Q _11213_/X _09659_/X _11214_/X vssd1 vssd1 vccd1 vccd1 _21207_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_3_6_0_HCLK_A clkbuf_3_7_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19861_ _21164_/CLK _19861_/D repeater226/X vssd1 vssd1 vccd1 vccd1 _19861_/Q sky130_fd_sc_hd__dfrtp_1
X_12196_ _12306_/A _20334_/Q _20952_/Q _12195_/Y vssd1 vssd1 vccd1 vccd1 _12196_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__17806__B _17807_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18812_ _18811_/X _14409_/Y _18897_/S vssd1 vssd1 vccd1 vccd1 _18812_/X sky130_fd_sc_hd__mux2_1
Xoutput82 _17883_/Y vssd1 vssd1 vccd1 vccd1 HRDATA[12] sky130_fd_sc_hd__clkbuf_2
Xoutput93 _18014_/X vssd1 vssd1 vccd1 vccd1 HRDATA[22] sky130_fd_sc_hd__clkbuf_2
X_11147_ _15638_/A _15466_/B vssd1 vssd1 vccd1 vccd1 _11172_/B sky130_fd_sc_hd__or2_1
X_19792_ _19820_/CLK _19792_/D vssd1 vssd1 vccd1 vccd1 _19792_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09605__A _17204_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18743_ _17545_/Y _20777_/Q _18885_/S vssd1 vssd1 vccd1 vccd1 _18743_/X sky130_fd_sc_hd__mux2_1
X_15955_ _15961_/A vssd1 vssd1 vccd1 vccd1 _15962_/A sky130_fd_sc_hd__inv_2
X_11078_ _11078_/A vssd1 vssd1 vccd1 vccd1 _21236_/D sky130_fd_sc_hd__inv_2
XFILLER_110_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14906_ _20573_/Q vssd1 vssd1 vccd1 vccd1 _14906_/Y sky130_fd_sc_hd__inv_2
X_10029_ _21406_/Q vssd1 vssd1 vccd1 vccd1 _10077_/A sky130_fd_sc_hd__inv_2
X_18674_ _17774_/X _20151_/Q _18928_/S vssd1 vssd1 vccd1 vccd1 _18674_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15886_ _15896_/A vssd1 vssd1 vccd1 vccd1 _15886_/X sky130_fd_sc_hd__buf_1
XFILLER_236_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17625_ _19459_/Q vssd1 vssd1 vccd1 vccd1 _17625_/Y sky130_fd_sc_hd__inv_2
X_14837_ _20096_/Q vssd1 vssd1 vccd1 vccd1 _14838_/A sky130_fd_sc_hd__inv_2
XANTENNA__17541__B _17542_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18129__S _18909_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17556_ _21048_/Q vssd1 vssd1 vccd1 vccd1 _17556_/Y sky130_fd_sc_hd__inv_2
X_14768_ _14755_/Y _14767_/X _14755_/Y _14767_/X vssd1 vssd1 vccd1 vccd1 _14769_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_32_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_95_HCLK clkbuf_4_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20592_/CLK sky130_fd_sc_hd__clkbuf_16
X_16507_ _16507_/A _16507_/B vssd1 vssd1 vccd1 vccd1 _16508_/A sky130_fd_sc_hd__or2_1
XFILLER_149_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13719_ input73/X _15758_/A _13725_/S vssd1 vssd1 vccd1 vccd1 _20331_/D sky130_fd_sc_hd__mux2_1
X_17487_ _19474_/Q vssd1 vssd1 vccd1 vccd1 _17487_/Y sky130_fd_sc_hd__inv_2
X_14699_ _18244_/X _14696_/X _20161_/Q _14688_/X vssd1 vssd1 vccd1 vccd1 _20161_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_177_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19226_ _19222_/X _19223_/X _19224_/X _19225_/X _21005_/Q _21006_/Q vssd1 vssd1 vccd1
+ vccd1 _19226_/X sky130_fd_sc_hd__mux4_2
XFILLER_176_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16438_ _19315_/Q _16434_/X _11502_/X _16436_/X vssd1 vssd1 vccd1 vccd1 _19315_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_192_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13395__B1 _13270_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19157_ _19684_/Q _19812_/Q _19804_/Q _19796_/Q _19285_/S0 _21017_/Q vssd1 vssd1
+ vccd1 vccd1 _19157_/X sky130_fd_sc_hd__mux4_2
X_16369_ _19353_/Q _16363_/X _16204_/X _16365_/X vssd1 vssd1 vccd1 vccd1 _19353_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_191_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18108_ _17506_/Y _17607_/Y _17423_/Y _17505_/X _18107_/X vssd1 vssd1 vccd1 vccd1
+ _18109_/B sky130_fd_sc_hd__o221a_2
X_19088_ _21045_/Q _21058_/Q _19872_/Q vssd1 vssd1 vccd1 vccd1 _19088_/X sky130_fd_sc_hd__mux2_1
XANTENNA__16333__B1 _16332_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18799__S _18929_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13147__B1 _13146_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_1_HCLK clkbuf_opt_0_HCLK/A vssd1 vssd1 vccd1 vccd1 _19789_/CLK sky130_fd_sc_hd__clkbuf_16
X_18039_ _18365_/X _17907_/A _18354_/X _17908_/A vssd1 vssd1 vccd1 vccd1 _18042_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_114_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21050_ _21164_/CLK _21050_/D repeater227/X vssd1 vssd1 vccd1 vccd1 _21050_/Q sky130_fd_sc_hd__dfrtp_1
X_20001_ _21164_/CLK _20001_/D repeater225/X vssd1 vssd1 vccd1 vccd1 _20001_/Q sky130_fd_sc_hd__dfrtp_1
X_09812_ _09812_/A _09812_/B vssd1 vssd1 vccd1 vccd1 _09827_/A sky130_fd_sc_hd__or2_4
XANTENNA__15517__A input63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20713__RESET_B repeater254/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09743_ _21233_/Q vssd1 vssd1 vccd1 vccd1 _11058_/A sky130_fd_sc_hd__inv_2
XFILLER_223_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09674_ input66/X vssd1 vssd1 vccd1 vccd1 _15382_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_228_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20903_ _21196_/CLK _20903_/D repeater217/X vssd1 vssd1 vccd1 vccd1 _20903_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_215_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20834_ _20930_/CLK _20834_/D repeater268/X vssd1 vssd1 vccd1 vccd1 _20834_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_82_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18010__B1 _18295_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20765_ _21342_/CLK _20765_/D repeater211/X vssd1 vssd1 vccd1 vccd1 _20765_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20696_ _20697_/CLK _20696_/D repeater193/X vssd1 vssd1 vccd1 vccd1 _20696_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_149_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17179__A _17193_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19967__RESET_B repeater184/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18313__A1 _10618_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16324__B1 _16016_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10380_ _10380_/A vssd1 vssd1 vccd1 vccd1 _10380_/Y sky130_fd_sc_hd__inv_2
XFILLER_164_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21317_ _21319_/CLK _21317_/D repeater191/X vssd1 vssd1 vccd1 vccd1 _21317_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_164_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18502__S _18896_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13689__A1 _20347_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12050_ _20969_/Q vssd1 vssd1 vccd1 vccd1 _12322_/A sky130_fd_sc_hd__inv_2
X_21248_ _21431_/CLK _21248_/D repeater237/X vssd1 vssd1 vccd1 vccd1 _21248_/Q sky130_fd_sc_hd__dfstp_4
X_11001_ _10991_/B _15396_/B _21016_/Q _15505_/B vssd1 vssd1 vccd1 vccd1 _11983_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_117_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15427__A _15588_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21179_ _21183_/CLK _21179_/D repeater216/X vssd1 vssd1 vccd1 vccd1 _21179_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_77_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_237_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_50_HCLK_A clkbuf_4_9_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13310__B1 _13154_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15740_ _19655_/Q _15736_/X _15703_/X _15737_/X vssd1 vssd1 vccd1 vccd1 _19655_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_93_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12952_ _20710_/Q _12948_/X _12950_/X _12951_/X vssd1 vssd1 vccd1 vccd1 _20710_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_45_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11903_ _11896_/A _10991_/B _19114_/X _21016_/Q vssd1 vssd1 vccd1 vccd1 _21016_/D
+ sky130_fd_sc_hd__o22a_1
X_15671_ _19686_/Q _15666_/X _15592_/X _15667_/X vssd1 vssd1 vccd1 vccd1 _19686_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12883_ _15354_/A vssd1 vssd1 vccd1 vccd1 _13714_/A sky130_fd_sc_hd__buf_4
XANTENNA__12786__A _12804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17410_ _19473_/Q vssd1 vssd1 vccd1 vccd1 _17410_/Y sky130_fd_sc_hd__inv_2
X_14622_ _14583_/A _14583_/B _14621_/X _14619_/Y vssd1 vssd1 vccd1 vccd1 _20194_/D
+ sky130_fd_sc_hd__a211oi_2
XPHY_4363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18390_ _17079_/Y _15221_/Y _18908_/S vssd1 vssd1 vccd1 vccd1 _18390_/X sky130_fd_sc_hd__mux2_1
X_11834_ _21218_/Q vssd1 vssd1 vccd1 vccd1 _11834_/X sky130_fd_sc_hd__buf_1
XPHY_4374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17341_ _19720_/Q vssd1 vssd1 vccd1 vccd1 _17341_/Y sky130_fd_sc_hd__inv_2
X_11765_ _11771_/A vssd1 vssd1 vccd1 vccd1 _11765_/X sky130_fd_sc_hd__buf_1
XFILLER_186_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14553_ _14553_/A vssd1 vssd1 vccd1 vccd1 _14553_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15312__D _15312_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10716_ _21317_/Q _10715_/Y _10706_/B _10712_/X vssd1 vssd1 vccd1 vccd1 _21317_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13504_ _20441_/Q _13499_/X _13313_/X _13500_/X vssd1 vssd1 vccd1 vccd1 _20441_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_9_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17272_ _19463_/Q vssd1 vssd1 vccd1 vccd1 _17272_/Y sky130_fd_sc_hd__inv_2
XFILLER_201_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14484_ _20228_/Q _14483_/Y _14472_/X _14372_/B vssd1 vssd1 vccd1 vccd1 _20228_/D
+ sky130_fd_sc_hd__o211a_1
X_11696_ _17286_/A _15312_/D vssd1 vssd1 vccd1 vccd1 _11704_/A sky130_fd_sc_hd__or2_2
XPHY_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19011_ _16947_/X _20412_/Q _19019_/S vssd1 vssd1 vccd1 vccd1 _19965_/D sky130_fd_sc_hd__mux2_1
XFILLER_201_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16223_ _16223_/A vssd1 vssd1 vccd1 vccd1 _16223_/X sky130_fd_sc_hd__buf_1
X_10647_ _10647_/A vssd1 vssd1 vccd1 vccd1 _10668_/B sky130_fd_sc_hd__inv_2
X_13435_ _20473_/Q _13428_/X _13313_/X _13430_/X vssd1 vssd1 vccd1 vccd1 _20473_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_173_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_repeater246_A repeater247/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11927__A1 _11916_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrebuffer4 rebuffer6/X vssd1 vssd1 vccd1 vccd1 _14964_/B sky130_fd_sc_hd__dlygate4sd1_1
X_16154_ _19461_/Q _16151_/X _16131_/X _16153_/X vssd1 vssd1 vccd1 vccd1 _19461_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16315__B1 _16231_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13366_ _13378_/A vssd1 vssd1 vccd1 vccd1 _13366_/X sky130_fd_sc_hd__buf_1
X_10578_ _20741_/Q vssd1 vssd1 vccd1 vccd1 _10578_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13129__B1 _12918_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15105_ _15103_/Y _15029_/A _20457_/Q _15104_/X vssd1 vssd1 vccd1 vccd1 _15105_/Y
+ sky130_fd_sc_hd__a22oi_1
X_12317_ _12317_/A _12317_/B vssd1 vssd1 vccd1 vccd1 _12366_/A sky130_fd_sc_hd__or2_1
XFILLER_6_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17817__A _17854_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16085_ _19491_/Q _16080_/X _15871_/X _16082_/X vssd1 vssd1 vccd1 vccd1 _19491_/D
+ sky130_fd_sc_hd__a22o_1
X_13297_ _20547_/Q _13293_/X _13221_/X _13294_/X vssd1 vssd1 vccd1 vccd1 _20547_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18412__S _18849_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19913_ _21055_/CLK _19913_/D repeater220/X vssd1 vssd1 vccd1 vccd1 _19913_/Q sky130_fd_sc_hd__dfrtp_1
X_15036_ _20066_/Q vssd1 vssd1 vccd1 vccd1 _15129_/A sky130_fd_sc_hd__inv_2
X_12248_ _12395_/B _20525_/Q _12396_/B _20500_/Q _12247_/X vssd1 vssd1 vccd1 vccd1
+ _12255_/C sky130_fd_sc_hd__o221a_1
XFILLER_96_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19844_ _21183_/CLK _19844_/D repeater219/X vssd1 vssd1 vccd1 vccd1 _19844_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_229_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12179_ _20345_/Q vssd1 vssd1 vccd1 vccd1 _12179_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20195__RESET_B repeater193/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19775_ _19776_/CLK _19775_/D vssd1 vssd1 vccd1 vccd1 _19775_/Q sky130_fd_sc_hd__dfxtp_1
X_16987_ _19974_/Q _16989_/B vssd1 vssd1 vccd1 vccd1 _16992_/B sky130_fd_sc_hd__or2_1
XFILLER_237_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18726_ _18725_/X _15132_/Y _18784_/S vssd1 vssd1 vccd1 vccd1 _18726_/X sky130_fd_sc_hd__mux2_2
X_15938_ _19565_/Q _15935_/X _15887_/X _15937_/X vssd1 vssd1 vccd1 vccd1 _19565_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_225_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18657_ _18081_/Y _20030_/Q _18669_/S vssd1 vssd1 vccd1 vccd1 _18657_/X sky130_fd_sc_hd__mux2_1
X_15869_ _15869_/A vssd1 vssd1 vccd1 vccd1 _15869_/X sky130_fd_sc_hd__buf_1
XFILLER_36_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17608_ _19603_/Q _17631_/B vssd1 vssd1 vccd1 vccd1 _17608_/X sky130_fd_sc_hd__or2_1
X_18588_ _17079_/Y _12140_/Y _18908_/S vssd1 vssd1 vccd1 vccd1 _18588_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17539_ _17539_/A _17542_/B vssd1 vssd1 vccd1 vccd1 _17539_/Y sky130_fd_sc_hd__nor2_1
X_20550_ _20947_/CLK _20550_/D repeater266/X vssd1 vssd1 vccd1 vccd1 _20550_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_193_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19209_ _17694_/Y _17695_/Y _17696_/Y _17697_/Y _20130_/Q _20131_/Q vssd1 vssd1 vccd1
+ vccd1 _19209_/X sky130_fd_sc_hd__mux4_1
XANTENNA__13368__B1 _13154_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20481_ _20944_/CLK _20481_/D repeater274/X vssd1 vssd1 vccd1 vccd1 _20481_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_145_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20965__RESET_B repeater186/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16631__A _16631_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18322__S _18835_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21102_ _21429_/CLK _21102_/D repeater229/X vssd1 vssd1 vccd1 vccd1 _21102_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_161_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_102_HCLK clkbuf_4_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20101_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_160_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21033_ _21218_/CLK _21033_/D repeater242/X vssd1 vssd1 vccd1 vccd1 _21033_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_219_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input1_A HADDR[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11494__B _17169_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09726_ _21238_/Q vssd1 vssd1 vccd1 vccd1 _11063_/A sky130_fd_sc_hd__inv_2
XFILLER_28_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09657_ _09657_/A vssd1 vssd1 vccd1 vccd1 _09657_/X sky130_fd_sc_hd__buf_1
XFILLER_103_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17585__A2 _17579_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20817_ _21141_/CLK _20817_/D repeater212/X vssd1 vssd1 vccd1 vccd1 _20817_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11550_ _17387_/A vssd1 vssd1 vccd1 vccd1 _17301_/A sky130_fd_sc_hd__buf_1
XPHY_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20748_ _21306_/CLK _20748_/D repeater207/X vssd1 vssd1 vccd1 vccd1 _20748_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10501_ _21289_/Q _10499_/Y _21297_/Q _17981_/A vssd1 vssd1 vccd1 vccd1 _10501_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11481_ _11481_/A vssd1 vssd1 vccd1 vccd1 _11481_/X sky130_fd_sc_hd__buf_1
XPHY_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20679_ _21357_/CLK _20679_/D repeater199/X vssd1 vssd1 vccd1 vccd1 _20679_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_155_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13220_ _20583_/Q _13215_/X _13219_/X _13217_/X vssd1 vssd1 vccd1 vccd1 _20583_/D
+ sky130_fd_sc_hd__a22o_1
X_10432_ _21296_/Q _10430_/Y _10767_/A _20680_/Q vssd1 vssd1 vccd1 vccd1 _10432_/X
+ sky130_fd_sc_hd__o22a_1
X_13151_ input40/X vssd1 vssd1 vccd1 vccd1 _13151_/X sky130_fd_sc_hd__buf_2
XFILLER_128_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10363_ _10395_/A vssd1 vssd1 vccd1 vccd1 _10381_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__18232__S _18236_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12102_ _20981_/Q _12100_/Y _12321_/A _20382_/Q vssd1 vssd1 vccd1 vccd1 _12102_/X
+ sky130_fd_sc_hd__o22a_1
X_13082_ _20649_/Q _13079_/X _12849_/X _13081_/X vssd1 vssd1 vccd1 vccd1 _20649_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_152_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input57_A HWDATA[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10294_ _10291_/Y _20734_/Q _21353_/Q _10292_/Y _10293_/X vssd1 vssd1 vccd1 vccd1
+ _10307_/A sky130_fd_sc_hd__o221a_1
XFILLER_88_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12033_ _19081_/X _12029_/X _20984_/Q _12030_/X vssd1 vssd1 vccd1 vccd1 _20984_/D
+ sky130_fd_sc_hd__a22o_1
X_16910_ _16910_/A _16910_/B vssd1 vssd1 vccd1 vccd1 _16910_/Y sky130_fd_sc_hd__nor2_1
XFILLER_111_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17890_ _18480_/X _18020_/A _18469_/X _17326_/X vssd1 vssd1 vccd1 vccd1 _17890_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__19375__CLK _19706_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_239_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18470__A0 _17281_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16841_ _16877_/A _16841_/B vssd1 vssd1 vccd1 vccd1 _16841_/Y sky130_fd_sc_hd__nor2_1
XFILLER_77_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19063__S _19910_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19560_ _19706_/CLK _19560_/D vssd1 vssd1 vccd1 vccd1 _19560_/Q sky130_fd_sc_hd__dfxtp_1
X_16772_ _19924_/Q vssd1 vssd1 vccd1 vccd1 _16774_/A sky130_fd_sc_hd__inv_2
X_13984_ _13893_/A _13983_/A _20316_/Q _13983_/Y _13980_/X vssd1 vssd1 vccd1 vccd1
+ _20316_/D sky130_fd_sc_hd__o221a_1
X_18511_ _17281_/X _18061_/Y _18909_/S vssd1 vssd1 vccd1 vccd1 _18511_/X sky130_fd_sc_hd__mux2_1
XFILLER_207_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15723_ _15736_/A vssd1 vssd1 vccd1 vccd1 _15723_/X sky130_fd_sc_hd__buf_1
XFILLER_19_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19491_ _21040_/CLK _19491_/D vssd1 vssd1 vccd1 vccd1 _19491_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12935_ _12960_/A vssd1 vssd1 vccd1 vccd1 _12935_/X sky130_fd_sc_hd__buf_1
XFILLER_18_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18442_ _17079_/Y _12090_/Y _18908_/S vssd1 vssd1 vccd1 vccd1 _18442_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09602__B _19986_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15654_ _16311_/A vssd1 vssd1 vccd1 vccd1 _15722_/A sky130_fd_sc_hd__buf_1
XPHY_4160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12866_ _20746_/Q _12859_/X _12699_/X _12861_/X vssd1 vssd1 vccd1 vccd1 _20746_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14605_ _14605_/A vssd1 vssd1 vccd1 vccd1 _14605_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13598__B1 _13452_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18373_ _18000_/Y _20354_/Q _18787_/S vssd1 vssd1 vccd1 vccd1 _18373_/X sky130_fd_sc_hd__mux2_1
X_11817_ _11817_/A vssd1 vssd1 vccd1 vccd1 _11817_/X sky130_fd_sc_hd__buf_1
XFILLER_14_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15585_ _15788_/A vssd1 vssd1 vccd1 vccd1 _15585_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__16716__A _16718_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18407__S _18906_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12797_ _12803_/A vssd1 vssd1 vccd1 vccd1 _12797_/X sky130_fd_sc_hd__buf_1
XFILLER_187_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17324_ _18065_/A vssd1 vssd1 vccd1 vccd1 _17324_/X sky130_fd_sc_hd__buf_2
XPHY_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14536_ _20136_/Q vssd1 vssd1 vccd1 vccd1 _14536_/X sky130_fd_sc_hd__buf_1
X_11748_ _16502_/A _11748_/B vssd1 vssd1 vccd1 vccd1 _11749_/A sky130_fd_sc_hd__or2_2
XFILLER_175_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_239_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17255_ _17829_/B vssd1 vssd1 vccd1 vccd1 _17533_/B sky130_fd_sc_hd__clkbuf_2
X_14467_ _14467_/A _14524_/C _14467_/C vssd1 vssd1 vccd1 vccd1 _20237_/D sky130_fd_sc_hd__nor3_1
X_11679_ _11689_/A vssd1 vssd1 vccd1 vccd1 _11679_/X sky130_fd_sc_hd__buf_1
X_16206_ _16206_/A vssd1 vssd1 vccd1 vccd1 _16206_/X sky130_fd_sc_hd__buf_1
XANTENNA__13140__A input44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13418_ input44/X vssd1 vssd1 vccd1 vccd1 _13418_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_125_HCLK clkbuf_4_4_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20413_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_127_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17186_ _21342_/Q vssd1 vssd1 vccd1 vccd1 _17186_/Y sky130_fd_sc_hd__inv_2
X_14398_ _21485_/Q _14463_/D _14397_/Y _20210_/Q vssd1 vssd1 vccd1 vccd1 _14398_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12573__A1 _10859_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16137_ _21451_/Q vssd1 vssd1 vccd1 vccd1 _16137_/X sky130_fd_sc_hd__buf_1
XANTENNA__12573__B2 _18242_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18142__S _18896_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13349_ _20519_/Q _13345_/X _13211_/X _13346_/X vssd1 vssd1 vccd1 vccd1 _20519_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20376__RESET_B repeater185/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16068_ _19500_/Q _16064_/X _15762_/X _16066_/X vssd1 vssd1 vccd1 vccd1 _19500_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_115_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15019_ _15019_/A _15019_/B _15019_/C vssd1 vssd1 vccd1 vccd1 _15022_/A sky130_fd_sc_hd__or3_4
XFILLER_130_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18461__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19827_ _19835_/CLK _19827_/D vssd1 vssd1 vccd1 vccd1 _19827_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17282__A _20774_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19758_ _21009_/CLK _19758_/D vssd1 vssd1 vccd1 vccd1 _19758_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_244_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18097__B _18097_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18709_ _17281_/X _17636_/Y _18835_/S vssd1 vssd1 vccd1 vccd1 _18709_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19689_ _19811_/CLK _19689_/D vssd1 vssd1 vccd1 vccd1 _19689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__21164__RESET_B repeater226/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_240_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18516__A1 _20755_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18317__S _18666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20602_ _20693_/CLK _20602_/D repeater195/X vssd1 vssd1 vccd1 vccd1 _20602_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_33_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20533_ _21366_/CLK _20533_/D repeater265/X vssd1 vssd1 vccd1 vccd1 _20533_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_220_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13050__A _13657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20464_ _20495_/CLK _20464_/D repeater273/X vssd1 vssd1 vccd1 vccd1 _20464_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_229_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_3_4_0_HCLK clkbuf_3_5_0_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_9_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_20395_ _20951_/CLK _20395_/D repeater272/X vssd1 vssd1 vccd1 vccd1 _20395_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_106_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20046__RESET_B repeater281/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13513__B1 _13442_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21016_ _21431_/CLK _21016_/D repeater238/X vssd1 vssd1 vccd1 vccd1 _21016_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__18452__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15705__A input38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13816__A1 _20611_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09709_ _21461_/Q _21460_/Q _21462_/Q vssd1 vssd1 vccd1 vccd1 _09770_/B sky130_fd_sc_hd__and3_1
X_10981_ _16594_/A _11875_/B vssd1 vssd1 vccd1 vccd1 _11883_/A sky130_fd_sc_hd__nand2_1
XFILLER_43_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12720_ _12898_/A vssd1 vssd1 vccd1 vccd1 _17177_/A sky130_fd_sc_hd__buf_4
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19982__RESET_B repeater276/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12651_ input62/X vssd1 vssd1 vccd1 vccd1 _12651_/X sky130_fd_sc_hd__clkbuf_4
XPHY_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18227__S _18236_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11602_ _18987_/X _11598_/X _21119_/Q _11600_/X vssd1 vssd1 vccd1 vccd1 _21119_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19911__RESET_B repeater220/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15370_ _19823_/Q _15366_/X _15352_/X _15367_/X vssd1 vssd1 vccd1 vccd1 _19823_/D
+ sky130_fd_sc_hd__a22o_1
X_12582_ _12582_/A vssd1 vssd1 vccd1 vccd1 _12601_/A sky130_fd_sc_hd__clkbuf_2
XPHY_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_148_HCLK clkbuf_opt_1_HCLK/A vssd1 vssd1 vccd1 vccd1 _21235_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14321_ _20128_/Q vssd1 vssd1 vccd1 vccd1 _16034_/A sky130_fd_sc_hd__buf_1
XPHY_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11533_ _21140_/Q _11527_/X _10892_/X _11529_/X vssd1 vssd1 vccd1 vccd1 _21140_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10584__A _20750_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17040_ _21413_/Q vssd1 vssd1 vccd1 vccd1 _17040_/Y sky130_fd_sc_hd__inv_2
XPHY_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14252_ _20254_/Q _14246_/A _20253_/Q _14249_/X vssd1 vssd1 vccd1 vccd1 _20254_/D
+ sky130_fd_sc_hd__a22o_1
X_11464_ _19091_/X _11461_/X _21167_/Q _11463_/X vssd1 vssd1 vccd1 vccd1 _21167_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_144_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19058__S _19058_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13203_ _20591_/Q _13200_/X _12999_/X _13201_/X vssd1 vssd1 vccd1 vccd1 _20591_/D
+ sky130_fd_sc_hd__a22o_1
X_10415_ _10415_/A vssd1 vssd1 vccd1 vccd1 _10415_/Y sky130_fd_sc_hd__inv_2
X_11395_ _19870_/Q _16507_/A vssd1 vssd1 vccd1 vccd1 _11395_/Y sky130_fd_sc_hd__nor2_2
X_14183_ _14191_/A vssd1 vssd1 vccd1 vccd1 _14183_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_164_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13134_ _20618_/Q _13132_/X _12925_/X _13133_/X vssd1 vssd1 vccd1 vccd1 _20618_/D
+ sky130_fd_sc_hd__a22o_1
X_10346_ _10346_/A vssd1 vssd1 vccd1 vccd1 _10346_/X sky130_fd_sc_hd__buf_1
X_18991_ _21262_/Q _21114_/Q _18992_/S vssd1 vssd1 vccd1 vccd1 _18991_/X sky130_fd_sc_hd__mux2_1
XANTENNA__18897__S _18897_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13504__B1 _13313_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17942_ _17942_/A _17943_/B vssd1 vssd1 vccd1 vccd1 _17942_/Y sky130_fd_sc_hd__nor2_1
X_13065_ _20658_/Q _13060_/X _13003_/X _13061_/X vssd1 vssd1 vccd1 vccd1 _20658_/D
+ sky130_fd_sc_hd__a22o_1
X_10277_ _10277_/A _10277_/B vssd1 vssd1 vccd1 vccd1 _10388_/A sky130_fd_sc_hd__or2_1
XFILLER_151_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_repeater209_A repeater211/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12016_ _19070_/X _12010_/X _20995_/Q _12012_/X vssd1 vssd1 vccd1 vccd1 _20995_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_39_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater208 repeater209/X vssd1 vssd1 vccd1 vccd1 repeater208/X sky130_fd_sc_hd__buf_6
X_17873_ _18570_/X _17861_/X _18552_/X _17862_/X _17872_/X vssd1 vssd1 vccd1 vccd1
+ _17873_/X sky130_fd_sc_hd__o221a_2
Xrepeater219 repeater220/X vssd1 vssd1 vccd1 vccd1 repeater219/X sky130_fd_sc_hd__buf_8
XANTENNA__20868__CLK _21452_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19612_ _21040_/CLK _19612_/D vssd1 vssd1 vccd1 vccd1 _19612_/Q sky130_fd_sc_hd__dfxtp_1
X_16824_ _16822_/A _16822_/C _19936_/Q vssd1 vssd1 vccd1 vccd1 _16824_/X sky130_fd_sc_hd__o21a_1
XFILLER_38_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19543_ _21462_/CLK _19543_/D vssd1 vssd1 vccd1 vccd1 _19543_/Q sky130_fd_sc_hd__dfxtp_1
X_16755_ _19920_/Q vssd1 vssd1 vccd1 vccd1 _16755_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13967_ _13990_/A vssd1 vssd1 vccd1 vccd1 _14037_/C sky130_fd_sc_hd__clkbuf_2
X_15706_ _16016_/A vssd1 vssd1 vccd1 vccd1 _15706_/X sky130_fd_sc_hd__buf_1
XFILLER_207_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12918_ input52/X vssd1 vssd1 vccd1 vccd1 _12918_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_74_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19474_ _21222_/CLK _19474_/D vssd1 vssd1 vccd1 vccd1 _19474_/Q sky130_fd_sc_hd__dfxtp_1
X_16686_ _16686_/A vssd1 vssd1 vccd1 vccd1 _16686_/Y sky130_fd_sc_hd__inv_2
X_13898_ _13898_/A vssd1 vssd1 vccd1 vccd1 _13898_/Y sky130_fd_sc_hd__inv_2
XFILLER_222_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18425_ _18424_/X _14895_/Y _18907_/S vssd1 vssd1 vccd1 vccd1 _18425_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15637_ _19702_/Q _15632_/X _15592_/X _15633_/X vssd1 vssd1 vccd1 vccd1 _19702_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_222_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12849_ _12849_/A vssd1 vssd1 vccd1 vccd1 _12849_/X sky130_fd_sc_hd__buf_2
XANTENNA__18137__S _18787_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12974__A _17178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15350__A _15588_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18356_ _18355_/X _13958_/Y _18849_/S vssd1 vssd1 vccd1 vccd1 _18356_/X sky130_fd_sc_hd__mux2_1
X_15568_ _15568_/A vssd1 vssd1 vccd1 vccd1 _15568_/X sky130_fd_sc_hd__buf_1
XFILLER_14_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17307_ _17305_/Y _17142_/A _17306_/Y _17154_/X vssd1 vssd1 vccd1 vccd1 _17307_/X
+ sky130_fd_sc_hd__o22a_1
X_14519_ _14351_/B _14521_/A _14351_/A vssd1 vssd1 vccd1 vccd1 _14520_/B sky130_fd_sc_hd__o21a_1
X_18287_ _18286_/X _10776_/A _18617_/S vssd1 vssd1 vccd1 vccd1 _18287_/X sky130_fd_sc_hd__mux2_1
X_15499_ _15499_/A vssd1 vssd1 vccd1 vccd1 _15499_/X sky130_fd_sc_hd__buf_1
XFILLER_175_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20557__RESET_B repeater267/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17238_ _19695_/Q vssd1 vssd1 vccd1 vccd1 _17238_/Y sky130_fd_sc_hd__inv_2
XFILLER_143_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17169_ _17169_/A _17169_/B _17169_/C _17169_/D vssd1 vssd1 vccd1 vccd1 _17560_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_89_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20180_ _21483_/CLK _20180_/D repeater200/X vssd1 vssd1 vccd1 vccd1 _20180_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_131_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09991_ _21420_/Q vssd1 vssd1 vccd1 vccd1 _09991_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15496__B1 _15454_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19690__CLK _19813_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18600__S _18902_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_29_HCLK clkbuf_opt_4_HCLK/A vssd1 vssd1 vccd1 vccd1 _21429_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_85_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11521__A2 _11497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21345__RESET_B repeater255/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_244_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12884__A _13714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_240_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20516_ _20944_/CLK _20516_/D repeater277/X vssd1 vssd1 vccd1 vccd1 _20516_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_181_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20227__RESET_B repeater200/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20447_ _20480_/CLK _20447_/D repeater183/X vssd1 vssd1 vccd1 vccd1 _20447_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_146_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10200_ _10221_/A _10220_/A _10200_/C vssd1 vssd1 vccd1 vccd1 _10218_/A sky130_fd_sc_hd__or3_1
XFILLER_180_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11180_ _21218_/Q vssd1 vssd1 vccd1 vccd1 _11180_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_109_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20378_ _20957_/CLK _20378_/D repeater185/X vssd1 vssd1 vccd1 vccd1 _20378_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_134_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10131_ _10154_/A _20790_/Q _10158_/A _20794_/Q _10130_/X vssd1 vssd1 vccd1 vccd1
+ _10136_/C sky130_fd_sc_hd__o221a_1
XANTENNA__18510__S _18898_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18425__A0 _18424_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10062_ _10158_/A _10157_/A _10150_/A _10149_/A vssd1 vssd1 vccd1 vccd1 _10068_/C
+ sky130_fd_sc_hd__or4_4
XFILLER_88_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11512__A2 _11497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14870_ _14961_/D _14870_/B vssd1 vssd1 vccd1 vccd1 _14987_/A sky130_fd_sc_hd__or2_1
XFILLER_236_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13821_ _20203_/Q vssd1 vssd1 vccd1 vccd1 _14592_/A sky130_fd_sc_hd__inv_2
XANTENNA__21015__RESET_B repeater238/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16540_ _21195_/Q _21194_/Q _21196_/Q vssd1 vssd1 vccd1 vccd1 _16561_/A sky130_fd_sc_hd__or3_4
XANTENNA__17650__A _21141_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13752_ _20623_/Q vssd1 vssd1 vccd1 vccd1 _18032_/A sky130_fd_sc_hd__inv_2
X_10964_ _11804_/C vssd1 vssd1 vccd1 vccd1 _10964_/X sky130_fd_sc_hd__buf_1
XFILLER_232_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12703_ _20818_/Q _12701_/X _12544_/X _12702_/X vssd1 vssd1 vccd1 vccd1 _20818_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_44_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_105_HCLK_A clkbuf_4_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17400__A1 _18810_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16471_ _19297_/Q _16466_/X _16283_/X _16468_/X vssd1 vssd1 vccd1 vccd1 _19297_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_204_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13683_ _20349_/Q _13679_/X _13487_/X _13680_/X vssd1 vssd1 vccd1 vccd1 _20349_/D
+ sky130_fd_sc_hd__a22o_1
X_10895_ _21253_/Q _10888_/X _10894_/X _10890_/X vssd1 vssd1 vccd1 vccd1 _21253_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_168_HCLK_A clkbuf_opt_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18210_ _18209_/X _12260_/Y _18910_/S vssd1 vssd1 vccd1 vccd1 _18210_/X sky130_fd_sc_hd__mux2_1
X_15422_ _19802_/Q _15415_/X _15421_/X _15417_/X vssd1 vssd1 vccd1 vccd1 _19802_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12634_ input30/X _12631_/X _20850_/Q _12632_/X vssd1 vssd1 vccd1 vccd1 _20850_/D
+ sky130_fd_sc_hd__o22a_1
X_19190_ _19305_/Q _19827_/Q _19835_/Q _19419_/Q _19280_/S0 _20122_/Q vssd1 vssd1
+ vccd1 vccd1 _19190_/X sky130_fd_sc_hd__mux4_2
XPHY_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18141_ _18140_/X _14573_/A _18748_/S vssd1 vssd1 vccd1 vccd1 _18141_/X sky130_fd_sc_hd__mux2_2
X_15353_ _19831_/Q _15345_/X _15352_/X _15347_/X vssd1 vssd1 vccd1 vccd1 _19831_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12565_ _12580_/A vssd1 vssd1 vccd1 vccd1 _12574_/A sky130_fd_sc_hd__buf_1
XPHY_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_repeater159_A _18850_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14304_ _14304_/A _17320_/A vssd1 vssd1 vccd1 vccd1 _14730_/B sky130_fd_sc_hd__or2_1
XFILLER_200_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18072_ _18670_/X _17205_/X _18622_/X _18045_/X vssd1 vssd1 vccd1 vccd1 _18072_/X
+ sky130_fd_sc_hd__o22a_2
XANTENNA__15175__C1 _15201_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11516_ _16340_/A vssd1 vssd1 vccd1 vccd1 _11516_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20540__CLK _20592_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15284_ _15284_/A _15284_/B _15284_/C _15284_/D vssd1 vssd1 vccd1 vccd1 _15285_/D
+ sky130_fd_sc_hd__and4_1
XPHY_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12496_ _12496_/A _12496_/B _12496_/C vssd1 vssd1 vccd1 vccd1 _20919_/D sky130_fd_sc_hd__nor3_2
XANTENNA__17809__B _17812_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17023_ _17023_/A _17023_/B vssd1 vssd1 vccd1 vccd1 _20009_/D sky130_fd_sc_hd__nor2_1
X_14235_ _19895_/Q _14235_/B vssd1 vssd1 vccd1 vccd1 _14236_/B sky130_fd_sc_hd__or2_1
X_11447_ _21159_/Q _11447_/B vssd1 vssd1 vccd1 vccd1 _11448_/B sky130_fd_sc_hd__or2_1
XFILLER_109_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11378_ _21170_/Q vssd1 vssd1 vccd1 vccd1 _11386_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA_output88_A _17966_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14166_ _14163_/Y _20265_/Q _14164_/Y _20275_/Q _14165_/X vssd1 vssd1 vccd1 vccd1
+ _14170_/C sky130_fd_sc_hd__o221a_1
XFILLER_125_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13117_ _20629_/Q _13112_/X _12989_/X _13115_/X vssd1 vssd1 vccd1 vccd1 _20629_/D
+ sky130_fd_sc_hd__a22o_1
X_10329_ _20706_/Q vssd1 vssd1 vccd1 vccd1 _10329_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14097_ _14097_/A _14097_/B vssd1 vssd1 vccd1 vccd1 _14179_/A sky130_fd_sc_hd__or2_1
XANTENNA__18420__S _18904_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18974_ _13182_/X _13177_/Y _18975_/S vssd1 vssd1 vccd1 vccd1 _18974_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17544__B _17807_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17925_ _17925_/A vssd1 vssd1 vccd1 vccd1 _17925_/X sky130_fd_sc_hd__buf_1
XFILLER_67_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13048_ _13048_/A _17209_/A vssd1 vssd1 vccd1 vccd1 _13262_/B sky130_fd_sc_hd__or2_2
X_17856_ _17856_/A vssd1 vssd1 vccd1 vccd1 _17856_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16807_ _16820_/A _16807_/B vssd1 vssd1 vccd1 vccd1 _16807_/Y sky130_fd_sc_hd__nor2_1
XFILLER_226_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17787_ _17783_/Y _11678_/A _16634_/A _17553_/X _17786_/X vssd1 vssd1 vccd1 vccd1
+ _17787_/X sky130_fd_sc_hd__o221a_1
XFILLER_53_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14999_ _15019_/A _15019_/B _14999_/C vssd1 vssd1 vccd1 vccd1 _15017_/A sky130_fd_sc_hd__or3_1
X_16738_ _21144_/Q _16738_/B vssd1 vssd1 vccd1 vccd1 _16738_/X sky130_fd_sc_hd__or2_1
X_19526_ _19784_/CLK _19526_/D vssd1 vssd1 vccd1 vccd1 _19526_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_241_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19457_ _20137_/CLK _19457_/D vssd1 vssd1 vccd1 vccd1 _19457_/Q sky130_fd_sc_hd__dfxtp_1
X_16669_ _21157_/Q _11445_/B _11446_/B vssd1 vssd1 vccd1 vccd1 _16669_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__20738__RESET_B repeater205/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18408_ _18407_/X _14919_/Y _18907_/S vssd1 vssd1 vccd1 vccd1 _18408_/X sky130_fd_sc_hd__mux2_2
X_19388_ _20432_/CLK _19388_/D vssd1 vssd1 vccd1 vccd1 _19388_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_27_HCLK_A clkbuf_opt_4_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18339_ _17984_/Y _16970_/Y _18680_/S vssd1 vssd1 vccd1 vccd1 _18339_/X sky130_fd_sc_hd__mux2_2
XANTENNA__12209__A _20501_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20391__RESET_B repeater278/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21350_ _21407_/CLK _21350_/D repeater252/X vssd1 vssd1 vccd1 vccd1 _21350_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_147_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20320__RESET_B repeater262/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20301_ _20693_/CLK _20301_/D repeater197/X vssd1 vssd1 vccd1 vccd1 _20301_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_162_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21281_ _21342_/CLK _21281_/D repeater211/X vssd1 vssd1 vccd1 vccd1 _21281_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18104__C1 _18103_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20232_ _21484_/CLK _20232_/D repeater203/X vssd1 vssd1 vccd1 vccd1 _20232_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_2_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17157__D _17157_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20163_ _21121_/CLK _20163_/D repeater237/X vssd1 vssd1 vccd1 vccd1 _20163_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18330__S _18669_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09974_ _21418_/Q _09968_/X _09676_/X _09970_/X vssd1 vssd1 vccd1 vccd1 _21418_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_39_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14141__B1 _20547_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20094_ _20101_/CLK _20094_/D repeater273/X vssd1 vssd1 vccd1 vccd1 _20094_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12879__A _13710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_218_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19887__SET_B repeater217/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20996_ _21185_/CLK _20996_/D repeater222/X vssd1 vssd1 vccd1 vccd1 _20996_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_72_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10680_ _10694_/A vssd1 vssd1 vccd1 vccd1 _10680_/X sky130_fd_sc_hd__buf_1
XANTENNA__12207__B1 _20982_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_213_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20408__RESET_B repeater184/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19230__S1 _20131_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18505__S _18884_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12350_ _12350_/A vssd1 vssd1 vccd1 vccd1 _12350_/X sky130_fd_sc_hd__buf_2
XFILLER_138_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20061__RESET_B repeater281/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_217_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11301_ _11301_/A _11301_/B vssd1 vssd1 vccd1 vccd1 _12500_/B sky130_fd_sc_hd__nand2_1
XFILLER_181_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12281_ _20929_/Q _20509_/Q _12398_/C _12280_/Y vssd1 vssd1 vccd1 vccd1 _12281_/X
+ sky130_fd_sc_hd__o22a_1
X_21479_ _21481_/CLK _21479_/D repeater206/X vssd1 vssd1 vccd1 vccd1 _21479_/Q sky130_fd_sc_hd__dfrtp_1
X_11232_ _19911_/Q vssd1 vssd1 vccd1 vccd1 _11233_/C sky130_fd_sc_hd__inv_2
X_14020_ _14020_/A vssd1 vssd1 vccd1 vccd1 _14020_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11194__B1 _10892_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11163_ _15638_/C vssd1 vssd1 vccd1 vccd1 _16593_/B sky130_fd_sc_hd__inv_2
XANTENNA__20004__SET_B repeater225/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18240__S _18242_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10114_ _21382_/Q _10081_/Y _10041_/A _20776_/Q _10113_/X vssd1 vssd1 vccd1 vccd1
+ _10114_/X sky130_fd_sc_hd__a221o_1
XFILLER_96_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15971_ _15979_/A vssd1 vssd1 vccd1 vccd1 _15971_/X sky130_fd_sc_hd__buf_1
XFILLER_49_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11094_ _11090_/B _11079_/X _11093_/X _11082_/X _11093_/A vssd1 vssd1 vccd1 vccd1
+ _11095_/A sky130_fd_sc_hd__o32a_1
XFILLER_248_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18949__A1 _21087_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14683__A1 _10985_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17710_ _20403_/Q vssd1 vssd1 vccd1 vccd1 _17710_/Y sky130_fd_sc_hd__inv_2
X_14922_ _20588_/Q vssd1 vssd1 vccd1 vccd1 _14922_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10045_ _21376_/Q vssd1 vssd1 vccd1 vccd1 _10199_/A sky130_fd_sc_hd__inv_2
X_18690_ _18689_/X _14424_/Y _18897_/S vssd1 vssd1 vccd1 vccd1 _18690_/X sky130_fd_sc_hd__mux2_1
XFILLER_248_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17641_ _21085_/Q vssd1 vssd1 vccd1 vccd1 _17641_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14853_ _14853_/A _14853_/B _15019_/C vssd1 vssd1 vccd1 vccd1 _14999_/C sky130_fd_sc_hd__or3_1
XFILLER_35_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output126_A _17089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19071__S _19908_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13804_ _20625_/Q _14591_/A _13800_/Y _20176_/Q _13803_/X vssd1 vssd1 vccd1 vccd1
+ _13811_/C sky130_fd_sc_hd__o221a_1
XANTENNA__12446__B1 _12445_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17572_ _18748_/X _17572_/B vssd1 vssd1 vccd1 vccd1 _17572_/Y sky130_fd_sc_hd__nand2_2
X_14784_ _14784_/A vssd1 vssd1 vccd1 vccd1 _14787_/A sky130_fd_sc_hd__inv_2
XFILLER_223_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11996_ _20990_/Q _11996_/B vssd1 vssd1 vccd1 vccd1 _11997_/B sky130_fd_sc_hd__or2_1
XFILLER_28_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19311_ _20142_/CLK _19311_/D vssd1 vssd1 vccd1 vccd1 _19311_/Q sky130_fd_sc_hd__dfxtp_1
X_16523_ _16523_/A vssd1 vssd1 vccd1 vccd1 _20002_/D sky130_fd_sc_hd__inv_2
X_13735_ _20631_/Q vssd1 vssd1 vccd1 vccd1 _13735_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10947_ _21207_/Q vssd1 vssd1 vccd1 vccd1 _10947_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19242_ _17407_/Y _17408_/Y _17409_/Y _17410_/Y _19275_/S0 _21004_/Q vssd1 vssd1
+ vccd1 vccd1 _19242_/X sky130_fd_sc_hd__mux4_2
X_16454_ _16460_/A vssd1 vssd1 vccd1 vccd1 _16454_/X sky130_fd_sc_hd__buf_1
XFILLER_31_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13666_ _20360_/Q _13659_/X _13547_/X _13662_/X vssd1 vssd1 vccd1 vccd1 _20360_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19126__A1 _14275_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10878_ _10880_/A vssd1 vssd1 vccd1 vccd1 _10888_/A sky130_fd_sc_hd__buf_1
XANTENNA__20149__RESET_B repeater250/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15405_ _15405_/A vssd1 vssd1 vccd1 vccd1 _15405_/X sky130_fd_sc_hd__buf_1
XPHY_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12617_ input10/X _12613_/X _20861_/Q _12614_/X vssd1 vssd1 vccd1 vccd1 _20861_/D
+ sky130_fd_sc_hd__o22a_1
X_19173_ _19544_/Q _19536_/Q _19528_/Q _19512_/Q _19280_/S0 _20122_/Q vssd1 vssd1
+ vccd1 vccd1 _19173_/X sky130_fd_sc_hd__mux4_1
XPHY_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16385_ _16385_/A vssd1 vssd1 vccd1 vccd1 _16385_/X sky130_fd_sc_hd__buf_1
XPHY_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19221__S1 _20133_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18415__S _18680_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13597_ _20399_/Q _13594_/X _13449_/X _13595_/X vssd1 vssd1 vccd1 vccd1 _20399_/D
+ sky130_fd_sc_hd__a22o_1
X_18124_ vssd1 vssd1 vccd1 vccd1 _18124_/HI _18124_/LO sky130_fd_sc_hd__conb_1
XFILLER_157_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15336_ _15448_/A _15967_/B _15999_/C vssd1 vssd1 vccd1 vccd1 _15345_/A sky130_fd_sc_hd__or3_4
X_12548_ _12548_/A vssd1 vssd1 vccd1 vccd1 _12548_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_118_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17539__B _17542_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18055_ _18133_/X _18021_/X _18338_/X _18045_/X vssd1 vssd1 vccd1 vccd1 _18055_/X
+ sky130_fd_sc_hd__o22a_2
X_15267_ _15266_/Y _20056_/Q _20473_/Q _15093_/X vssd1 vssd1 vccd1 vccd1 _15267_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__14244__A _14246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12479_ _12479_/A vssd1 vssd1 vccd1 vccd1 _12479_/Y sky130_fd_sc_hd__inv_2
XFILLER_144_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17006_ _17013_/A _17006_/B vssd1 vssd1 vccd1 vccd1 _17006_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__18637__A0 _18848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14218_ _14078_/A _14078_/B _14216_/Y _14207_/X vssd1 vssd1 vccd1 vccd1 _20267_/D
+ sky130_fd_sc_hd__a211oi_2
X_15198_ _15198_/A vssd1 vssd1 vccd1 vccd1 _15201_/A sky130_fd_sc_hd__inv_2
XANTENNA__18101__A2 _17205_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14149_ _14147_/Y _20284_/Q _14148_/Y _20270_/Q vssd1 vssd1 vccd1 vccd1 _14149_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__18150__S _18787_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18957_ _16644_/X _21079_/Q _18962_/S vssd1 vssd1 vccd1 vccd1 _18957_/X sky130_fd_sc_hd__mux2_1
XFILLER_112_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17908_ _17908_/A vssd1 vssd1 vccd1 vccd1 _17908_/X sky130_fd_sc_hd__buf_1
XFILLER_239_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09690_ _15329_/A vssd1 vssd1 vccd1 vccd1 _09690_/X sky130_fd_sc_hd__buf_1
X_18888_ _18887_/X _10421_/Y _18910_/S vssd1 vssd1 vccd1 vccd1 _18888_/X sky130_fd_sc_hd__mux2_1
XFILLER_66_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17839_ _17839_/A vssd1 vssd1 vccd1 vccd1 _17839_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_26_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14426__B2 _21486_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17290__A _17290_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_212_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20850_ _20857_/CLK _20850_/D repeater243/X vssd1 vssd1 vccd1 vccd1 _20850_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12988__A1 _20697_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19509_ _20327_/CLK _19509_/D vssd1 vssd1 vccd1 vccd1 _19509_/Q sky130_fd_sc_hd__dfxtp_1
X_20781_ _21406_/CLK _20781_/D repeater213/X vssd1 vssd1 vccd1 vccd1 _20781_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17915__A2 _18024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11660__A1 _11486_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19117__A1 _11123_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_151_HCLK_A clkbuf_4_4_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18325__S _18784_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19212__S1 _21004_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21402_ _21405_/CLK _21402_/D repeater255/X vssd1 vssd1 vccd1 vccd1 _21402_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_157_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21333_ _21476_/CLK _21333_/D repeater204/X vssd1 vssd1 vccd1 vccd1 _21333_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__18628__A0 _17079_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21264_ _21417_/CLK _21264_/D repeater234/X vssd1 vssd1 vccd1 vccd1 _21264_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_116_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20215_ _20220_/CLK _20215_/D repeater202/X vssd1 vssd1 vccd1 vccd1 _20215_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_173_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17465__A _21144_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21195_ _21196_/CLK _21195_/D repeater220/X vssd1 vssd1 vccd1 vccd1 _21195_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__21360__RESET_B repeater254/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20146_ _21239_/CLK _20146_/D repeater250/X vssd1 vssd1 vccd1 vccd1 _20146_/Q sky130_fd_sc_hd__dfrtp_1
X_09957_ _09957_/A vssd1 vssd1 vccd1 vccd1 _09957_/X sky130_fd_sc_hd__buf_1
XANTENNA__19279__S1 _20122_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18995__S _19026_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12676__B1 _09621_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20077_ _20107_/CLK _20077_/D repeater259/X vssd1 vssd1 vccd1 vccd1 _20077_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_100_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09888_ _20012_/Q _09887_/B _09887_/Y vssd1 vssd1 vccd1 vccd1 _17026_/A sky130_fd_sc_hd__o21ai_1
XFILLER_245_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_245_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11850_ _11850_/A vssd1 vssd1 vccd1 vccd1 _11851_/B sky130_fd_sc_hd__inv_2
XFILLER_122_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10801_ _10801_/A vssd1 vssd1 vccd1 vccd1 _10801_/Y sky130_fd_sc_hd__inv_2
XPHY_4567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11781_ _11781_/A vssd1 vssd1 vccd1 vccd1 _21043_/D sky130_fd_sc_hd__inv_2
XPHY_3833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20979_ _20981_/CLK _20979_/D repeater187/X vssd1 vssd1 vccd1 vccd1 _20979_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_3855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17906__A2 _17200_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13520_ _11973_/A _18975_/S _18973_/X vssd1 vssd1 vccd1 vccd1 _13520_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_241_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10732_ _19943_/Q _19942_/Q vssd1 vssd1 vccd1 vccd1 _10748_/C sky130_fd_sc_hd__or2_1
XPHY_3877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13451_ _15523_/A vssd1 vssd1 vccd1 vccd1 _15429_/A sky130_fd_sc_hd__clkbuf_2
X_10663_ _10663_/A _10663_/B vssd1 vssd1 vccd1 vccd1 _10675_/A sky130_fd_sc_hd__or2_2
XANTENNA__18235__S _18236_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19203__S1 _21004_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12402_ _12425_/A _12424_/A _12426_/A _12423_/A vssd1 vssd1 vccd1 vccd1 _12403_/D
+ sky130_fd_sc_hd__or4_4
XANTENNA_clkbuf_leaf_10_HCLK_A clkbuf_opt_2_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16170_ _19452_/Q _16166_/X _16135_/X _16168_/X vssd1 vssd1 vccd1 vccd1 _19452_/D
+ sky130_fd_sc_hd__a22o_1
X_10594_ _10707_/A _20747_/Q _21319_/Q _10593_/Y vssd1 vssd1 vccd1 vccd1 _10594_/X
+ sky130_fd_sc_hd__o22a_1
X_13382_ _20498_/Q _13377_/X _13173_/X _13378_/X vssd1 vssd1 vccd1 vccd1 _20498_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_139_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_73_HCLK_A clkbuf_opt_7_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15121_ _20433_/Q _15059_/A _15097_/Y _15098_/X _15120_/X vssd1 vssd1 vccd1 vccd1
+ _15121_/X sky130_fd_sc_hd__o221a_1
X_12333_ _12333_/A _12333_/B vssd1 vssd1 vccd1 vccd1 _12334_/A sky130_fd_sc_hd__or2_1
XANTENNA__21448__RESET_B repeater248/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15052_ _20050_/Q vssd1 vssd1 vccd1 vccd1 _15065_/A sky130_fd_sc_hd__inv_2
XFILLER_142_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12264_ _20508_/Q vssd1 vssd1 vccd1 vccd1 _12264_/Y sky130_fd_sc_hd__inv_2
XFILLER_147_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14003_ _20306_/Q _14002_/Y _13883_/B _13988_/X vssd1 vssd1 vccd1 vccd1 _20306_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__19066__S _19910_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17375__A _21082_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11215_ _21208_/Q _11213_/X _09655_/X _11214_/X vssd1 vssd1 vccd1 vccd1 _21208_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11200__B _17838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19860_ _21164_/CLK _19860_/D repeater226/X vssd1 vssd1 vccd1 vccd1 _19860_/Q sky130_fd_sc_hd__dfrtp_1
X_12195_ _20334_/Q vssd1 vssd1 vccd1 vccd1 _12195_/Y sky130_fd_sc_hd__inv_2
XFILLER_122_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18811_ _18845_/A0 _13763_/Y _18896_/S vssd1 vssd1 vccd1 vccd1 _18811_/X sky130_fd_sc_hd__mux2_1
XANTENNA__19751__CLK _19765_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput83 _17892_/Y vssd1 vssd1 vccd1 vccd1 HRDATA[13] sky130_fd_sc_hd__clkbuf_2
XANTENNA__17842__B2 _18019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11146_ _21220_/Q vssd1 vssd1 vccd1 vccd1 _15638_/A sky130_fd_sc_hd__inv_2
Xoutput94 _18027_/Y vssd1 vssd1 vccd1 vccd1 HRDATA[23] sky130_fd_sc_hd__clkbuf_2
X_19791_ _19820_/CLK _19791_/D vssd1 vssd1 vccd1 vccd1 _19791_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__21030__RESET_B repeater242/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18742_ _17546_/Y _16766_/A _18880_/S vssd1 vssd1 vccd1 vccd1 _18742_/X sky130_fd_sc_hd__mux2_2
X_15954_ _15961_/A vssd1 vssd1 vccd1 vccd1 _15954_/X sky130_fd_sc_hd__buf_1
X_11077_ _11072_/B _11051_/X _11075_/Y _11076_/X _11061_/A vssd1 vssd1 vccd1 vccd1
+ _11078_/A sky130_fd_sc_hd__o32a_1
XANTENNA__12667__B1 _12666_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14905_ _14902_/Y _20089_/Q _20578_/Q _14960_/C _14904_/X vssd1 vssd1 vccd1 vccd1
+ _14918_/A sky130_fd_sc_hd__o221a_1
X_10028_ _09931_/X _21408_/Q _10028_/S vssd1 vssd1 vccd1 vccd1 _21408_/D sky130_fd_sc_hd__mux2_1
X_18673_ _17775_/Y _19201_/X _18930_/S vssd1 vssd1 vccd1 vccd1 _18673_/X sky130_fd_sc_hd__mux2_2
XANTENNA__14408__A1 _21471_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15885_ _15885_/A _16485_/A vssd1 vssd1 vccd1 vccd1 _15896_/A sky130_fd_sc_hd__or2_2
XFILLER_63_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17624_ _19443_/Q vssd1 vssd1 vccd1 vccd1 _17624_/Y sky130_fd_sc_hd__inv_2
X_14836_ _20097_/Q vssd1 vssd1 vccd1 vccd1 _14960_/A sky130_fd_sc_hd__inv_2
XFILLER_17_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09621__A input52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19870__SET_B repeater225/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17555_ _21076_/Q vssd1 vssd1 vccd1 vccd1 _17555_/Y sky130_fd_sc_hd__inv_2
X_14767_ _20132_/Q _14758_/B _15816_/A _15799_/A _14753_/B vssd1 vssd1 vccd1 vccd1
+ _14767_/X sky130_fd_sc_hd__a32o_1
XFILLER_44_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11979_ _21001_/Q _11978_/Y _11975_/X vssd1 vssd1 vccd1 vccd1 _21001_/D sky130_fd_sc_hd__o21a_1
XFILLER_189_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16506_ _16503_/A _16494_/X _16505_/X vssd1 vssd1 vccd1 vccd1 _20001_/D sky130_fd_sc_hd__o21ai_1
X_13718_ _13727_/A vssd1 vssd1 vccd1 vccd1 _13725_/S sky130_fd_sc_hd__clkbuf_2
X_17486_ _19698_/Q vssd1 vssd1 vccd1 vccd1 _17486_/Y sky130_fd_sc_hd__inv_2
X_14698_ _18245_/X _14696_/X _20162_/Q _14688_/X vssd1 vssd1 vccd1 vccd1 _20162_/D
+ sky130_fd_sc_hd__o22a_1
X_16437_ _19316_/Q _16434_/X _11486_/X _16436_/X vssd1 vssd1 vccd1 vccd1 _19316_/D
+ sky130_fd_sc_hd__a22o_1
X_19225_ _17600_/Y _17601_/Y _17602_/Y _17603_/Y _19275_/S0 _21004_/Q vssd1 vssd1
+ vccd1 vccd1 _19225_/X sky130_fd_sc_hd__mux4_1
XFILLER_177_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13649_ _20369_/Q _13645_/X _13511_/X _13646_/X vssd1 vssd1 vccd1 vccd1 _20369_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_20_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18145__S _18884_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19156_ _19152_/X _19153_/X _19154_/X _19155_/X _21018_/Q _21019_/Q vssd1 vssd1 vccd1
+ vccd1 _19156_/X sky130_fd_sc_hd__mux4_2
X_16368_ _19354_/Q _16363_/X _16202_/X _16365_/X vssd1 vssd1 vccd1 vccd1 _19354_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_191_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18107_ _21223_/Q _17346_/Y _17252_/Y _20999_/Q vssd1 vssd1 vccd1 vccd1 _18107_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_191_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15319_ _09840_/X _15320_/B _09851_/X _15318_/A vssd1 vssd1 vccd1 vccd1 _20034_/D
+ sky130_fd_sc_hd__a22o_1
X_19087_ _21046_/Q _21059_/Q _19872_/Q vssd1 vssd1 vccd1 vccd1 _19087_/X sky130_fd_sc_hd__mux2_1
XFILLER_184_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16299_ _16305_/A vssd1 vssd1 vccd1 vccd1 _16306_/A sky130_fd_sc_hd__inv_2
XANTENNA__13147__A1 _20612_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18038_ _18351_/X _17947_/X _18252_/X _17948_/X vssd1 vssd1 vccd1 vccd1 _18042_/A
+ sky130_fd_sc_hd__o22ai_2
XFILLER_133_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21118__RESET_B repeater233/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20000_ _21167_/CLK _20000_/D repeater225/X vssd1 vssd1 vccd1 vccd1 _20000_/Q sky130_fd_sc_hd__dfrtp_1
X_09811_ _21453_/Q vssd1 vssd1 vccd1 vccd1 _15865_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_87_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19989_ _21055_/CLK _19989_/D repeater218/X vssd1 vssd1 vccd1 vccd1 _19989_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_141_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09742_ _09732_/X _09742_/B _09742_/C _09742_/D vssd1 vssd1 vccd1 vccd1 _09769_/C
+ sky130_fd_sc_hd__and4b_1
XANTENNA__19130__S0 _19285_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09673_ _15329_/A vssd1 vssd1 vccd1 vccd1 _09673_/X sky130_fd_sc_hd__buf_1
XFILLER_27_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20753__RESET_B repeater210/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20902_ _20908_/CLK _20902_/D repeater217/X vssd1 vssd1 vccd1 vccd1 _20902_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_82_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20833_ _20949_/CLK _20833_/D repeater269/X vssd1 vssd1 vccd1 vccd1 _20833_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__13083__B1 _12853_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20764_ _21342_/CLK _20764_/D repeater211/X vssd1 vssd1 vccd1 vccd1 _20764_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20695_ _20697_/CLK _20695_/D repeater196/X vssd1 vssd1 vccd1 vccd1 _20695_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12892__A _13106_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19197__S0 _20130_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_248_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21316_ _21321_/CLK _21316_/D repeater222/X vssd1 vssd1 vccd1 vccd1 _21316_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_123_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17195__A _17195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21247_ _21433_/CLK _21247_/D repeater233/X vssd1 vssd1 vccd1 vccd1 _21247_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__19936__RESET_B repeater251/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20751__CLK _21342_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11000_ _21012_/Q vssd1 vssd1 vccd1 vccd1 _15505_/B sky130_fd_sc_hd__buf_1
X_21178_ _21183_/CLK _21178_/D repeater216/X vssd1 vssd1 vccd1 vccd1 _21178_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_77_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20129_ _21235_/CLK _20129_/D repeater249/X vssd1 vssd1 vccd1 vccd1 _20129_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_89_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13310__A1 _20540_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12951_ _12961_/A vssd1 vssd1 vccd1 vccd1 _12951_/X sky130_fd_sc_hd__buf_1
XANTENNA__10124__A1 _10154_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11902_ _19114_/X _10992_/X _11901_/X vssd1 vssd1 vccd1 vccd1 _21017_/D sky130_fd_sc_hd__a21oi_1
XFILLER_93_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15670_ _19687_/Q _15666_/X _15590_/X _15667_/X vssd1 vssd1 vccd1 vccd1 _19687_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12882_ _20739_/Q _12874_/X _12881_/X _12876_/X vssd1 vssd1 vccd1 vccd1 _20739_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_46_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14621_ _14639_/A vssd1 vssd1 vccd1 vccd1 _14621_/X sky130_fd_sc_hd__clkbuf_2
XPHY_4353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11833_ _21035_/Q _11833_/B vssd1 vssd1 vccd1 vccd1 _11833_/Y sky130_fd_sc_hd__nor2_1
XPHY_4364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13074__B1 _12925_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17340_ _19504_/Q vssd1 vssd1 vccd1 vccd1 _17340_/Y sky130_fd_sc_hd__inv_2
XPHY_4397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10427__A2 _20697_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14552_ _20131_/Q vssd1 vssd1 vccd1 vccd1 _14751_/A sky130_fd_sc_hd__inv_2
XPHY_3663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11764_ _11770_/A vssd1 vssd1 vccd1 vccd1 _11764_/X sky130_fd_sc_hd__buf_1
XPHY_3674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13503_ _20442_/Q _13499_/X _13311_/X _13500_/X vssd1 vssd1 vccd1 vccd1 _20442_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10715_ _10715_/A vssd1 vssd1 vccd1 vccd1 _10715_/Y sky130_fd_sc_hd__inv_2
XFILLER_159_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17271_ _19455_/Q vssd1 vssd1 vccd1 vccd1 _17271_/Y sky130_fd_sc_hd__inv_2
XFILLER_202_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14483_ _14483_/A vssd1 vssd1 vccd1 vccd1 _14483_/Y sky130_fd_sc_hd__inv_2
XPHY_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11695_ _12715_/A vssd1 vssd1 vccd1 vccd1 _17286_/A sky130_fd_sc_hd__buf_1
XPHY_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19010_ _16952_/X _20413_/Q _19019_/S vssd1 vssd1 vccd1 vccd1 _19966_/D sky130_fd_sc_hd__mux2_1
XPHY_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19188__S0 _19280_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16222_ _19426_/Q _16216_/X _16117_/X _16218_/X vssd1 vssd1 vccd1 vccd1 _19426_/D
+ sky130_fd_sc_hd__a22o_1
X_13434_ _20474_/Q _13428_/X _13311_/X _13430_/X vssd1 vssd1 vccd1 vccd1 _20474_/D
+ sky130_fd_sc_hd__a22o_1
X_10646_ _20699_/Q _10685_/A vssd1 vssd1 vccd1 vccd1 _10647_/A sky130_fd_sc_hd__or2_1
XFILLER_173_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17089__B _20700_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16153_ _16159_/A vssd1 vssd1 vccd1 vccd1 _16153_/X sky130_fd_sc_hd__buf_1
Xrebuffer5 rebuffer7/X vssd1 vssd1 vccd1 vccd1 _14954_/A sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_166_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13365_ _13377_/A vssd1 vssd1 vccd1 vccd1 _13365_/X sky130_fd_sc_hd__buf_1
X_10577_ _21341_/Q vssd1 vssd1 vccd1 vccd1 _10577_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21282__RESET_B repeater207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15104_ _15104_/A vssd1 vssd1 vccd1 vccd1 _15104_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12316_ _12316_/A _12369_/A vssd1 vssd1 vccd1 vccd1 _12317_/B sky130_fd_sc_hd__or2_1
X_16084_ _19492_/Q _16080_/X _15869_/X _16082_/X vssd1 vssd1 vccd1 vccd1 _19492_/D
+ sky130_fd_sc_hd__a22o_1
X_13296_ _20548_/Q _13293_/X _13219_/X _13294_/X vssd1 vssd1 vccd1 vccd1 _20548_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_181_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19912_ _21185_/CLK _19912_/D repeater221/X vssd1 vssd1 vccd1 vccd1 _19912_/Q sky130_fd_sc_hd__dfrtp_1
X_15035_ _20067_/Q vssd1 vssd1 vccd1 vccd1 _15081_/A sky130_fd_sc_hd__inv_2
X_12247_ _12428_/A _20519_/Q _12423_/A _20514_/Q vssd1 vssd1 vccd1 vccd1 _12247_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_123_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19843_ _21196_/CLK _19843_/D repeater219/X vssd1 vssd1 vccd1 vccd1 _19843_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__09616__A _20875_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12178_ _20979_/Q _12176_/Y _12139_/X _20341_/Q _12177_/X vssd1 vssd1 vccd1 vccd1
+ _12190_/A sky130_fd_sc_hd__o221a_1
XFILLER_96_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11129_ _21222_/Q vssd1 vssd1 vccd1 vccd1 _16465_/A sky130_fd_sc_hd__inv_2
X_19774_ _19774_/CLK _19774_/D vssd1 vssd1 vccd1 vccd1 _19774_/Q sky130_fd_sc_hd__dfxtp_1
X_16986_ _19974_/Q vssd1 vssd1 vccd1 vccd1 _16986_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_62_HCLK clkbuf_4_14_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _21476_/CLK sky130_fd_sc_hd__clkbuf_16
X_18725_ _17079_/Y _15270_/Y _18908_/S vssd1 vssd1 vccd1 vccd1 _18725_/X sky130_fd_sc_hd__mux2_1
XFILLER_237_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15937_ _15945_/A vssd1 vssd1 vccd1 vccd1 _15937_/X sky130_fd_sc_hd__buf_1
XFILLER_76_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15868_ _19597_/Q _15864_/X _15865_/X _15867_/X vssd1 vssd1 vccd1 vccd1 _19597_/D
+ sky130_fd_sc_hd__a22o_1
X_18656_ _18655_/X _12251_/Y _18910_/S vssd1 vssd1 vccd1 vccd1 _18656_/X sky130_fd_sc_hd__mux2_1
XFILLER_225_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17607_ _21010_/Q _17425_/X _17605_/X _17606_/X _17504_/Y vssd1 vssd1 vccd1 vccd1
+ _17607_/Y sky130_fd_sc_hd__o221ai_4
X_14819_ _14819_/A vssd1 vssd1 vccd1 vccd1 _14823_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__13065__B1 _13003_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_212_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15799_ _15799_/A _15833_/B _16405_/C vssd1 vssd1 vccd1 vccd1 _15807_/A sky130_fd_sc_hd__or3_4
X_18587_ _18586_/X _14896_/Y _18907_/S vssd1 vssd1 vccd1 vccd1 _18587_/X sky130_fd_sc_hd__mux2_1
XFILLER_240_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17538_ _17808_/A vssd1 vssd1 vccd1 vccd1 _17542_/B sky130_fd_sc_hd__buf_4
XFILLER_60_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17469_ _17464_/Y _17387_/X _17465_/Y _17378_/X _17468_/X vssd1 vssd1 vccd1 vccd1
+ _17469_/X sky130_fd_sc_hd__o221a_1
XANTENNA__19179__S0 _19280_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19208_ _17690_/Y _17691_/Y _17692_/Y _17693_/Y _20130_/Q _20131_/Q vssd1 vssd1 vccd1
+ vccd1 _19208_/X sky130_fd_sc_hd__mux4_2
X_20480_ _20480_/CLK _20480_/D repeater183/X vssd1 vssd1 vccd1 vccd1 _20480_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_193_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19139_ _19688_/Q _19376_/Q _19672_/Q _19664_/Q _19285_/S0 _21017_/Q vssd1 vssd1
+ vccd1 vccd1 _19139_/X sky130_fd_sc_hd__mux4_1
XFILLER_192_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18603__S _18928_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21101_ _21429_/CLK _21101_/D repeater229/X vssd1 vssd1 vccd1 vccd1 _21101_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_161_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21032_ _21218_/CLK _21032_/D repeater242/X vssd1 vssd1 vccd1 vccd1 _21032_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__20004__CLK _20004_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09725_ _20159_/Q vssd1 vssd1 vccd1 vccd1 _09725_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11791__A _11794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09656_ _21474_/Q _09643_/X _09655_/X _09646_/X vssd1 vssd1 vccd1 vccd1 _21474_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_227_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16242__B1 _16009_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13056__B1 _12984_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20816_ _21319_/CLK _20816_/D repeater191/X vssd1 vssd1 vccd1 vccd1 _20816_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20747_ _21319_/CLK _20747_/D repeater191/X vssd1 vssd1 vccd1 vccd1 _20747_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13511__A _14264_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10500_ _20686_/Q vssd1 vssd1 vccd1 vccd1 _17981_/A sky130_fd_sc_hd__inv_2
XPHY_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11480_ _11480_/A vssd1 vssd1 vccd1 vccd1 _11480_/X sky130_fd_sc_hd__buf_1
XFILLER_155_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20678_ _21357_/CLK _20678_/D repeater199/X vssd1 vssd1 vccd1 vccd1 _20678_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_12_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10431_ _21291_/Q vssd1 vssd1 vccd1 vccd1 _10767_/A sky130_fd_sc_hd__inv_2
XFILLER_195_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18513__S _18902_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13150_ _13165_/A vssd1 vssd1 vccd1 vccd1 _13150_/X sky130_fd_sc_hd__buf_1
X_10362_ _10366_/A vssd1 vssd1 vccd1 vccd1 _10395_/A sky130_fd_sc_hd__inv_2
XFILLER_163_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12101_ _20968_/Q vssd1 vssd1 vccd1 vccd1 _12321_/A sky130_fd_sc_hd__inv_2
XFILLER_3_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10293_ _10268_/A _20711_/Q _10276_/A _20720_/Q vssd1 vssd1 vccd1 vccd1 _10293_/X
+ sky130_fd_sc_hd__o22a_1
X_13081_ _13099_/A vssd1 vssd1 vccd1 vccd1 _13081_/X sky130_fd_sc_hd__buf_1
X_12032_ _19080_/X _12029_/X _20985_/Q _12030_/X vssd1 vssd1 vccd1 vccd1 _20985_/D
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_85_HCLK clkbuf_4_12_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _21294_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__20675__RESET_B repeater208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_238_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16840_ _19939_/Q _16834_/A _16829_/A _16839_/Y _16836_/Y vssd1 vssd1 vccd1 vccd1
+ _16841_/B sky130_fd_sc_hd__o32a_1
X_16771_ _16774_/B _16770_/Y _16762_/X vssd1 vssd1 vccd1 vccd1 _16771_/X sky130_fd_sc_hd__o21a_1
XFILLER_219_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13295__B1 _13216_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13983_ _13983_/A vssd1 vssd1 vccd1 vccd1 _13983_/Y sky130_fd_sc_hd__inv_2
XFILLER_234_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18510_ _18509_/X _14581_/A _18898_/S vssd1 vssd1 vccd1 vccd1 _18510_/X sky130_fd_sc_hd__mux2_1
X_15722_ _15722_/A _15778_/B _15722_/C vssd1 vssd1 vccd1 vccd1 _15736_/A sky130_fd_sc_hd__or3_4
XFILLER_46_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12934_ _12934_/A vssd1 vssd1 vccd1 vccd1 _12960_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_207_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19490_ _21449_/CLK _19490_/D vssd1 vssd1 vccd1 vccd1 _19490_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18441_ _18440_/X _20512_/Q _18910_/S vssd1 vssd1 vccd1 vccd1 _18441_/X sky130_fd_sc_hd__mux2_1
X_15653_ _15653_/A vssd1 vssd1 vccd1 vccd1 _16311_/A sky130_fd_sc_hd__buf_1
X_12865_ _20747_/Q _12859_/X _12697_/X _12861_/X vssd1 vssd1 vccd1 vccd1 _20747_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_repeater189_A repeater270/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14604_ _14593_/A _14593_/B _14636_/A _14602_/Y vssd1 vssd1 vccd1 vccd1 _20204_/D
+ sky130_fd_sc_hd__a211oi_2
XPHY_4183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18372_ _18371_/X _20522_/Q _18910_/S vssd1 vssd1 vccd1 vccd1 _18372_/X sky130_fd_sc_hd__mux2_1
X_11816_ _11816_/A vssd1 vssd1 vccd1 vccd1 _11816_/Y sky130_fd_sc_hd__inv_2
XPHY_4194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15584_ _15584_/A vssd1 vssd1 vccd1 vccd1 _15584_/X sky130_fd_sc_hd__buf_1
XPHY_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12796_ _20781_/Q _12791_/X _12699_/X _12792_/X vssd1 vssd1 vccd1 vccd1 _20781_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17323_ _17323_/A vssd1 vssd1 vccd1 vccd1 _18065_/A sky130_fd_sc_hd__buf_1
XFILLER_202_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14535_ _20132_/Q vssd1 vssd1 vccd1 vccd1 _14535_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11747_ _16680_/B vssd1 vssd1 vccd1 vccd1 _11748_/B sky130_fd_sc_hd__inv_2
XPHY_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17733__B1 _18703_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21463__RESET_B repeater205/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17254_ _17254_/A vssd1 vssd1 vccd1 vccd1 _17829_/B sky130_fd_sc_hd__inv_2
XPHY_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14466_ _14410_/Y _14378_/A _14465_/X _14421_/Y vssd1 vssd1 vccd1 vccd1 _14467_/C
+ sky130_fd_sc_hd__o31a_1
XPHY_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11678_ _11678_/A _15312_/D vssd1 vssd1 vccd1 vccd1 _11689_/A sky130_fd_sc_hd__or2_2
X_16205_ _19434_/Q _16195_/X _16204_/X _16198_/X vssd1 vssd1 vccd1 vccd1 _19434_/D
+ sky130_fd_sc_hd__a22o_1
X_13417_ _13444_/A vssd1 vssd1 vccd1 vccd1 _13417_/X sky130_fd_sc_hd__buf_1
X_17185_ _20700_/Q _17187_/B vssd1 vssd1 vccd1 vccd1 _17185_/Y sky130_fd_sc_hd__nor2_1
X_10629_ _20740_/Q vssd1 vssd1 vccd1 vccd1 _10629_/Y sky130_fd_sc_hd__inv_2
X_14397_ _21464_/Q vssd1 vssd1 vccd1 vccd1 _14397_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18423__S _18908_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12573__A2 _12566_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16136_ _19468_/Q _16130_/X _16135_/X _16133_/X vssd1 vssd1 vccd1 vccd1 _19468_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09974__B1 _09676_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13348_ _20520_/Q _13345_/X _13209_/X _13346_/X vssd1 vssd1 vccd1 vccd1 _20520_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17547__B _18835_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16067_ _19501_/Q _16064_/X _15758_/X _16066_/X vssd1 vssd1 vccd1 vccd1 _19501_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_142_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13279_ _20557_/Q _13276_/X _13277_/X _13278_/X vssd1 vssd1 vccd1 vccd1 _20557_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15018_ _20080_/Q _15021_/A _15015_/A _14952_/X vssd1 vssd1 vccd1 vccd1 _20080_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__11533__B1 _10892_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19826_ _19835_/CLK _19826_/D vssd1 vssd1 vccd1 vccd1 _19826_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19757_ _19765_/CLK _19757_/D vssd1 vssd1 vccd1 vccd1 _19757_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_244_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16969_ _19970_/Q vssd1 vssd1 vccd1 vccd1 _16970_/A sky130_fd_sc_hd__buf_1
XFILLER_110_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18708_ _17682_/X _19588_/Q _18926_/S vssd1 vssd1 vccd1 vccd1 _18708_/X sky130_fd_sc_hd__mux2_1
XFILLER_204_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19688_ _19811_/CLK _19688_/D vssd1 vssd1 vccd1 vccd1 _19688_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13038__B1 _12957_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18639_ _18638_/X _14099_/A _18904_/S vssd1 vssd1 vccd1 vccd1 _18639_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17972__B1 _18300_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20601_ _20693_/CLK _20601_/D repeater196/X vssd1 vssd1 vccd1 vccd1 _20601_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_177_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20532_ _21366_/CLK _20532_/D repeater265/X vssd1 vssd1 vccd1 vccd1 _20532_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_138_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_opt_1_HCLK_A clkbuf_opt_1_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20463_ _20495_/CLK _20463_/D repeater273/X vssd1 vssd1 vccd1 vccd1 _20463_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__13210__B1 _13209_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18333__S _18667_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10024__B1 _21410_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20394_ _20951_/CLK _20394_/D repeater270/X vssd1 vssd1 vccd1 vccd1 _20394_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_165_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14710__B1 _12857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20898__SET_B repeater212/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21015_ _21121_/CLK _21015_/D repeater238/X vssd1 vssd1 vccd1 vccd1 _21015_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13506__A _14258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09708_ _09812_/B vssd1 vssd1 vccd1 vccd1 _16617_/A sky130_fd_sc_hd__buf_1
XFILLER_28_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10980_ _15505_/C vssd1 vssd1 vccd1 vccd1 _11875_/B sky130_fd_sc_hd__inv_2
XFILLER_243_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09639_ _21479_/Q _09632_/X _09638_/X _09634_/X vssd1 vssd1 vccd1 vccd1 _21479_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13029__B1 _12863_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18508__S _18896_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12650_ _12679_/A vssd1 vssd1 vccd1 vccd1 _12650_/X sky130_fd_sc_hd__buf_1
XPHY_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11601_ _18986_/X _11598_/X _21120_/Q _11600_/X vssd1 vssd1 vccd1 vccd1 _21120_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12581_ _12600_/A vssd1 vssd1 vccd1 vccd1 _12581_/X sky130_fd_sc_hd__buf_1
XPHY_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14320_ _14293_/X _14319_/Y _14293_/X _14319_/Y vssd1 vssd1 vccd1 vccd1 _14324_/C
+ sky130_fd_sc_hd__a2bb2o_1
XPHY_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11532_ _21141_/Q _11527_/X _10889_/X _11529_/X vssd1 vssd1 vccd1 vccd1 _21141_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14251_ _20255_/Q _14246_/X _20254_/Q _14249_/X vssd1 vssd1 vccd1 vccd1 _20255_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11463_ _11481_/A vssd1 vssd1 vccd1 vccd1 _11463_/X sky130_fd_sc_hd__buf_1
XANTENNA__19951__RESET_B repeater270/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13202_ _20592_/Q _13200_/X _12996_/X _13201_/X vssd1 vssd1 vccd1 vccd1 _20592_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_125_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09956__B1 _09685_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17479__C1 _17478_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10414_ _10264_/A _10264_/B _10412_/Y _10375_/X vssd1 vssd1 vccd1 vccd1 _21348_/D
+ sky130_fd_sc_hd__a211oi_2
X_14182_ _14182_/A vssd1 vssd1 vccd1 vccd1 _14182_/Y sky130_fd_sc_hd__inv_2
X_11394_ _19844_/Q vssd1 vssd1 vccd1 vccd1 _16507_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__20856__RESET_B repeater243/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13133_ _13133_/A vssd1 vssd1 vccd1 vccd1 _13133_/X sky130_fd_sc_hd__buf_1
XFILLER_124_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10345_ _21348_/Q _17545_/A _10263_/A _20706_/Q _10344_/X vssd1 vssd1 vccd1 vccd1
+ _10360_/A sky130_fd_sc_hd__o221a_1
X_18990_ _21263_/Q _21115_/Q _18992_/S vssd1 vssd1 vccd1 vccd1 _18990_/X sky130_fd_sc_hd__mux2_1
XFILLER_125_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13504__A1 _20441_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17941_ _17941_/A _17943_/B vssd1 vssd1 vccd1 vccd1 _17941_/Y sky130_fd_sc_hd__nor2_1
XFILLER_140_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_128_HCLK_A clkbuf_4_4_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13064_ _20659_/Q _13060_/X _13001_/X _13061_/X vssd1 vssd1 vccd1 vccd1 _20659_/D
+ sky130_fd_sc_hd__a22o_1
X_10276_ _10276_/A _10391_/A vssd1 vssd1 vccd1 vccd1 _10277_/B sky130_fd_sc_hd__or2_2
XFILLER_155_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12015_ _19069_/X _12010_/X _20996_/Q _12012_/X vssd1 vssd1 vccd1 vccd1 _20996_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19074__S _19908_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_238_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17872_ _18549_/X _17839_/X _18581_/X _17840_/X vssd1 vssd1 vccd1 vccd1 _17872_/X
+ sky130_fd_sc_hd__o22a_1
Xrepeater209 repeater211/X vssd1 vssd1 vccd1 vccd1 repeater209/X sky130_fd_sc_hd__buf_8
X_19611_ _21452_/CLK _19611_/D vssd1 vssd1 vccd1 vccd1 _19611_/Q sky130_fd_sc_hd__dfxtp_1
X_16823_ _16827_/B vssd1 vssd1 vccd1 vccd1 _16830_/B sky130_fd_sc_hd__inv_2
XFILLER_171_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19542_ _19784_/CLK _19542_/D vssd1 vssd1 vccd1 vccd1 _19542_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16754_ _16756_/A _16753_/X _16835_/A vssd1 vssd1 vccd1 vccd1 _16754_/Y sky130_fd_sc_hd__a21oi_1
X_13966_ _20322_/Q _13898_/Y _13899_/Y _13898_/A _13965_/X vssd1 vssd1 vccd1 vccd1
+ _20322_/D sky130_fd_sc_hd__o221a_1
XFILLER_234_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15705_ input38/X vssd1 vssd1 vccd1 vccd1 _16016_/A sky130_fd_sc_hd__clkbuf_2
X_12917_ _20726_/Q _12915_/X _12673_/X _12916_/X vssd1 vssd1 vccd1 vccd1 _20726_/D
+ sky130_fd_sc_hd__a22o_1
X_16685_ _16503_/Y _16510_/A _16684_/A vssd1 vssd1 vccd1 vccd1 _19873_/D sky130_fd_sc_hd__o21a_1
X_19473_ _19521_/CLK _19473_/D vssd1 vssd1 vccd1 vccd1 _19473_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18418__S _18875_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13897_ _13897_/A _13897_/B vssd1 vssd1 vccd1 vccd1 _13898_/A sky130_fd_sc_hd__or2_1
XFILLER_222_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18424_ _18423_/X _15151_/Y _18784_/S vssd1 vssd1 vccd1 vccd1 _18424_/X sky130_fd_sc_hd__mux2_2
XFILLER_61_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12848_ _12874_/A vssd1 vssd1 vccd1 vccd1 _12848_/X sky130_fd_sc_hd__buf_1
X_15636_ _19703_/Q _15632_/X _15590_/X _15633_/X vssd1 vssd1 vccd1 vccd1 _19703_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_222_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15567_ _19738_/Q _15561_/X _15514_/X _15563_/X vssd1 vssd1 vccd1 vccd1 _19738_/D
+ sky130_fd_sc_hd__a22o_1
X_18355_ _18848_/A0 _14108_/Y _18902_/S vssd1 vssd1 vccd1 vccd1 _18355_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13440__B1 _13245_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12779_ _20792_/Q _12777_/X _09630_/X _12778_/X vssd1 vssd1 vccd1 vccd1 _20792_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13151__A input40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14518_ _14518_/A _14518_/B _14518_/C vssd1 vssd1 vccd1 vccd1 _14521_/A sky130_fd_sc_hd__or3_4
X_17306_ _21187_/Q vssd1 vssd1 vccd1 vccd1 _17306_/Y sky130_fd_sc_hd__inv_2
XFILLER_174_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18286_ _18285_/X _10602_/Y _18891_/S vssd1 vssd1 vccd1 vccd1 _18286_/X sky130_fd_sc_hd__mux2_1
X_15498_ _19770_/Q _15492_/X _15421_/X _15494_/X vssd1 vssd1 vccd1 vccd1 _19770_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_159_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14449_ _14437_/X _14449_/B _14449_/C _14449_/D vssd1 vssd1 vccd1 vccd1 _14450_/D
+ sky130_fd_sc_hd__and4b_1
X_17237_ _19639_/Q vssd1 vssd1 vccd1 vccd1 _17237_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18153__S _18907_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17168_ _17164_/Y _17147_/X _17165_/Y _17150_/X _17167_/X vssd1 vssd1 vccd1 vccd1
+ _17168_/X sky130_fd_sc_hd__o221a_1
XANTENNA__18131__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16119_ _16119_/A vssd1 vssd1 vccd1 vccd1 _16119_/X sky130_fd_sc_hd__buf_1
XANTENNA__20597__RESET_B repeater235/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17099_ _19390_/Q vssd1 vssd1 vccd1 vccd1 _17099_/Y sky130_fd_sc_hd__inv_2
X_09990_ _21421_/Q _17038_/A _21421_/Q _17038_/A vssd1 vssd1 vccd1 vccd1 _10017_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_130_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19985__CLK _19985_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19809_ _19820_/CLK _19809_/D vssd1 vssd1 vccd1 vccd1 _19809_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18198__A0 _18848_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20242__SET_B repeater247/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18328__S _18841_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13431__B1 _13429_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13061__A _13073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20515_ _20944_/CLK _20515_/D repeater275/X vssd1 vssd1 vccd1 vccd1 _20515_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_181_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17187__B _17187_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20446_ _20480_/CLK _20446_/D repeater183/X vssd1 vssd1 vccd1 vccd1 _20446_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_180_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18998__S _19026_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18673__A1 _19201_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20377_ _20957_/CLK _20377_/D repeater186/X vssd1 vssd1 vccd1 vccd1 _20377_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_122_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20267__RESET_B repeater263/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10130_ _21391_/Q _10129_/Y _10152_/A _20788_/Q vssd1 vssd1 vccd1 vccd1 _10130_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_79_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13498__B1 _13426_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10061_ _21388_/Q vssd1 vssd1 vccd1 vccd1 _10149_/A sky130_fd_sc_hd__inv_2
XFILLER_87_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13820_ _20177_/Q vssd1 vssd1 vccd1 vccd1 _14567_/A sky130_fd_sc_hd__inv_2
XANTENNA__17931__A _18024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18189__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_115_HCLK clkbuf_opt_3_HCLK/A vssd1 vssd1 vccd1 vccd1 _20470_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_244_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13751_ _20205_/Q vssd1 vssd1 vccd1 vccd1 _14594_/A sky130_fd_sc_hd__inv_2
XFILLER_55_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10963_ _21026_/Q vssd1 vssd1 vccd1 vccd1 _11804_/C sky130_fd_sc_hd__inv_2
XANTENNA__13670__B1 _13553_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18238__S _18242_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12702_ _12708_/A vssd1 vssd1 vccd1 vccd1 _12702_/X sky130_fd_sc_hd__buf_1
XFILLER_204_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16470_ _19298_/Q _16466_/X _16281_/X _16468_/X vssd1 vssd1 vccd1 vccd1 _19298_/D
+ sky130_fd_sc_hd__a22o_1
X_13682_ _20350_/Q _13679_/X _13485_/X _13680_/X vssd1 vssd1 vccd1 vccd1 _20350_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__21055__RESET_B repeater220/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10894_ _10894_/A vssd1 vssd1 vccd1 vccd1 _10894_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_71_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15421_ _15421_/A vssd1 vssd1 vccd1 vccd1 _15421_/X sky130_fd_sc_hd__clkbuf_2
XPHY_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12633_ input31/X _12631_/X _20851_/Q _12632_/X vssd1 vssd1 vccd1 vccd1 _20851_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_43_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18140_ _18139_/X _14427_/Y _18897_/S vssd1 vssd1 vccd1 vccd1 _18140_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15352_ _15429_/A vssd1 vssd1 vccd1 vccd1 _15352_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_156_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12564_ _19984_/D _16527_/B vssd1 vssd1 vccd1 vccd1 _12580_/A sky130_fd_sc_hd__or2b_2
XFILLER_157_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14303_ _20890_/Q _20889_/Q _14303_/C vssd1 vssd1 vccd1 vccd1 _17320_/A sky130_fd_sc_hd__or3_4
XANTENNA__19069__S _19908_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18071_ _20425_/Q vssd1 vssd1 vccd1 vccd1 _18071_/Y sky130_fd_sc_hd__inv_2
X_11515_ input49/X vssd1 vssd1 vccd1 vccd1 _16340_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_156_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15283_ _20482_/Q _15075_/A _18030_/A _20068_/Q _15282_/X vssd1 vssd1 vccd1 vccd1
+ _15284_/D sky130_fd_sc_hd__o221a_1
XPHY_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12495_ _12490_/A _12490_/B _12490_/C vssd1 vssd1 vccd1 vccd1 _12496_/B sky130_fd_sc_hd__o21a_1
XFILLER_200_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17022_ _17022_/A _17023_/B vssd1 vssd1 vccd1 vccd1 _20008_/D sky130_fd_sc_hd__nor2_1
XANTENNA__09929__A0 _20014_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14234_ _19894_/Q _14234_/B vssd1 vssd1 vccd1 vccd1 _14235_/B sky130_fd_sc_hd__or2_1
XANTENNA__13725__A1 _15766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11446_ _21158_/Q _11446_/B vssd1 vssd1 vccd1 vccd1 _11447_/B sky130_fd_sc_hd__or2_1
XFILLER_109_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20835__CLK _20930_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18664__A1 _20594_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14165_ _20538_/Q _14078_/A _20555_/Q _14094_/A vssd1 vssd1 vccd1 vccd1 _14165_/X
+ sky130_fd_sc_hd__o22a_1
X_11377_ _21171_/Q vssd1 vssd1 vccd1 vccd1 _11388_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_124_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13116_ _20630_/Q _13112_/X _12984_/X _13115_/X vssd1 vssd1 vccd1 vccd1 _20630_/D
+ sky130_fd_sc_hd__a22o_1
X_10328_ _21365_/Q _10324_/Y _21361_/Q _17943_/A _10327_/X vssd1 vssd1 vccd1 vccd1
+ _10340_/A sky130_fd_sc_hd__o221a_1
X_14096_ _14096_/A _14182_/A vssd1 vssd1 vccd1 vccd1 _14097_/B sky130_fd_sc_hd__or2_2
X_18973_ _16524_/Y _13177_/Y _18975_/S vssd1 vssd1 vccd1 vccd1 _18973_/X sky130_fd_sc_hd__mux2_1
XFILLER_239_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15626__A _15632_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17924_ _18018_/A vssd1 vssd1 vccd1 vccd1 _17925_/A sky130_fd_sc_hd__buf_1
X_13047_ _13047_/A _13047_/B _13047_/C vssd1 vssd1 vccd1 vccd1 _17209_/A sky130_fd_sc_hd__or3_4
X_10259_ _21344_/Q vssd1 vssd1 vccd1 vccd1 _10260_/A sky130_fd_sc_hd__inv_2
XANTENNA__14530__A _20208_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17855_ _18603_/X _17853_/X _18607_/X _17854_/X vssd1 vssd1 vccd1 vccd1 _17855_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_120_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16806_ _19932_/Q _16801_/A _16805_/Y _16801_/Y vssd1 vssd1 vccd1 vccd1 _16807_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__13146__A input42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17786_ _17784_/Y _17141_/A _17785_/Y _17390_/X vssd1 vssd1 vccd1 vccd1 _17786_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_226_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14998_ _14998_/A vssd1 vssd1 vccd1 vccd1 _15019_/B sky130_fd_sc_hd__buf_1
X_19525_ _20327_/CLK _19525_/D vssd1 vssd1 vccd1 vccd1 _19525_/Q sky130_fd_sc_hd__dfxtp_1
X_16737_ _16737_/A _19995_/Q vssd1 vssd1 vccd1 vccd1 _18931_/S sky130_fd_sc_hd__nor2_1
XFILLER_47_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18148__S _18903_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13949_ _20648_/Q _13971_/C _20648_/Q _13857_/A vssd1 vssd1 vccd1 vccd1 _13949_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_207_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19456_ _21234_/CLK _19456_/D vssd1 vssd1 vccd1 vccd1 _19456_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16668_ _21156_/Q _11444_/B _11445_/B vssd1 vssd1 vccd1 vccd1 _16668_/X sky130_fd_sc_hd__a21bo_1
X_18407_ _18406_/X _15119_/Y _18906_/S vssd1 vssd1 vccd1 vccd1 _18407_/X sky130_fd_sc_hd__mux2_2
XFILLER_62_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15619_ _15619_/A vssd1 vssd1 vccd1 vccd1 _15619_/X sky130_fd_sc_hd__buf_1
XANTENNA__19873__RESET_B repeater225/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13413__B1 _13219_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19387_ _20432_/CLK _19387_/D vssd1 vssd1 vccd1 vccd1 _19387_/Q sky130_fd_sc_hd__dfxtp_1
X_16599_ _21256_/Q vssd1 vssd1 vccd1 vccd1 _16599_/Y sky130_fd_sc_hd__inv_2
XFILLER_203_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18338_ _18337_/X _10779_/A _18898_/S vssd1 vssd1 vccd1 vccd1 _18338_/X sky130_fd_sc_hd__mux2_1
XFILLER_175_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18269_ _18268_/X _21366_/Q _18850_/S vssd1 vssd1 vccd1 vccd1 _18269_/X sky130_fd_sc_hd__mux2_1
XFILLER_175_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20300_ _20316_/CLK _20300_/D repeater197/X vssd1 vssd1 vccd1 vccd1 _20300_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__20707__RESET_B repeater210/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21280_ _21342_/CLK _21280_/D repeater207/X vssd1 vssd1 vccd1 vccd1 _21280_/Q sky130_fd_sc_hd__dfrtp_1
X_20231_ _21484_/CLK _20231_/D repeater203/X vssd1 vssd1 vccd1 vccd1 _20231_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18611__S _18835_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20162_ _21121_/CLK _20162_/D repeater237/X vssd1 vssd1 vccd1 vccd1 _20162_/Q sky130_fd_sc_hd__dfrtp_1
X_09973_ _21419_/Q _09968_/X _09670_/X _09970_/X vssd1 vssd1 vccd1 vccd1 _21419_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_130_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14141__A1 _20551_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20093_ _20496_/CLK _20093_/D repeater273/X vssd1 vssd1 vccd1 vccd1 _20093_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_97_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_138_HCLK clkbuf_4_12_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _21405_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_245_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14444__A2 _14442_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20995_ _21185_/CLK _20995_/D repeater222/X vssd1 vssd1 vccd1 vccd1 _20995_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12895__A _13108_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_213_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15271__A _20482_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18591__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11300_ _11300_/A _20908_/Q _11310_/D _11310_/C vssd1 vssd1 vccd1 vccd1 _11301_/B
+ sky130_fd_sc_hd__or4b_4
XFILLER_126_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12280_ _20509_/Q vssd1 vssd1 vccd1 vccd1 _12280_/Y sky130_fd_sc_hd__inv_2
X_21478_ _21480_/CLK _21478_/D repeater206/X vssd1 vssd1 vccd1 vccd1 _21478_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_112_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11231_ _21194_/Q vssd1 vssd1 vccd1 vccd1 _11241_/A sky130_fd_sc_hd__buf_1
XFILLER_20_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17926__A _18019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20429_ _21001_/CLK _20429_/D repeater190/X vssd1 vssd1 vccd1 vccd1 _20429_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18521__S _18680_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11162_ _21011_/Q _16524_/A _11964_/A vssd1 vssd1 vccd1 vccd1 _15638_/C sky130_fd_sc_hd__or3_4
X_10113_ _10201_/A _20777_/Q _10034_/A _20801_/Q vssd1 vssd1 vccd1 vccd1 _10113_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_121_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15970_ _15978_/A vssd1 vssd1 vccd1 vccd1 _15979_/A sky130_fd_sc_hd__inv_2
X_11093_ _11093_/A _11093_/B vssd1 vssd1 vccd1 vccd1 _11093_/X sky130_fd_sc_hd__and2_1
XFILLER_49_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input32_A HADDR[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19071__A1 _21139_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14921_ _20568_/Q _14853_/A _14919_/Y _20104_/Q _14920_/X vssd1 vssd1 vccd1 vccd1
+ _14933_/A sky130_fd_sc_hd__o221a_1
X_10044_ _21381_/Q vssd1 vssd1 vccd1 vccd1 _10202_/A sky130_fd_sc_hd__inv_2
XFILLER_88_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17640_ _17638_/Y _17639_/X _17044_/Y _17142_/A vssd1 vssd1 vccd1 vccd1 _17640_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_36_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_33_HCLK_A clkbuf_opt_4_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14852_ _20077_/Q vssd1 vssd1 vccd1 vccd1 _15019_/C sky130_fd_sc_hd__inv_2
XFILLER_208_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_96_HCLK_A clkbuf_4_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13803_ _13801_/Y _20201_/Q _13802_/Y _20187_/Q vssd1 vssd1 vccd1 vccd1 _13803_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_223_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14783_ _14783_/A _14783_/B vssd1 vssd1 vccd1 vccd1 _14784_/A sky130_fd_sc_hd__or2_1
X_17571_ _17955_/A vssd1 vssd1 vccd1 vccd1 _17572_/B sky130_fd_sc_hd__clkbuf_2
X_11995_ _20989_/Q _11995_/B vssd1 vssd1 vccd1 vccd1 _11996_/B sky130_fd_sc_hd__or2_1
XANTENNA__13643__B1 _13584_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17909__B1 _18410_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output119_A _18112_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19310_ _20241_/CLK _19310_/D vssd1 vssd1 vccd1 vccd1 _19310_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16522_ _16495_/Y _16632_/B _16686_/A _16498_/A _16494_/X vssd1 vssd1 vccd1 vccd1
+ _16523_/A sky130_fd_sc_hd__o32a_1
X_13734_ _15774_/A _16127_/A _13734_/S vssd1 vssd1 vccd1 vccd1 _20324_/D sky130_fd_sc_hd__mux2_1
XFILLER_244_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10946_ _21027_/Q vssd1 vssd1 vccd1 vccd1 _11804_/D sky130_fd_sc_hd__inv_2
XFILLER_204_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18582__A0 _18845_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19241_ _19237_/X _19238_/X _19239_/X _19240_/X _20132_/Q _20133_/Q vssd1 vssd1 vccd1
+ vccd1 _19241_/X sky130_fd_sc_hd__mux4_2
XFILLER_43_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13665_ _20361_/Q _13659_/X _13545_/X _13662_/X vssd1 vssd1 vccd1 vccd1 _20361_/D
+ sky130_fd_sc_hd__a22o_1
X_16453_ _16459_/A vssd1 vssd1 vccd1 vccd1 _16460_/A sky130_fd_sc_hd__inv_2
XFILLER_188_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_repeater171_A _18891_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09610__C _13383_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10877_ _10877_/A _15312_/A _12605_/A _10908_/B vssd1 vssd1 vccd1 vccd1 _10880_/A
+ sky130_fd_sc_hd__or4_4
XANTENNA_repeater269_A repeater270/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12616_ input11/X _12613_/X _20862_/Q _12614_/X vssd1 vssd1 vccd1 vccd1 _20862_/D
+ sky130_fd_sc_hd__o22a_1
X_15404_ _19810_/Q _15398_/X _15343_/X _15400_/X vssd1 vssd1 vccd1 vccd1 _19810_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13946__A1 _13942_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16384_ _19345_/Q _16378_/X _16204_/X _16380_/X vssd1 vssd1 vccd1 vccd1 _19345_/D
+ sky130_fd_sc_hd__a22o_1
X_19172_ _19704_/Q _19568_/Q _19560_/Q _19552_/Q _19280_/S0 _20122_/Q vssd1 vssd1
+ vccd1 vccd1 _19172_/X sky130_fd_sc_hd__mux4_2
XPHY_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13596_ _20400_/Q _13594_/X _13446_/X _13595_/X vssd1 vssd1 vccd1 vccd1 _20400_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_84_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_19_HCLK clkbuf_4_3_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _21431_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18123_ vssd1 vssd1 vccd1 vccd1 _18123_/HI _18123_/LO sky130_fd_sc_hd__conb_1
X_15335_ _15335_/A _15335_/B _16481_/A vssd1 vssd1 vccd1 vccd1 _15999_/C sky130_fd_sc_hd__or3_4
X_12547_ _20900_/Q _12543_/X _12544_/X _12546_/X vssd1 vssd1 vccd1 vccd1 _20900_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_157_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20189__RESET_B repeater200/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20800__RESET_B repeater255/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15266_ _20477_/Q vssd1 vssd1 vccd1 vccd1 _15266_/Y sky130_fd_sc_hd__inv_2
X_18054_ _20423_/Q vssd1 vssd1 vccd1 vccd1 _18054_/Y sky130_fd_sc_hd__inv_2
XFILLER_145_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12478_ _12476_/A _12476_/B _12445_/A _12476_/Y vssd1 vssd1 vccd1 vccd1 _20928_/D
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__20118__RESET_B repeater247/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17005_ _19978_/Q _17004_/A _17003_/Y _17004_/Y vssd1 vssd1 vccd1 vccd1 _17006_/B
+ sky130_fd_sc_hd__o22a_1
X_14217_ _14103_/X _14216_/A _20268_/Q _14216_/Y _14174_/X vssd1 vssd1 vccd1 vccd1
+ _20268_/D sky130_fd_sc_hd__o221a_1
X_11429_ _11379_/B _11401_/X _11409_/B _11404_/X vssd1 vssd1 vccd1 vccd1 _21174_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_160_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15197_ _15070_/A _15070_/B _15195_/Y _15193_/X vssd1 vssd1 vccd1 vccd1 _20056_/D
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__18431__S _18841_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14148_ _20541_/Q vssd1 vssd1 vccd1 vccd1 _14148_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18956_ _16647_/X _21080_/Q _18962_/S vssd1 vssd1 vccd1 vccd1 _18956_/X sky130_fd_sc_hd__mux2_1
X_14079_ _14079_/A _14103_/A _14216_/A vssd1 vssd1 vccd1 vccd1 _14212_/A sky130_fd_sc_hd__or3_1
XFILLER_112_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17907_ _17907_/A vssd1 vssd1 vccd1 vccd1 _17907_/X sky130_fd_sc_hd__buf_1
X_18887_ _17185_/Y _10723_/B _18899_/S vssd1 vssd1 vccd1 vccd1 _18887_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17838_ _17838_/A _17838_/B vssd1 vssd1 vccd1 vccd1 _17838_/X sky130_fd_sc_hd__or2_2
XFILLER_82_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17769_ _19332_/Q vssd1 vssd1 vccd1 vccd1 _17769_/Y sky130_fd_sc_hd__inv_2
XFILLER_212_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19508_ _20327_/CLK _19508_/D vssd1 vssd1 vccd1 vccd1 _19508_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_212_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20780_ _21147_/CLK _20780_/D repeater215/X vssd1 vssd1 vccd1 vccd1 _20780_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_50_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20959__RESET_B repeater186/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19439_ _20137_/CLK _19439_/D vssd1 vssd1 vccd1 vccd1 _19439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_211_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18606__S _18748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11124__A _21006_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21401_ _21401_/CLK _21401_/D repeater253/X vssd1 vssd1 vccd1 vccd1 _21401_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18876__A1 _16758_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21332_ _21476_/CLK _21332_/D repeater203/X vssd1 vssd1 vccd1 vccd1 _21332_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_108_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19403__CLK _21009_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21263_ _21417_/CLK _21263_/D repeater234/X vssd1 vssd1 vccd1 vccd1 _21263_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_190_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18341__S _18748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20214_ _20220_/CLK _20214_/D repeater202/X vssd1 vssd1 vccd1 vccd1 _20214_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_132_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21194_ _21196_/CLK _21194_/D repeater220/X vssd1 vssd1 vccd1 vccd1 _21194_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_173_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11794__A _11794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09956_ _21426_/Q _09950_/X _09685_/X _09952_/X vssd1 vssd1 vccd1 vccd1 _21426_/D
+ sky130_fd_sc_hd__a22o_1
X_20145_ _21239_/CLK _20145_/D repeater250/X vssd1 vssd1 vccd1 vccd1 _20145_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__19553__CLK _19706_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20076_ _20107_/CLK _20076_/D repeater259/X vssd1 vssd1 vccd1 vccd1 _20076_/Q sky130_fd_sc_hd__dfrtp_4
X_09887_ _20012_/Q _09887_/B vssd1 vssd1 vccd1 vccd1 _09887_/Y sky130_fd_sc_hd__nand2_1
XFILLER_57_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18800__A1 _19246_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10800_ _10777_/A _10777_/B _10795_/X _10797_/Y vssd1 vssd1 vccd1 vccd1 _21301_/D
+ sky130_fd_sc_hd__a211oi_2
XPHY_4557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11780_ _11776_/X _11457_/A _11780_/S vssd1 vssd1 vccd1 vccd1 _11781_/A sky130_fd_sc_hd__mux2_1
XPHY_3823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20978_ _20980_/CLK _20978_/D repeater271/X vssd1 vssd1 vccd1 vccd1 _20978_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_53_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10731_ _20770_/Q vssd1 vssd1 vccd1 vccd1 _10731_/Y sky130_fd_sc_hd__inv_2
XPHY_3867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18516__S _18775_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_241_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20629__RESET_B repeater193/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13450_ _20467_/Q _13444_/X _13449_/X _13447_/X vssd1 vssd1 vccd1 vccd1 _20467_/D
+ sky130_fd_sc_hd__a22o_1
X_10662_ _10662_/A _10679_/A vssd1 vssd1 vccd1 vccd1 _10663_/B sky130_fd_sc_hd__or2_1
XFILLER_185_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12401_ _12428_/A _12427_/A _12420_/A _12419_/A vssd1 vssd1 vccd1 vccd1 _12403_/C
+ sky130_fd_sc_hd__or4_4
X_13381_ _20499_/Q _13377_/X _13171_/X _13378_/X vssd1 vssd1 vccd1 vccd1 _20499_/D
+ sky130_fd_sc_hd__a22o_1
X_10593_ _20747_/Q vssd1 vssd1 vccd1 vccd1 _10593_/Y sky130_fd_sc_hd__inv_2
X_15120_ _20461_/Q _15086_/A _15119_/Y _20072_/Q vssd1 vssd1 vccd1 vccd1 _15120_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__20282__RESET_B repeater264/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12332_ _12332_/A _12339_/A vssd1 vssd1 vccd1 vccd1 _12333_/B sky130_fd_sc_hd__or2_2
XFILLER_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20211__RESET_B repeater203/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15051_ _20051_/Q vssd1 vssd1 vccd1 vccd1 _15066_/A sky130_fd_sc_hd__inv_2
X_12263_ _20514_/Q vssd1 vssd1 vccd1 vccd1 _12263_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18619__A1 _20288_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18251__S _18907_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14002_ _14002_/A vssd1 vssd1 vccd1 vccd1 _14002_/Y sky130_fd_sc_hd__inv_2
X_11214_ _11226_/A vssd1 vssd1 vccd1 vccd1 _11214_/X sky130_fd_sc_hd__buf_1
XFILLER_141_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18095__A2 _17862_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12194_ _20363_/Q vssd1 vssd1 vccd1 vccd1 _12194_/Y sky130_fd_sc_hd__inv_2
X_18810_ _18809_/X _10756_/A _18880_/S vssd1 vssd1 vccd1 vccd1 _18810_/X sky130_fd_sc_hd__mux2_2
X_11145_ _21220_/Q vssd1 vssd1 vccd1 vccd1 _15609_/A sky130_fd_sc_hd__buf_1
Xoutput84 _17911_/Y vssd1 vssd1 vccd1 vccd1 HRDATA[14] sky130_fd_sc_hd__clkbuf_2
X_19790_ _19820_/CLK _19790_/D vssd1 vssd1 vccd1 vccd1 _19790_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17842__A2 _18024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput95 _18042_/X vssd1 vssd1 vccd1 vccd1 HRDATA[24] sky130_fd_sc_hd__clkbuf_2
X_18741_ _17547_/Y _16902_/A _18875_/S vssd1 vssd1 vccd1 vccd1 _18741_/X sky130_fd_sc_hd__mux2_2
XFILLER_89_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15953_ _15985_/A _16325_/B _16229_/C vssd1 vssd1 vccd1 vccd1 _15961_/A sky130_fd_sc_hd__or3_4
X_11076_ _11101_/A vssd1 vssd1 vccd1 vccd1 _11076_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_237_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19082__S _19908_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10678__B1 _10677_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14904_ _14903_/Y _20085_/Q _20574_/Q _15005_/A vssd1 vssd1 vccd1 vccd1 _14904_/X
+ sky130_fd_sc_hd__o22a_1
X_10027_ _10898_/A _21409_/Q _10028_/S vssd1 vssd1 vccd1 vccd1 _21409_/D sky130_fd_sc_hd__mux2_1
XFILLER_237_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18672_ _17776_/Y _09895_/Y _20870_/Q vssd1 vssd1 vccd1 vccd1 _18672_/X sky130_fd_sc_hd__mux2_1
XFILLER_248_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15884_ _15884_/A _17153_/A vssd1 vssd1 vccd1 vccd1 _16485_/A sky130_fd_sc_hd__or2_4
X_17623_ _19330_/Q vssd1 vssd1 vccd1 vccd1 _17623_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14835_ _14835_/A vssd1 vssd1 vccd1 vccd1 _14963_/D sky130_fd_sc_hd__buf_1
XFILLER_29_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13616__B1 _13553_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13424__A input42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17554_ _21060_/Q vssd1 vssd1 vccd1 vccd1 _17554_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14766_ _14536_/X _14765_/Y _14536_/X _14765_/Y vssd1 vssd1 vccd1 vccd1 _14769_/C
+ sky130_fd_sc_hd__a2bb2o_1
X_11978_ _11978_/A _11978_/B vssd1 vssd1 vccd1 vccd1 _11978_/Y sky130_fd_sc_hd__nor2_1
XFILLER_205_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16505_ _16597_/A _16505_/B vssd1 vssd1 vccd1 vccd1 _16505_/X sky130_fd_sc_hd__or2_1
XFILLER_189_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10929_ _21038_/Q vssd1 vssd1 vccd1 vccd1 _11815_/A sky130_fd_sc_hd__inv_2
X_13717_ _16515_/A _13717_/B _13717_/C vssd1 vssd1 vccd1 vccd1 _13727_/A sky130_fd_sc_hd__or3_4
X_17485_ _19642_/Q vssd1 vssd1 vccd1 vccd1 _17485_/Y sky130_fd_sc_hd__inv_2
X_14697_ _18246_/X _14696_/X _20163_/Q _14692_/X vssd1 vssd1 vccd1 vccd1 _20163_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_205_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18426__S _18928_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19224_ _17596_/Y _17597_/Y _17598_/Y _17599_/Y _19275_/S0 _21004_/Q vssd1 vssd1
+ vccd1 vccd1 _19224_/X sky130_fd_sc_hd__mux4_2
XFILLER_20_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16436_ _16442_/A vssd1 vssd1 vccd1 vccd1 _16436_/X sky130_fd_sc_hd__buf_1
XFILLER_158_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13648_ _20370_/Q _13645_/X _13509_/X _13646_/X vssd1 vssd1 vccd1 vccd1 _20370_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_20_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19155_ _19659_/Q _19651_/Q _19635_/Q _19819_/Q _19285_/S0 _21017_/Q vssd1 vssd1
+ vccd1 vccd1 _19155_/X sky130_fd_sc_hd__mux4_2
X_16367_ _19355_/Q _16363_/X _16200_/X _16365_/X vssd1 vssd1 vccd1 vccd1 _19355_/D
+ sky130_fd_sc_hd__a22o_1
X_13579_ _20409_/Q _13573_/X _13426_/X _13575_/X vssd1 vssd1 vccd1 vccd1 _20409_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_158_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14255__A _20251_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18106_ hold9/A _19291_/Q vssd1 vssd1 vccd1 vccd1 _19982_/D sky130_fd_sc_hd__or2_1
X_15318_ _15318_/A vssd1 vssd1 vccd1 vccd1 _15320_/B sky130_fd_sc_hd__inv_2
X_19086_ _21047_/Q _21060_/Q _19872_/Q vssd1 vssd1 vccd1 vccd1 _19086_/X sky130_fd_sc_hd__mux2_1
X_16298_ _16305_/A vssd1 vssd1 vccd1 vccd1 _16298_/X sky130_fd_sc_hd__buf_1
XFILLER_184_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18037_ _20421_/Q _18084_/B vssd1 vssd1 vccd1 vccd1 _18037_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__18161__S _18669_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15249_ _15246_/Y _20069_/Q _17807_/A _20052_/Q _15248_/X vssd1 vssd1 vccd1 vccd1
+ _15250_/D sky130_fd_sc_hd__o221a_1
XFILLER_132_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09810_ _09806_/A _09806_/B _21454_/Q _09809_/X vssd1 vssd1 vccd1 vccd1 _21454_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_87_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19988_ _21196_/CLK _19988_/D repeater218/X vssd1 vssd1 vccd1 vccd1 _19988_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_98_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09741_ _09739_/X _20146_/Q _21226_/Q _09740_/Y vssd1 vssd1 vccd1 vccd1 _09742_/D
+ sky130_fd_sc_hd__o22a_1
X_18939_ _16706_/X _21137_/Q _18946_/S vssd1 vssd1 vccd1 vccd1 _18939_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19130__S1 _21017_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09672_ _09672_/A vssd1 vssd1 vccd1 vccd1 _15329_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_82_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20901_ _21196_/CLK _20901_/D repeater217/X vssd1 vssd1 vccd1 vccd1 _20901_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_36_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20832_ _21372_/CLK _20832_/D repeater268/X vssd1 vssd1 vccd1 vccd1 _20832_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_82_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13083__A1 _20648_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20793__RESET_B repeater252/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20763_ _21342_/CLK _20763_/D repeater211/X vssd1 vssd1 vccd1 vccd1 _20763_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18336__S _18896_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16645__A _16663_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20722__RESET_B repeater264/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20694_ _20697_/CLK _20694_/D repeater193/X vssd1 vssd1 vccd1 vccd1 _20694_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_50_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19197__S1 _20131_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18849__A1 _13942_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_248_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21315_ _21319_/CLK _21315_/D repeater222/X vssd1 vssd1 vccd1 vccd1 _21315_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__15532__B1 _15450_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21246_ _21433_/CLK _21246_/D repeater236/X vssd1 vssd1 vccd1 vccd1 _21246_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_117_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13509__A _14262_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21177_ _21183_/CLK _21177_/D repeater216/X vssd1 vssd1 vccd1 vccd1 _21177_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_104_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20128_ _21273_/CLK _20128_/D repeater245/X vssd1 vssd1 vccd1 vccd1 _20128_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_77_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09939_ _11654_/A _17231_/A vssd1 vssd1 vccd1 vccd1 _10026_/B sky130_fd_sc_hd__or2_2
XFILLER_219_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15724__A input67/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12950_ _14258_/A vssd1 vssd1 vccd1 vccd1 _12950_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__19905__RESET_B repeater217/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_219_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20059_ _20066_/CLK _20059_/D repeater281/X vssd1 vssd1 vccd1 vccd1 _20059_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_46_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18785__A0 _18784_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10124__A2 _20790_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11901_ _11896_/A _10991_/B _10991_/A vssd1 vssd1 vccd1 vccd1 _11901_/X sky130_fd_sc_hd__o21a_1
XFILLER_245_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12881_ _13171_/A vssd1 vssd1 vccd1 vccd1 _12881_/X sky130_fd_sc_hd__buf_2
XPHY_4310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14620_ _20195_/Q _14619_/Y _14610_/X _14585_/B vssd1 vssd1 vccd1 vccd1 _20195_/D
+ sky130_fd_sc_hd__o211a_1
X_11832_ _11832_/A vssd1 vssd1 vccd1 vccd1 _11833_/B sky130_fd_sc_hd__inv_2
XPHY_4354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14271__B1 _13712_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14551_ _15832_/A _15798_/B _15902_/B vssd1 vssd1 vccd1 vccd1 _14553_/A sky130_fd_sc_hd__o21ai_2
X_11763_ _19872_/Q _11763_/B vssd1 vssd1 vccd1 vccd1 _21052_/D sky130_fd_sc_hd__or2_1
XPHY_3653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10714_ _10706_/A _10706_/B _10711_/Y _10677_/X vssd1 vssd1 vccd1 vccd1 _21318_/D
+ sky130_fd_sc_hd__a211oi_2
XPHY_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13502_ _20443_/Q _13499_/X _13432_/X _13500_/X vssd1 vssd1 vccd1 vccd1 _20443_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14482_ _14460_/B _14372_/B _14480_/Y _14474_/X vssd1 vssd1 vccd1 vccd1 _20229_/D
+ sky130_fd_sc_hd__a211oi_2
XPHY_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17270_ _19439_/Q vssd1 vssd1 vccd1 vccd1 _17270_/Y sky130_fd_sc_hd__inv_2
XFILLER_198_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11694_ _21080_/Q _11689_/X _11573_/X _11690_/X vssd1 vssd1 vccd1 vccd1 _21080_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19288__D _21185_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19188__S1 _20122_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13433_ _20475_/Q _13428_/X _13432_/X _13430_/X vssd1 vssd1 vccd1 vccd1 _20475_/D
+ sky130_fd_sc_hd__a22o_1
X_16221_ _19427_/Q _16216_/X _16115_/X _16218_/X vssd1 vssd1 vccd1 vccd1 _19427_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_201_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10645_ _10677_/A vssd1 vssd1 vccd1 vccd1 _10729_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_174_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16152_ _16158_/A vssd1 vssd1 vccd1 vccd1 _16159_/A sky130_fd_sc_hd__inv_2
X_13364_ _20510_/Q _13358_/X _13148_/X _13360_/X vssd1 vssd1 vccd1 vccd1 _20510_/D
+ sky130_fd_sc_hd__a22o_1
X_10576_ _10576_/A vssd1 vssd1 vccd1 vccd1 _10649_/A sky130_fd_sc_hd__inv_2
XFILLER_154_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrebuffer6 _14950_/A vssd1 vssd1 vccd1 vccd1 rebuffer6/X sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_127_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19077__S _19908_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12315_ _12315_/A _12315_/B vssd1 vssd1 vccd1 vccd1 _12369_/A sky130_fd_sc_hd__or2_1
X_15103_ _20462_/Q vssd1 vssd1 vccd1 vccd1 _15103_/Y sky130_fd_sc_hd__inv_2
X_16083_ _19493_/Q _16080_/X _15865_/X _16082_/X vssd1 vssd1 vccd1 vccd1 _19493_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_181_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13295_ _20549_/Q _13293_/X _13216_/X _13294_/X vssd1 vssd1 vccd1 vccd1 _20549_/D
+ sky130_fd_sc_hd__a22o_1
X_19911_ _21055_/CLK _19911_/D repeater220/X vssd1 vssd1 vccd1 vccd1 _19911_/Q sky130_fd_sc_hd__dfrtp_1
X_15034_ _20068_/Q vssd1 vssd1 vccd1 vccd1 _15104_/A sky130_fd_sc_hd__inv_2
XFILLER_108_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12246_ _20934_/Q vssd1 vssd1 vccd1 vccd1 _12423_/A sky130_fd_sc_hd__inv_2
X_19842_ _21134_/CLK _19842_/D repeater212/X vssd1 vssd1 vccd1 vccd1 _19842_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__10899__B1 _10898_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12177_ _12332_/A _20361_/Q _12073_/X _12147_/Y vssd1 vssd1 vccd1 vccd1 _12177_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_111_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11128_ _11131_/B vssd1 vssd1 vccd1 vccd1 _11128_/X sky130_fd_sc_hd__buf_1
X_19773_ _19789_/CLK _19773_/D vssd1 vssd1 vccd1 vccd1 _19773_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16985_ _19973_/Q _16980_/Y _16983_/Y _16980_/A _16984_/X vssd1 vssd1 vccd1 vccd1
+ _16985_/X sky130_fd_sc_hd__o221a_1
X_18724_ _18723_/X _14075_/A _18850_/S vssd1 vssd1 vccd1 vccd1 _18724_/X sky130_fd_sc_hd__mux2_1
X_11059_ _11059_/A _11085_/A vssd1 vssd1 vccd1 vccd1 _11080_/A sky130_fd_sc_hd__or2_1
X_15936_ _15943_/A vssd1 vssd1 vccd1 vccd1 _15945_/A sky130_fd_sc_hd__inv_2
XANTENNA__10115__A2 _20777_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_237_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18655_ _18654_/X _12194_/Y _18787_/S vssd1 vssd1 vccd1 vccd1 _18655_/X sky130_fd_sc_hd__mux2_1
XFILLER_92_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_237_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15867_ _15877_/A vssd1 vssd1 vccd1 vccd1 _15867_/X sky130_fd_sc_hd__buf_1
XFILLER_18_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13154__A input39/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17606_ _11940_/A _17348_/X _21010_/Q _17425_/X vssd1 vssd1 vccd1 vccd1 _17606_/X
+ sky130_fd_sc_hd__a22o_1
X_14818_ _20112_/Q _20113_/Q _14818_/S vssd1 vssd1 vccd1 vccd1 _20113_/D sky130_fd_sc_hd__mux2_1
XFILLER_240_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18586_ _18585_/X _15127_/Y _18784_/S vssd1 vssd1 vccd1 vccd1 _18586_/X sky130_fd_sc_hd__mux2_2
XFILLER_92_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15798_ _15832_/A _15798_/B _16484_/B vssd1 vssd1 vccd1 vccd1 _16405_/C sky130_fd_sc_hd__or3_4
XFILLER_205_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17537_ _17777_/A _20113_/Q vssd1 vssd1 vccd1 vccd1 _17537_/Y sky130_fd_sc_hd__nand2_1
X_14749_ _14747_/A _14747_/B _14747_/Y vssd1 vssd1 vccd1 vccd1 _20134_/D sky130_fd_sc_hd__a21oi_1
XFILLER_233_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18156__S _18617_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12993__A input58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17468_ _17466_/Y _14256_/A _17467_/Y _17390_/X vssd1 vssd1 vccd1 vccd1 _17468_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_177_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20133__RESET_B repeater249/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19207_ _17686_/Y _17687_/Y _17688_/Y _17689_/Y _20130_/Q _20131_/Q vssd1 vssd1 vccd1
+ vccd1 _19207_/X sky130_fd_sc_hd__mux4_1
X_16419_ _16419_/A _16419_/B _16419_/C vssd1 vssd1 vccd1 vccd1 _16427_/A sky130_fd_sc_hd__or3_4
XANTENNA__19179__S1 _20122_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13601__B _13601_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17399_ _18834_/X _17315_/X _18802_/X _17844_/A vssd1 vssd1 vccd1 vccd1 _17399_/X
+ sky130_fd_sc_hd__o22a_2
X_19138_ _19760_/Q _19752_/Q _19744_/Q _19736_/Q _19285_/S0 _21017_/Q vssd1 vssd1
+ vccd1 vccd1 _19138_/X sky130_fd_sc_hd__mux4_2
XFILLER_192_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18700__A0 _18699_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19069_ _16734_/X _21141_/Q _19908_/D vssd1 vssd1 vccd1 vccd1 _19069_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21100_ _21429_/CLK _21100_/D repeater229/X vssd1 vssd1 vccd1 vccd1 _21100_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_105_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13329__A _13329_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21031_ _21207_/CLK _21031_/D repeater242/X vssd1 vssd1 vccd1 vccd1 _21031_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_234_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13048__B _17209_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09724_ _21239_/Q vssd1 vssd1 vccd1 vccd1 _09724_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15544__A _15657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18767__A0 _17281_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20974__RESET_B repeater278/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09655_ _12860_/A vssd1 vssd1 vccd1 vccd1 _09655_/X sky130_fd_sc_hd__buf_4
XFILLER_227_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20903__RESET_B repeater217/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_227_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_242_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20815_ _21141_/CLK _20815_/D repeater212/X vssd1 vssd1 vccd1 vccd1 _20815_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_24_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20746_ _21342_/CLK _20746_/D repeater207/X vssd1 vssd1 vccd1 vccd1 _20746_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20677_ _21480_/CLK _20677_/D repeater208/X vssd1 vssd1 vccd1 vccd1 _20677_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_195_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10430_ _20685_/Q vssd1 vssd1 vccd1 vccd1 _10430_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10361_ _10361_/A _10361_/B _10361_/C _10361_/D vssd1 vssd1 vccd1 vccd1 _10366_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_128_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12100_ _20395_/Q vssd1 vssd1 vccd1 vccd1 _12100_/Y sky130_fd_sc_hd__inv_2
XFILLER_163_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13080_ _13080_/A vssd1 vssd1 vccd1 vccd1 _13099_/A sky130_fd_sc_hd__buf_1
X_10292_ _20712_/Q vssd1 vssd1 vccd1 vccd1 _10292_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21009__RESET_B repeater235/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12031_ _19079_/X _12029_/X _20986_/Q _12030_/X vssd1 vssd1 vccd1 vccd1 _20986_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_2_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21229_ _21235_/CLK _21229_/D repeater249/X vssd1 vssd1 vccd1 vccd1 _21229_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_2_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15454__A _15661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16770_ _16770_/A _16770_/B vssd1 vssd1 vccd1 vccd1 _16770_/Y sky130_fd_sc_hd__nor2_1
XFILLER_46_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13982_ _20317_/Q _13977_/C _13969_/X _13979_/A vssd1 vssd1 vccd1 vccd1 _20317_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_219_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15721_ _19662_/Q _15716_/X _15706_/X _15717_/X vssd1 vssd1 vccd1 vccd1 _19662_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_234_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12933_ _20719_/Q _12924_/X _12932_/X _12926_/X vssd1 vssd1 vccd1 vccd1 _20719_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_219_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18440_ _17895_/Y _20346_/Q _18909_/S vssd1 vssd1 vccd1 vccd1 _18440_/X sky130_fd_sc_hd__mux2_1
X_15652_ _19694_/Q _15647_/X _15487_/X _15648_/X vssd1 vssd1 vccd1 vccd1 _19694_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_73_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12864_ _20748_/Q _12859_/X _12863_/X _12861_/X vssd1 vssd1 vccd1 vccd1 _20748_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14603_ _20205_/Q _14602_/Y _14599_/X _14595_/B vssd1 vssd1 vccd1 vccd1 _20205_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_4173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18371_ _18029_/Y _20356_/Q _18909_/S vssd1 vssd1 vccd1 vccd1 _18371_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11815_ _11815_/A _11822_/A vssd1 vssd1 vccd1 vccd1 _11815_/X sky130_fd_sc_hd__or2_1
XPHY_4184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output101_A _17406_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15583_ _19730_/Q _15576_/X _15582_/X _15578_/X vssd1 vssd1 vccd1 vccd1 _19730_/D
+ sky130_fd_sc_hd__a22o_1
X_12795_ _20782_/Q _12791_/X _12697_/X _12792_/X vssd1 vssd1 vccd1 vccd1 _20782_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17322_ _18850_/X _17211_/A _18853_/X _17319_/X _17321_/X vssd1 vssd1 vccd1 vccd1
+ _17322_/X sky130_fd_sc_hd__o221a_2
X_11746_ _19999_/Q vssd1 vssd1 vccd1 vccd1 _16680_/B sky130_fd_sc_hd__clkbuf_2
X_14534_ _14663_/A vssd1 vssd1 vccd1 vccd1 _14534_/X sky130_fd_sc_hd__buf_1
XPHY_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09671__B1 _09670_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17253_ _19583_/Q vssd1 vssd1 vccd1 vccd1 _17253_/Y sky130_fd_sc_hd__inv_2
XPHY_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14465_ _14465_/A _14465_/B _14465_/C _14464_/X vssd1 vssd1 vccd1 vccd1 _14465_/X
+ sky130_fd_sc_hd__or4b_4
XFILLER_169_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11677_ _11726_/B vssd1 vssd1 vccd1 vccd1 _15312_/D sky130_fd_sc_hd__clkbuf_2
XPHY_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18704__S _18928_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12558__B1 _11743_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16204_ _21450_/Q vssd1 vssd1 vccd1 vccd1 _16204_/X sky130_fd_sc_hd__buf_1
X_10628_ _10664_/A _20763_/Q _21328_/Q _10626_/Y _10627_/X vssd1 vssd1 vccd1 vccd1
+ _10638_/B sky130_fd_sc_hd__o221a_1
X_13416_ _13416_/A vssd1 vssd1 vccd1 vccd1 _13444_/A sky130_fd_sc_hd__clkbuf_2
X_14396_ _21473_/Q vssd1 vssd1 vccd1 vccd1 _14396_/Y sky130_fd_sc_hd__inv_2
X_17184_ _21343_/Q vssd1 vssd1 vccd1 vccd1 _17184_/Y sky130_fd_sc_hd__inv_2
XFILLER_190_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16135_ _21452_/Q vssd1 vssd1 vccd1 vccd1 _16135_/X sky130_fd_sc_hd__clkbuf_2
X_13347_ _20521_/Q _13345_/X _13287_/X _13346_/X vssd1 vssd1 vccd1 vccd1 _20521_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11230__B1 _10900_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10559_ _21322_/Q vssd1 vssd1 vccd1 vccd1 _10651_/A sky130_fd_sc_hd__inv_2
XFILLER_155_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13278_ _13294_/A vssd1 vssd1 vccd1 vccd1 _13278_/X sky130_fd_sc_hd__buf_1
X_16066_ _16072_/A vssd1 vssd1 vccd1 vccd1 _16066_/X sky130_fd_sc_hd__buf_1
XFILLER_170_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12229_ _20519_/Q vssd1 vssd1 vccd1 vccd1 _12229_/Y sky130_fd_sc_hd__inv_2
X_15017_ _15017_/A vssd1 vssd1 vccd1 vccd1 _15021_/A sky130_fd_sc_hd__inv_2
XFILLER_151_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19825_ _19835_/CLK _19825_/D vssd1 vssd1 vccd1 vccd1 _19825_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19756_ _19813_/CLK _19756_/D vssd1 vssd1 vccd1 vccd1 _19756_/Q sky130_fd_sc_hd__dfxtp_1
X_16968_ _16965_/Y _16966_/Y _16967_/X vssd1 vssd1 vccd1 vccd1 _16968_/X sky130_fd_sc_hd__o21a_1
XFILLER_96_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18707_ _17683_/X _21203_/Q _18928_/S vssd1 vssd1 vccd1 vccd1 _18707_/X sky130_fd_sc_hd__mux2_1
X_15919_ _15919_/A _16325_/B _16325_/C vssd1 vssd1 vccd1 vccd1 _15927_/A sky130_fd_sc_hd__or3_4
XFILLER_37_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19687_ _19765_/CLK _19687_/D vssd1 vssd1 vccd1 vccd1 _19687_/Q sky130_fd_sc_hd__dfxtp_1
X_16899_ _16902_/B _16897_/X _16898_/X vssd1 vssd1 vccd1 vccd1 _16899_/X sky130_fd_sc_hd__o21a_1
XFILLER_224_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18638_ _18637_/X _13944_/Y _18849_/S vssd1 vssd1 vccd1 vccd1 _18638_/X sky130_fd_sc_hd__mux2_1
XFILLER_224_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19764__CLK _19765_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_212_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18569_ _18568_/X _10623_/Y _18891_/S vssd1 vssd1 vccd1 vccd1 _18569_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_220_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20600_ _20622_/CLK _20600_/D repeater196/X vssd1 vssd1 vccd1 vccd1 _20600_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_220_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20531_ _21366_/CLK _20531_/D repeater265/X vssd1 vssd1 vccd1 vccd1 _20531_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18614__S _18667_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12549__B1 _12548_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20462_ _20944_/CLK _20462_/D repeater274/X vssd1 vssd1 vccd1 vccd1 _20462_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__11221__B1 _10884_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20393_ _20951_/CLK _20393_/D repeater272/X vssd1 vssd1 vccd1 vccd1 _20393_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__10971__A _11800_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21173__RESET_B repeater220/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20121__CLK _21452_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21014_ _21121_/CLK _21014_/D repeater238/X vssd1 vssd1 vccd1 vccd1 _21014_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_248_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12898__A _12898_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17660__B1 _18735_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09707_ _09780_/A _09783_/A vssd1 vssd1 vccd1 vccd1 _09812_/B sky130_fd_sc_hd__or2_1
XFILLER_244_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12485__C1 _12445_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09638_ input45/X vssd1 vssd1 vccd1 vccd1 _09638_/X sky130_fd_sc_hd__buf_4
XFILLER_243_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20055__RESET_B repeater281/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12788__B1 _09645_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11600_ _11605_/A vssd1 vssd1 vccd1 vccd1 _11600_/X sky130_fd_sc_hd__buf_1
XFILLER_212_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12580_ _12580_/A vssd1 vssd1 vccd1 vccd1 _12600_/A sky130_fd_sc_hd__clkbuf_2
XPHY_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09653__B1 _09652_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19260__S0 _20130_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11531_ _21142_/Q _11527_/X _10886_/X _11529_/X vssd1 vssd1 vccd1 vccd1 _21142_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20729_ _21375_/CLK _20729_/D repeater257/X vssd1 vssd1 vccd1 vccd1 _20729_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18524__S _18910_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14250_ _20256_/Q _14246_/X _19907_/Q _14249_/X vssd1 vssd1 vccd1 vccd1 _20256_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11462_ _11462_/A vssd1 vssd1 vccd1 vccd1 _11481_/A sky130_fd_sc_hd__inv_2
XPHY_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_52_HCLK clkbuf_4_14_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _21141_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13201_ _13217_/A vssd1 vssd1 vccd1 vccd1 _13201_/X sky130_fd_sc_hd__buf_1
XFILLER_137_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17479__B1 _18785_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11212__B1 _09652_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10413_ _21349_/Q _10412_/Y _10266_/B _10381_/X vssd1 vssd1 vccd1 vccd1 _21349_/D
+ sky130_fd_sc_hd__o211a_1
X_14181_ _14097_/A _14097_/B _14179_/Y _14215_/B vssd1 vssd1 vccd1 vccd1 _20287_/D
+ sky130_fd_sc_hd__a211oi_2
X_11393_ _11408_/A vssd1 vssd1 vccd1 vccd1 _11393_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13132_ _13132_/A vssd1 vssd1 vccd1 vccd1 _13132_/X sky130_fd_sc_hd__buf_1
XANTENNA__11696__B _15312_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input62_A HWDATA[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10344_ _21356_/Q _10342_/Y _21364_/Q _17982_/A vssd1 vssd1 vccd1 vccd1 _10344_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_155_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13063_ _20660_/Q _13060_/X _12999_/X _13061_/X vssd1 vssd1 vccd1 vccd1 _20660_/D
+ sky130_fd_sc_hd__a22o_1
X_17940_ _17940_/A _17943_/B vssd1 vssd1 vccd1 vccd1 _17940_/Y sky130_fd_sc_hd__nor2_1
X_10275_ _10275_/A _10275_/B vssd1 vssd1 vccd1 vccd1 _10391_/A sky130_fd_sc_hd__or2_1
XANTENNA__19920__RESET_B repeater212/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12014_ _19068_/X _12010_/X _20997_/Q _12012_/X vssd1 vssd1 vccd1 vccd1 _20997_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12712__B1 _11743_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17871_ _18572_/X _17856_/X _18559_/X _17569_/X _17870_/X vssd1 vssd1 vccd1 vccd1
+ _17871_/X sky130_fd_sc_hd__o221a_1
Xclkbuf_4_6_0_HCLK clkbuf_4_7_0_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_6_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_238_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19610_ _19626_/CLK _19610_/D vssd1 vssd1 vccd1 vccd1 _19610_/Q sky130_fd_sc_hd__dfxtp_1
X_16822_ _16822_/A _19936_/Q _16822_/C vssd1 vssd1 vccd1 vccd1 _16827_/B sky130_fd_sc_hd__or3_1
XFILLER_238_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19541_ _19789_/CLK _19541_/D vssd1 vssd1 vccd1 vccd1 _19541_/Q sky130_fd_sc_hd__dfxtp_1
X_16753_ _16753_/A _16753_/B vssd1 vssd1 vccd1 vccd1 _16753_/X sky130_fd_sc_hd__or2_1
X_13965_ _13987_/A vssd1 vssd1 vccd1 vccd1 _13965_/X sky130_fd_sc_hd__buf_1
XFILLER_171_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15704_ _19671_/Q _15696_/X _15703_/X _15698_/X vssd1 vssd1 vccd1 vccd1 _19671_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17403__B1 _18819_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19472_ _19813_/CLK _19472_/D vssd1 vssd1 vccd1 vccd1 _19472_/Q sky130_fd_sc_hd__dfxtp_1
X_12916_ _12926_/A vssd1 vssd1 vccd1 vccd1 _12916_/X sky130_fd_sc_hd__buf_1
XFILLER_234_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16684_ _16684_/A _18947_/X vssd1 vssd1 vccd1 vccd1 _19874_/D sky130_fd_sc_hd__and2_1
XFILLER_206_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20764__CLK _21342_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13896_ _20320_/Q _13896_/B vssd1 vssd1 vccd1 vccd1 _13897_/B sky130_fd_sc_hd__nand2_1
XFILLER_61_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18423_ _17079_/Y _15222_/Y _18908_/S vssd1 vssd1 vccd1 vccd1 _18423_/X sky130_fd_sc_hd__mux2_1
X_15635_ _19704_/Q _15632_/X _15588_/X _15633_/X vssd1 vssd1 vccd1 vccd1 _19704_/D
+ sky130_fd_sc_hd__a22o_1
X_12847_ _12847_/A vssd1 vssd1 vccd1 vccd1 _12874_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__15965__B1 _15949_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13432__A input39/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12779__B1 _09630_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18354_ _18353_/X _21368_/Q _18850_/S vssd1 vssd1 vccd1 vccd1 _18354_/X sky130_fd_sc_hd__mux2_1
XANTENNA__19251__S0 _20132_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15566_ _19739_/Q _15561_/X _15550_/X _15563_/X vssd1 vssd1 vccd1 vccd1 _19739_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12778_ _12778_/A vssd1 vssd1 vccd1 vccd1 _12778_/X sky130_fd_sc_hd__buf_1
XPHY_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17305_ _19879_/Q vssd1 vssd1 vccd1 vccd1 _17305_/Y sky130_fd_sc_hd__inv_2
X_14517_ _14517_/A vssd1 vssd1 vccd1 vccd1 _14518_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_230_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11729_ _11737_/A vssd1 vssd1 vccd1 vccd1 _11729_/X sky130_fd_sc_hd__clkbuf_2
X_18285_ _18845_/A0 _10480_/Y _18896_/S vssd1 vssd1 vccd1 vccd1 _18285_/X sky130_fd_sc_hd__mux2_1
XFILLER_202_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18434__S _18680_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15497_ _19771_/Q _15492_/X _15456_/X _15494_/X vssd1 vssd1 vccd1 vccd1 _19771_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_174_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17236_ _19495_/Q vssd1 vssd1 vccd1 vccd1 _17236_/Y sky130_fd_sc_hd__inv_2
X_14448_ _20236_/Q _14446_/Y _14396_/Y _20219_/Q _14447_/X vssd1 vssd1 vccd1 vccd1
+ _14449_/D sky130_fd_sc_hd__o221a_1
XFILLER_80_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17167_ _17064_/A _17151_/X _17166_/Y _17154_/X vssd1 vssd1 vccd1 vccd1 _17167_/X
+ sky130_fd_sc_hd__o22a_1
X_14379_ _14379_/A vssd1 vssd1 vccd1 vccd1 _14380_/C sky130_fd_sc_hd__inv_2
XFILLER_115_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16118_ _19474_/Q _16108_/X _16117_/X _16111_/X vssd1 vssd1 vccd1 vccd1 _19474_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_127_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17098_ _19422_/Q vssd1 vssd1 vccd1 vccd1 _17098_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16049_ _16056_/A vssd1 vssd1 vccd1 vccd1 _16049_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__17890__B1 _18469_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11506__A1 _10892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12703__B1 _12544_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10714__C1 _10677_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19808_ _20172_/CLK _19808_/D vssd1 vssd1 vccd1 vccd1 _19808_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_226_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19739_ _19765_/CLK _19739_/D vssd1 vssd1 vccd1 vccd1 _19739_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__18609__S _18906_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09635__B1 _09633_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19242__S0 _19275_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_75_HCLK clkbuf_4_13_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20316_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_193_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18344__S _18907_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_134_HCLK_A clkbuf_4_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21354__RESET_B repeater252/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20514_ _20944_/CLK _20514_/D repeater275/X vssd1 vssd1 vccd1 vccd1 _20514_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_154_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20445_ _20480_/CLK _20445_/D repeater183/X vssd1 vssd1 vccd1 vccd1 _20445_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_134_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20376_ _20957_/CLK _20376_/D repeater185/X vssd1 vssd1 vccd1 vccd1 _20376_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_192_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17881__B1 _18474_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10060_ _21389_/Q vssd1 vssd1 vccd1 vccd1 _10150_/A sky130_fd_sc_hd__inv_2
XFILLER_102_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20236__RESET_B repeater204/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18519__S _18849_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15732__A input65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13750_ _20190_/Q vssd1 vssd1 vccd1 vccd1 _14579_/A sky130_fd_sc_hd__inv_2
X_10962_ _21199_/Q vssd1 vssd1 vccd1 vccd1 _10962_/Y sky130_fd_sc_hd__inv_2
XFILLER_244_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12701_ _12707_/A vssd1 vssd1 vccd1 vccd1 _12701_/X sky130_fd_sc_hd__buf_1
X_13681_ _20351_/Q _13679_/X _13482_/X _13680_/X vssd1 vssd1 vccd1 vccd1 _20351_/D
+ sky130_fd_sc_hd__a22o_1
X_10893_ _21254_/Q _10888_/X _10892_/X _10890_/X vssd1 vssd1 vccd1 vccd1 _21254_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_204_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_14_0_HCLK clkbuf_3_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_14_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_15420_ _19803_/Q _15415_/X _15386_/X _15417_/X vssd1 vssd1 vccd1 vccd1 _19803_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12632_ _12638_/A vssd1 vssd1 vccd1 vccd1 _12632_/X sky130_fd_sc_hd__buf_1
XPHY_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19233__S0 _19275_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12563_ _19983_/Q _12561_/B input37/X _11795_/A vssd1 vssd1 vccd1 vccd1 _16527_/B
+ sky130_fd_sc_hd__o211a_1
X_15351_ _19832_/Q _15345_/X _15350_/X _15347_/X vssd1 vssd1 vccd1 vccd1 _19832_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18254__S _18891_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21095__RESET_B repeater226/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11514_ _21146_/Q vssd1 vssd1 vccd1 vccd1 _11514_/Y sky130_fd_sc_hd__inv_2
X_14302_ _14302_/A _14302_/B _14302_/C _14324_/A vssd1 vssd1 vccd1 vccd1 _14302_/X
+ sky130_fd_sc_hd__or4b_1
XPHY_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18070_ _20839_/Q vssd1 vssd1 vccd1 vccd1 _18070_/Y sky130_fd_sc_hd__inv_2
XFILLER_200_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15282_ _20489_/Q _15104_/X _20467_/Q _15061_/A vssd1 vssd1 vccd1 vccd1 _15282_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_11_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12494_ _12396_/B _12493_/A _20920_/Q _12496_/A _12438_/X vssd1 vssd1 vccd1 vccd1
+ _20920_/D sky130_fd_sc_hd__o221a_1
XPHY_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17021_ _17021_/A _17023_/B vssd1 vssd1 vccd1 vccd1 _20007_/D sky130_fd_sc_hd__nor2_1
X_11445_ _21157_/Q _11445_/B vssd1 vssd1 vccd1 vccd1 _11446_/B sky130_fd_sc_hd__or2_1
X_14233_ _19893_/Q _14233_/B vssd1 vssd1 vccd1 vccd1 _14234_/B sky130_fd_sc_hd__or2_1
XFILLER_109_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_56_HCLK_A clkbuf_4_12_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12933__B1 _12932_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14164_ _20546_/Q vssd1 vssd1 vccd1 vccd1 _14164_/Y sky130_fd_sc_hd__inv_2
X_11376_ _11410_/A _16595_/B _11376_/C _11376_/D vssd1 vssd1 vccd1 vccd1 _11376_/X
+ sky130_fd_sc_hd__and4bb_1
XFILLER_180_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13115_ _13133_/A vssd1 vssd1 vccd1 vccd1 _13115_/X sky130_fd_sc_hd__buf_1
X_10327_ _10274_/A _20718_/Q _21359_/Q _10326_/Y vssd1 vssd1 vccd1 vccd1 _10327_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__17872__B1 _18581_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14095_ _14095_/A _14095_/B vssd1 vssd1 vccd1 vccd1 _14182_/A sky130_fd_sc_hd__or2_1
X_18972_ _16525_/X _16515_/Y _18975_/S vssd1 vssd1 vccd1 vccd1 _18972_/X sky130_fd_sc_hd__mux2_1
XFILLER_140_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17923_ _17315_/X _17853_/A _18928_/S _17852_/A _17830_/X vssd1 vssd1 vccd1 vccd1
+ _18018_/A sky130_fd_sc_hd__a2111oi_2
X_13046_ _13046_/A vssd1 vssd1 vccd1 vccd1 _13657_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_59_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10258_ _21345_/Q vssd1 vssd1 vccd1 vccd1 _10261_/A sky130_fd_sc_hd__inv_2
XFILLER_39_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17854_ _17854_/A vssd1 vssd1 vccd1 vccd1 _17854_/X sky130_fd_sc_hd__buf_1
XFILLER_79_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10189_ _10155_/A _10155_/B _10185_/X _10187_/Y vssd1 vssd1 vccd1 vccd1 _21394_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_94_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16805_ _19932_/Q vssd1 vssd1 vccd1 vccd1 _16805_/Y sky130_fd_sc_hd__inv_2
XFILLER_208_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17785_ _21051_/Q vssd1 vssd1 vccd1 vccd1 _17785_/Y sky130_fd_sc_hd__inv_2
X_14997_ _14997_/A vssd1 vssd1 vccd1 vccd1 _15019_/A sky130_fd_sc_hd__buf_1
XANTENNA__18429__S _18884_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16738__A _21144_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19524_ _20327_/CLK _19524_/D vssd1 vssd1 vccd1 vccd1 _19524_/Q sky130_fd_sc_hd__dfxtp_1
X_16736_ _20998_/Q _12003_/X _20998_/Q _12003_/X vssd1 vssd1 vccd1 vccd1 _16736_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_81_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13948_ _20646_/Q vssd1 vssd1 vccd1 vccd1 _13948_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_1_1_0_HCLK clkbuf_0_HCLK/X vssd1 vssd1 vccd1 vccd1 clkbuf_1_1_1_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_223_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_98_HCLK clkbuf_4_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20661_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__09640__A input44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19455_ _21234_/CLK _19455_/D vssd1 vssd1 vccd1 vccd1 _19455_/Q sky130_fd_sc_hd__dfxtp_1
X_16667_ _21155_/Q _11443_/B _11444_/B vssd1 vssd1 vccd1 vccd1 _16667_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__15938__B1 _15887_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14258__A _14258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13879_ _13972_/C _13879_/B vssd1 vssd1 vccd1 vccd1 _14006_/A sky130_fd_sc_hd__or2_1
XFILLER_234_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18406_ _17079_/Y _15238_/Y _18908_/S vssd1 vssd1 vccd1 vccd1 _18406_/X sky130_fd_sc_hd__mux2_1
XFILLER_222_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15618_ _15618_/A vssd1 vssd1 vccd1 vccd1 _15618_/X sky130_fd_sc_hd__buf_1
XANTENNA__19224__S0 _19275_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19386_ _20331_/CLK _19386_/D vssd1 vssd1 vccd1 vccd1 _19386_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16598_ _21418_/Q vssd1 vssd1 vccd1 vccd1 _16598_/Y sky130_fd_sc_hd__inv_2
X_18337_ _18336_/X _10614_/Y _18897_/S vssd1 vssd1 vccd1 vccd1 _18337_/X sky130_fd_sc_hd__mux2_1
X_15549_ _19748_/Q _15543_/X _15548_/X _15546_/X vssd1 vssd1 vccd1 vccd1 _19748_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16473__A _16473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18164__S _18903_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18268_ _18006_/Y _20795_/Q _18885_/S vssd1 vssd1 vccd1 vccd1 _18268_/X sky130_fd_sc_hd__mux2_1
XFILLER_136_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_4_HCLK clkbuf_opt_2_HCLK/A vssd1 vssd1 vccd1 vccd1 _19813_/CLK sky130_fd_sc_hd__clkbuf_16
X_17219_ _17857_/A vssd1 vssd1 vccd1 vccd1 _17219_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_190_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19842__RESET_B repeater212/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18199_ _18198_/X _16821_/Y _18667_/S vssd1 vssd1 vccd1 vccd1 _18199_/X sky130_fd_sc_hd__mux2_1
X_20230_ _21485_/CLK _20230_/D repeater203/X vssd1 vssd1 vccd1 vccd1 _20230_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_144_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20161_ _21121_/CLK _20161_/D repeater237/X vssd1 vssd1 vccd1 vccd1 _20161_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17863__B1 _18562_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09972_ _21420_/Q _09968_/X _09666_/X _09970_/X vssd1 vssd1 vccd1 vccd1 _21420_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_143_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20092_ _20496_/CLK _20092_/D repeater273/X vssd1 vssd1 vccd1 vccd1 _20092_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__12152__A1 _12036_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18339__S _18680_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13101__B1 _12879_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_226_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20994_ _21338_/CLK _20994_/D repeater222/X vssd1 vssd1 vccd1 vccd1 _20994_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_26_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17918__B2 _17203_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_241_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15929__B1 _15788_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_241_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13072__A _13072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19215__S0 _19275_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_213_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19135__A3 _19815_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13168__B1 _13166_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21477_ _21477_/CLK _21477_/D repeater201/X vssd1 vssd1 vccd1 vccd1 _21477_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__18802__S _18875_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11230_ _21197_/Q _11225_/X _10900_/X _11226_/X vssd1 vssd1 vccd1 vccd1 _21197_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16106__B1 _15916_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20428_ _20428_/CLK _20428_/D repeater269/X vssd1 vssd1 vccd1 vccd1 _20428_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_20_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11161_ _13182_/A _20597_/Q _16525_/C vssd1 vssd1 vccd1 vccd1 _16524_/A sky130_fd_sc_hd__or3_4
XFILLER_136_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20359_ _20982_/CLK _20359_/D repeater279/X vssd1 vssd1 vccd1 vccd1 _20359_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_161_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20417__RESET_B repeater187/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10112_ _10102_/X _10112_/B _10112_/C _10112_/D vssd1 vssd1 vccd1 vccd1 _10137_/B
+ sky130_fd_sc_hd__and4b_1
X_11092_ _11092_/A vssd1 vssd1 vccd1 vccd1 _21233_/D sky130_fd_sc_hd__inv_2
XFILLER_49_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14920_ _20569_/Q _15000_/A _20582_/Q _14961_/B vssd1 vssd1 vccd1 vccd1 _14920_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_76_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10043_ _21382_/Q vssd1 vssd1 vccd1 vccd1 _10203_/A sky130_fd_sc_hd__inv_2
XFILLER_49_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20070__RESET_B repeater276/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input25_A HADDR[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14851_ _20078_/Q vssd1 vssd1 vccd1 vccd1 _14853_/B sky130_fd_sc_hd__inv_2
XFILLER_64_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13802_ _20610_/Q vssd1 vssd1 vccd1 vccd1 _13802_/Y sky130_fd_sc_hd__inv_2
XFILLER_91_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17570_ _18021_/A vssd1 vssd1 vccd1 vccd1 _17955_/A sky130_fd_sc_hd__inv_2
X_14782_ _19126_/X vssd1 vssd1 vccd1 vccd1 _14783_/A sky130_fd_sc_hd__inv_2
XFILLER_63_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11994_ _20988_/Q _11994_/B vssd1 vssd1 vccd1 vccd1 _11995_/B sky130_fd_sc_hd__or2_1
XFILLER_29_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16521_ _16576_/B _16521_/B vssd1 vssd1 vccd1 vccd1 _16686_/A sky130_fd_sc_hd__or2_2
XFILLER_44_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13733_ _20324_/Q vssd1 vssd1 vccd1 vccd1 _16127_/A sky130_fd_sc_hd__buf_1
XFILLER_90_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10945_ _21025_/Q vssd1 vssd1 vccd1 vccd1 _11863_/A sky130_fd_sc_hd__inv_2
XFILLER_216_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__21276__RESET_B repeater245/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19240_ _17440_/Y _17441_/Y _17442_/Y _17443_/Y _20130_/Q _20131_/Q vssd1 vssd1 vccd1
+ vccd1 _19240_/X sky130_fd_sc_hd__mux4_2
XFILLER_45_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16452_ _16459_/A vssd1 vssd1 vccd1 vccd1 _16452_/X sky130_fd_sc_hd__buf_1
XFILLER_231_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13664_ _20362_/Q _13659_/X _13543_/X _13662_/X vssd1 vssd1 vccd1 vccd1 _20362_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19206__S0 _21005_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10876_ _21260_/Q _10871_/X _09702_/X _10872_/X vssd1 vssd1 vccd1 vccd1 _21260_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_188_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15403_ _19811_/Q _15398_/X _15386_/X _15400_/X vssd1 vssd1 vccd1 vccd1 _19811_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_231_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19171_ _19167_/X _19168_/X _19169_/X _19170_/X _20123_/Q _20124_/Q vssd1 vssd1 vccd1
+ vccd1 _19171_/X sky130_fd_sc_hd__mux4_2
X_12615_ input13/X _12613_/X _20863_/Q _12614_/X vssd1 vssd1 vccd1 vccd1 _20863_/D
+ sky130_fd_sc_hd__o22a_1
XPHY_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16383_ _19346_/Q _16378_/X _16202_/X _16380_/X vssd1 vssd1 vccd1 vccd1 _19346_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_197_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_repeater164_A _18835_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13595_ _13595_/A vssd1 vssd1 vccd1 vccd1 _13595_/X sky130_fd_sc_hd__buf_1
XPHY_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18122_ vssd1 vssd1 vccd1 vccd1 _18122_/HI _18122_/LO sky130_fd_sc_hd__conb_1
XANTENNA__13710__A _13710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15334_ _15574_/C vssd1 vssd1 vccd1 vccd1 _16481_/A sky130_fd_sc_hd__buf_1
X_12546_ _12554_/A vssd1 vssd1 vccd1 vccd1 _12546_/X sky130_fd_sc_hd__buf_1
XFILLER_8_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18053_ _20837_/Q vssd1 vssd1 vccd1 vccd1 _18053_/Y sky130_fd_sc_hd__inv_2
XFILLER_177_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15265_ _20491_/Q vssd1 vssd1 vccd1 vccd1 _15265_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18712__S _18880_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12477_ _20929_/Q _12476_/Y _12480_/A _12419_/B vssd1 vssd1 vccd1 vccd1 _20929_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_138_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17004_ _17004_/A vssd1 vssd1 vccd1 vccd1 _17004_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12906__B1 _12656_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output93_A _18014_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14216_ _14216_/A vssd1 vssd1 vccd1 vccd1 _14216_/Y sky130_fd_sc_hd__inv_2
X_11428_ _11387_/A _11420_/X _11389_/B _11421_/X vssd1 vssd1 vccd1 vccd1 _21175_/D
+ sky130_fd_sc_hd__o22a_1
X_15196_ _20057_/Q _15195_/Y _15185_/X _15072_/B vssd1 vssd1 vccd1 vccd1 _20057_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_153_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20840__RESET_B repeater251/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17845__B1 _18612_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11359_ _11359_/A vssd1 vssd1 vccd1 vccd1 _11411_/A sky130_fd_sc_hd__inv_2
XFILLER_140_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14147_ _20555_/Q vssd1 vssd1 vccd1 vccd1 _14147_/Y sky130_fd_sc_hd__inv_2
XFILLER_193_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18955_ _16649_/X _21081_/Q _18962_/S vssd1 vssd1 vccd1 vccd1 _18955_/X sky130_fd_sc_hd__mux2_1
X_14078_ _14078_/A _14078_/B vssd1 vssd1 vccd1 vccd1 _14216_/A sky130_fd_sc_hd__or2_2
X_13029_ _20676_/Q _13026_/X _12863_/X _13027_/X vssd1 vssd1 vccd1 vccd1 _20676_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17906_ _18445_/X _17200_/X _18434_/X _17224_/X _17905_/Y vssd1 vssd1 vccd1 vccd1
+ _17906_/X sky130_fd_sc_hd__o221a_1
XFILLER_67_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18886_ _18885_/X _10260_/A _18886_/S vssd1 vssd1 vccd1 vccd1 _18886_/X sky130_fd_sc_hd__mux2_1
X_17837_ _17835_/Y _17472_/A _17836_/Y _17474_/A vssd1 vssd1 vccd1 vccd1 _17838_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_239_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18159__S _18666_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12996__A input57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16468__A _16474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_242_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17768_ _19356_/Q vssd1 vssd1 vccd1 vccd1 _17768_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16719_ _19903_/Q _14243_/B _18946_/S vssd1 vssd1 vccd1 vccd1 _16719_/X sky130_fd_sc_hd__a21o_1
X_19507_ _20327_/CLK _19507_/D vssd1 vssd1 vccd1 vccd1 _19507_/Q sky130_fd_sc_hd__dfxtp_1
X_17699_ _19444_/Q vssd1 vssd1 vccd1 vccd1 _17699_/Y sky130_fd_sc_hd__inv_2
XFILLER_212_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19438_ _20137_/CLK _19438_/D vssd1 vssd1 vccd1 vccd1 _19438_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19369_ _19828_/CLK _19369_/D vssd1 vssd1 vccd1 vccd1 _19369_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21400_ _21405_/CLK _21400_/D repeater253/X vssd1 vssd1 vccd1 vccd1 _21400_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__13620__A _13626_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11948__B2 _11932_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21331_ _21476_/CLK _21331_/D repeater204/X vssd1 vssd1 vccd1 vccd1 _21331_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_191_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10620__B2 _20767_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18622__S _18898_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_21262_ _21433_/CLK _21262_/D repeater234/X vssd1 vssd1 vccd1 vccd1 _21262_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_144_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_105_HCLK clkbuf_4_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20946_/CLK sky130_fd_sc_hd__clkbuf_16
X_20213_ _20220_/CLK _20213_/D repeater203/X vssd1 vssd1 vccd1 vccd1 _20213_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_104_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21193_ _21193_/CLK _21193_/D repeater224/X vssd1 vssd1 vccd1 vccd1 _21193_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_143_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20510__RESET_B repeater267/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20144_ _21239_/CLK _20144_/D repeater250/X vssd1 vssd1 vccd1 vccd1 _20144_/Q sky130_fd_sc_hd__dfrtp_1
X_09955_ _21427_/Q _09950_/X _09682_/X _09952_/X vssd1 vssd1 vccd1 vccd1 _21427_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_131_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13067__A _13073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20075_ _20075_/CLK _20075_/D repeater276/X vssd1 vssd1 vccd1 vccd1 _20075_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_131_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09886_ _09886_/A vssd1 vssd1 vccd1 vccd1 _09887_/B sky130_fd_sc_hd__inv_2
XFILLER_106_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18013__B1 _18162_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20977_ _20982_/CLK _20977_/D repeater278/X vssd1 vssd1 vccd1 vccd1 _20977_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_4569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10730_ _10723_/A _10723_/B _21310_/Q _10647_/A _10670_/X vssd1 vssd1 vccd1 vccd1
+ _21310_/D sky130_fd_sc_hd__o221a_1
XFILLER_241_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10661_ _10661_/A _10661_/B vssd1 vssd1 vccd1 vccd1 _10679_/A sky130_fd_sc_hd__or2_1
XFILLER_9_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12400_ _20932_/Q vssd1 vssd1 vccd1 vccd1 _12421_/A sky130_fd_sc_hd__inv_2
XFILLER_167_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13380_ _20500_/Q _13377_/X _13169_/X _13378_/X vssd1 vssd1 vccd1 vccd1 _20500_/D
+ sky130_fd_sc_hd__a22o_1
X_10592_ _20751_/Q vssd1 vssd1 vccd1 vccd1 _10592_/Y sky130_fd_sc_hd__inv_2
XFILLER_222_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20669__RESET_B repeater207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12331_ _12331_/A _12331_/B vssd1 vssd1 vccd1 vccd1 _12339_/A sky130_fd_sc_hd__or2_1
XANTENNA__18532__S _18875_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15050_ _20052_/Q vssd1 vssd1 vccd1 vccd1 _15093_/A sky130_fd_sc_hd__inv_2
X_12262_ _12472_/A _20504_/Q _12427_/A _20518_/Q _12261_/X vssd1 vssd1 vccd1 vccd1
+ _12262_/X sky130_fd_sc_hd__a221o_1
XFILLER_141_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14001_ _13883_/A _13883_/B _13999_/Y _13991_/X vssd1 vssd1 vccd1 vccd1 _20307_/D
+ sky130_fd_sc_hd__a211oi_2
X_11213_ _11225_/A vssd1 vssd1 vccd1 vccd1 _11213_/X sky130_fd_sc_hd__buf_1
X_12193_ _20976_/Q _12191_/Y _12314_/A _20343_/Q _12192_/X vssd1 vssd1 vccd1 vccd1
+ _12193_/X sky130_fd_sc_hd__a221o_1
X_11144_ _11141_/X _11143_/Y _11141_/X _11143_/Y vssd1 vssd1 vccd1 vccd1 _11151_/C
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_68_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput85 _17919_/Y vssd1 vssd1 vccd1 vccd1 HRDATA[15] sky130_fd_sc_hd__clkbuf_2
XFILLER_122_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput96 _18051_/Y vssd1 vssd1 vccd1 vccd1 HRDATA[25] sky130_fd_sc_hd__clkbuf_2
X_18740_ _17608_/X _19587_/Q _18926_/S vssd1 vssd1 vccd1 vccd1 _18740_/X sky130_fd_sc_hd__mux2_1
X_15952_ _19558_/Q _15943_/X _15951_/X _15945_/X vssd1 vssd1 vccd1 vccd1 _19558_/D
+ sky130_fd_sc_hd__a22o_1
X_11075_ _21236_/Q _11075_/B vssd1 vssd1 vccd1 vccd1 _11075_/Y sky130_fd_sc_hd__nor2_1
XFILLER_237_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14903_ _20574_/Q vssd1 vssd1 vccd1 vccd1 _14903_/Y sky130_fd_sc_hd__inv_2
X_10026_ _10908_/A _10026_/B _17060_/C vssd1 vssd1 vccd1 vccd1 _10028_/S sky130_fd_sc_hd__or3_4
X_18671_ _17777_/Y _09996_/Y _20870_/Q vssd1 vssd1 vccd1 vccd1 _18671_/X sky130_fd_sc_hd__mux2_1
XANTENNA_output131_A _20004_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15883_ _19590_/Q _15875_/X _15812_/X _15877_/X vssd1 vssd1 vccd1 vccd1 _19590_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_49_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__21457__RESET_B repeater245/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17622_ _19354_/Q vssd1 vssd1 vccd1 vccd1 _17622_/Y sky130_fd_sc_hd__inv_2
X_14834_ _20098_/Q vssd1 vssd1 vccd1 vccd1 _14835_/A sky130_fd_sc_hd__inv_2
XFILLER_63_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17553_ _17553_/A vssd1 vssd1 vccd1 vccd1 _17553_/X sky130_fd_sc_hd__buf_1
X_14765_ _20132_/Q _14758_/B _14753_/B vssd1 vssd1 vccd1 vccd1 _14765_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_17_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18707__S _18928_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11977_ _21000_/Q vssd1 vssd1 vccd1 vccd1 _11978_/A sky130_fd_sc_hd__inv_2
X_16504_ _21093_/Q _16499_/X _16501_/X _16503_/Y vssd1 vssd1 vccd1 vccd1 _16505_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_60_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15920__A _15927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13716_ _20331_/Q vssd1 vssd1 vccd1 vccd1 _15758_/A sky130_fd_sc_hd__buf_1
X_10928_ _21211_/Q vssd1 vssd1 vccd1 vccd1 _10928_/Y sky130_fd_sc_hd__inv_2
X_17484_ _19498_/Q vssd1 vssd1 vccd1 vccd1 _17484_/Y sky130_fd_sc_hd__inv_2
X_14696_ _14696_/A vssd1 vssd1 vccd1 vccd1 _14696_/X sky130_fd_sc_hd__buf_1
X_19223_ _17592_/Y _17593_/Y _17594_/Y _17595_/Y _19275_/S0 _21004_/Q vssd1 vssd1
+ vccd1 vccd1 _19223_/X sky130_fd_sc_hd__mux4_2
XFILLER_177_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16435_ _16441_/A vssd1 vssd1 vccd1 vccd1 _16442_/A sky130_fd_sc_hd__inv_2
X_13647_ _20371_/Q _13645_/X _13506_/X _13646_/X vssd1 vssd1 vccd1 vccd1 _20371_/D
+ sky130_fd_sc_hd__a22o_1
X_10859_ _13188_/A _10859_/B _13327_/C vssd1 vssd1 vccd1 vccd1 _17195_/A sky130_fd_sc_hd__or3_4
XFILLER_158_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19154_ _19691_/Q _19379_/Q _19675_/Q _19667_/Q _19285_/S0 _21017_/Q vssd1 vssd1
+ vccd1 vccd1 _19154_/X sky130_fd_sc_hd__mux4_2
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16366_ _19356_/Q _16363_/X _16196_/X _16365_/X vssd1 vssd1 vccd1 vccd1 _19356_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_13_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16318__B1 _16006_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13578_ _20410_/Q _13573_/X _13424_/X _13575_/X vssd1 vssd1 vccd1 vccd1 _20410_/D
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_128_HCLK clkbuf_4_4_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20809_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_157_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18105_ _17925_/A _18105_/B _18105_/C vssd1 vssd1 vccd1 vccd1 _18105_/Y sky130_fd_sc_hd__nand3b_4
XFILLER_173_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15317_ _18281_/S _09870_/A _09852_/Y _15315_/Y _15316_/X vssd1 vssd1 vccd1 vccd1
+ _15318_/A sky130_fd_sc_hd__o311a_1
XFILLER_8_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12529_ _11541_/B _12527_/X _11272_/A _12528_/X vssd1 vssd1 vccd1 vccd1 _20913_/D
+ sky130_fd_sc_hd__o22ai_1
X_19085_ _21048_/Q _21061_/Q _19872_/Q vssd1 vssd1 vccd1 vccd1 _19085_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18442__S _18908_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16297_ _16297_/A _21221_/Q _16297_/C vssd1 vssd1 vccd1 vccd1 _16305_/A sky130_fd_sc_hd__or3_4
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18036_ _20835_/Q _18084_/B vssd1 vssd1 vccd1 vccd1 _18036_/Y sky130_fd_sc_hd__nand2_1
XFILLER_117_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15248_ _20490_/Q _15083_/A _20484_/Q _15077_/A vssd1 vssd1 vccd1 vccd1 _15248_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_172_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21130__CLK _21134_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13552__B1 _13550_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15179_ _15179_/A vssd1 vssd1 vccd1 vccd1 _15179_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_59_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19987_ _21196_/CLK _19987_/D repeater218/X vssd1 vssd1 vccd1 vccd1 _19987_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_86_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13304__B1 _13144_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09740_ _20146_/Q vssd1 vssd1 vccd1 vccd1 _09740_/Y sky130_fd_sc_hd__inv_2
X_18938_ _16708_/X _21138_/Q _18946_/S vssd1 vssd1 vccd1 vccd1 _18938_/X sky130_fd_sc_hd__mux2_1
.ends

