magic
tech sky130A
magscale 1 2
timestamp 1621801760
<< nwell >>
rect 1066 277157 218906 277478
rect 1066 276069 218906 276635
rect 1066 274981 218906 275547
rect 1066 273903 218906 274459
rect 1066 273893 90911 273903
rect 1066 273361 65532 273371
rect 1066 272815 218906 273361
rect 1066 272805 22936 272815
rect 1066 272273 54939 272283
rect 1066 271727 218906 272273
rect 1066 271717 25407 271727
rect 1066 271185 21267 271195
rect 1066 270639 218906 271185
rect 1066 270629 35251 270639
rect 1066 270097 8492 270107
rect 1066 269551 218906 270097
rect 1066 269541 7296 269551
rect 1066 269009 17219 269019
rect 1066 268463 218906 269009
rect 1066 268453 4352 268463
rect 1066 267921 4904 267931
rect 1066 267375 218906 267921
rect 1066 267365 5180 267375
rect 1066 266833 23107 266843
rect 1066 266287 218906 266833
rect 1066 266277 17955 266287
rect 1066 265745 56871 265755
rect 1066 265199 218906 265745
rect 1066 265189 13815 265199
rect 1066 264657 44543 264667
rect 1066 264111 218906 264657
rect 1066 264101 35816 264111
rect 1066 263569 48223 263579
rect 1066 263023 218906 263569
rect 1066 263013 4720 263023
rect 1066 262481 16943 262491
rect 1066 261935 218906 262481
rect 1066 261925 8111 261935
rect 1066 261393 11988 261403
rect 1066 260847 218906 261393
rect 1066 260837 8308 260847
rect 1066 260305 4996 260315
rect 1066 259759 218906 260305
rect 1066 259749 47211 259759
rect 1066 259217 36815 259227
rect 1066 258671 218906 259217
rect 1066 258661 47211 258671
rect 1066 258129 5088 258139
rect 1066 257583 218906 258129
rect 1066 257573 14472 257583
rect 1066 257041 4983 257051
rect 1066 256495 218906 257041
rect 1066 256485 37104 256495
rect 1066 255953 41336 255963
rect 1066 255407 218906 255953
rect 1066 255397 25683 255407
rect 1066 254865 36999 254875
rect 1066 254319 218906 254865
rect 1066 254309 9964 254319
rect 1066 253777 17035 253787
rect 1066 253231 218906 253777
rect 1066 253221 5456 253231
rect 1066 252689 36092 252699
rect 1066 252143 218906 252689
rect 1066 252133 22831 252143
rect 1066 251601 68831 251611
rect 1066 251055 218906 251601
rect 1066 251045 19887 251055
rect 1066 250513 53559 250523
rect 1066 249967 218906 250513
rect 1066 249957 4523 249967
rect 1066 249425 4904 249435
rect 1066 248879 218906 249425
rect 1066 248869 9031 248879
rect 1066 248337 26143 248347
rect 1066 247791 218906 248337
rect 1066 247781 9964 247791
rect 1066 247249 12803 247259
rect 1066 246703 218906 247249
rect 1066 246693 22371 246703
rect 1066 246161 7099 246171
rect 1066 245615 218906 246161
rect 1066 245605 17127 245615
rect 1066 245073 4628 245083
rect 1066 244527 218906 245073
rect 1066 244517 48683 244527
rect 1066 243985 36092 243995
rect 1066 243439 218906 243985
rect 1066 243429 4260 243439
rect 1066 242897 44924 242907
rect 1066 242351 218906 242897
rect 1066 242341 17127 242351
rect 1066 241809 6468 241819
rect 1066 241263 218906 241809
rect 1066 241253 12448 241263
rect 1066 240721 23672 240731
rect 1066 240175 218906 240721
rect 1066 240165 23107 240175
rect 1066 239633 4904 239643
rect 1066 239087 218906 239633
rect 1066 239077 9044 239087
rect 1066 238545 23291 238555
rect 1066 237999 218906 238545
rect 1066 237989 21188 237999
rect 1066 237457 9307 237467
rect 1066 236911 218906 237457
rect 1066 236901 169571 236911
rect 1066 236369 5732 236379
rect 1066 235823 218906 236369
rect 1066 235813 177312 235823
rect 1066 235281 23199 235291
rect 1066 234735 218906 235281
rect 1066 234725 9675 234735
rect 1066 234193 20347 234203
rect 1066 233647 218906 234193
rect 1066 233637 5088 233647
rect 1066 233105 44543 233115
rect 1066 232559 218906 233105
rect 1066 232549 15747 232559
rect 1066 232017 194976 232027
rect 1066 231471 218906 232017
rect 1066 231461 4983 231471
rect 1066 230929 4615 230939
rect 1066 230383 218906 230929
rect 1066 230373 4352 230383
rect 1066 229841 21727 229851
rect 1066 229295 218906 229841
rect 1066 229285 5180 229295
rect 1066 228753 16483 228763
rect 1066 228207 218906 228753
rect 1066 228197 4352 228207
rect 1066 227665 25039 227675
rect 1066 227119 218906 227665
rect 1066 227109 12448 227119
rect 1066 226577 41047 226587
rect 1066 226031 218906 226577
rect 1066 226021 85299 226031
rect 1066 225489 71144 225499
rect 1066 224943 218906 225489
rect 1066 224933 28443 224943
rect 1066 224401 12816 224411
rect 1066 223855 218906 224401
rect 1066 223845 81711 223855
rect 1066 223313 9872 223323
rect 1066 222767 218906 223313
rect 1066 222757 10516 222767
rect 1066 222225 124675 222235
rect 1066 221679 218906 222225
rect 1066 221669 37288 221679
rect 1066 221137 122927 221147
rect 1066 220591 218906 221137
rect 1066 220581 47027 220591
rect 1066 220049 42979 220059
rect 1066 219503 218906 220049
rect 1066 219493 36723 219503
rect 1066 218961 70868 218971
rect 1066 218415 218906 218961
rect 1066 218405 41244 218415
rect 1066 217873 69488 217883
rect 1066 217327 218906 217873
rect 1066 217317 35251 217327
rect 1066 216785 44372 216795
rect 1066 216239 218906 216785
rect 1066 216229 35724 216239
rect 1066 215697 104435 215707
rect 1066 215151 218906 215697
rect 1066 215141 102884 215151
rect 1066 214609 191467 214619
rect 1066 214063 218906 214609
rect 1066 214053 18507 214063
rect 1066 213521 25039 213531
rect 1066 212975 218906 213521
rect 1066 212965 10976 212975
rect 1066 212433 4628 212443
rect 1066 211887 218906 212433
rect 1066 211877 5259 211887
rect 1066 211345 83643 211355
rect 1066 210799 218906 211345
rect 1066 210789 72695 210799
rect 1066 210257 66176 210267
rect 1066 209711 218906 210257
rect 1066 209701 4352 209711
rect 1066 209169 97088 209179
rect 1066 208623 218906 209169
rect 1066 208613 4983 208623
rect 1066 208081 9872 208091
rect 1066 207535 218906 208081
rect 1066 207525 13999 207535
rect 1066 206993 14551 207003
rect 1066 206447 218906 206993
rect 1066 206437 5548 206447
rect 1066 205905 53467 205915
rect 1066 205359 218906 205905
rect 1066 205349 65979 205359
rect 1066 204817 49984 204827
rect 1066 204271 218906 204817
rect 1066 204261 13631 204271
rect 1066 203729 5364 203739
rect 1066 203183 218906 203729
rect 1066 203173 5075 203183
rect 1066 202641 9399 202651
rect 1066 202095 218906 202641
rect 1066 202085 76191 202095
rect 1066 201553 137384 201563
rect 1066 201007 218906 201553
rect 1066 200997 37288 201007
rect 1066 200465 32583 200475
rect 1066 199919 218906 200465
rect 1066 199909 65979 199919
rect 1066 199377 39391 199387
rect 1066 198831 218906 199377
rect 1066 198821 70224 198831
rect 1066 198289 22463 198299
rect 1066 197743 218906 198289
rect 1066 197733 10608 197743
rect 1066 197201 11712 197211
rect 1066 196655 218906 197201
rect 1066 196645 5548 196655
rect 1066 196113 4720 196123
rect 1066 195567 218906 196113
rect 1066 195557 5732 195567
rect 1066 195025 196711 195035
rect 1066 194479 218906 195025
rect 1066 194469 14275 194479
rect 1066 193937 5719 193947
rect 1066 193391 218906 193937
rect 1066 193381 40508 193391
rect 1066 192849 21635 192859
rect 1066 192303 218906 192849
rect 1066 192293 4352 192303
rect 1066 191761 4628 191771
rect 1066 191215 218906 191761
rect 1066 191205 66820 191215
rect 1066 190673 37091 190683
rect 1066 190127 218906 190673
rect 1066 190117 14183 190127
rect 1066 189585 5088 189595
rect 1066 189039 218906 189585
rect 1066 189029 40968 189039
rect 1066 188497 10516 188507
rect 1066 187951 218906 188497
rect 1066 187941 5548 187951
rect 1066 187409 32412 187419
rect 1066 186863 218906 187409
rect 1066 186853 50812 186863
rect 1066 186321 9872 186331
rect 1066 185775 218906 186321
rect 1066 185765 12159 185775
rect 1066 185233 21359 185243
rect 1066 184687 218906 185233
rect 1066 184677 83827 184687
rect 1066 184145 11883 184155
rect 1066 183599 218906 184145
rect 1066 183589 5272 183599
rect 1066 183057 4628 183067
rect 1066 182511 218906 183057
rect 1066 182501 49971 182511
rect 1066 181969 18415 181979
rect 1066 181423 218906 181969
rect 1066 181413 37288 181423
rect 1066 180881 33595 180891
rect 1066 180335 218906 180881
rect 1066 180325 4536 180335
rect 1066 179793 12803 179803
rect 1066 179247 218906 179793
rect 1066 179237 25499 179247
rect 1066 178705 69396 178715
rect 1066 178159 218906 178705
rect 1066 178149 43531 178159
rect 1066 177617 69015 177627
rect 1066 177071 218906 177617
rect 1066 177061 5640 177071
rect 1066 176529 15747 176539
rect 1066 175983 218906 176529
rect 1066 175973 5732 175983
rect 1066 175441 5995 175451
rect 1066 174895 218906 175441
rect 1066 174885 22936 174895
rect 1066 174353 37275 174363
rect 1066 173807 218906 174353
rect 1066 173797 4983 173807
rect 1066 173265 53467 173275
rect 1066 172719 218906 173265
rect 1066 172709 43807 172719
rect 1066 172177 32215 172187
rect 1066 171631 218906 172177
rect 1066 171621 117315 171631
rect 1066 171089 46751 171099
rect 1066 170543 218906 171089
rect 1066 170533 33424 170543
rect 1066 170001 34712 170011
rect 1066 169455 218906 170001
rect 1066 169445 96536 169455
rect 1066 168913 4904 168923
rect 1066 168367 218906 168913
rect 1066 168357 10608 168367
rect 1066 167825 5075 167835
rect 1066 167279 218906 167825
rect 1066 167269 5732 167279
rect 1066 166737 53007 166747
rect 1066 166191 218906 166737
rect 1066 166181 14275 166191
rect 1066 165649 130484 165659
rect 1066 165103 218906 165649
rect 1066 165093 96628 165103
rect 1066 164561 32872 164571
rect 1066 164015 218906 164561
rect 1066 164005 14367 164015
rect 1066 163473 6560 163483
rect 1066 162927 218906 163473
rect 1066 162917 47684 162927
rect 1066 162385 20991 162395
rect 1066 161839 218906 162385
rect 1066 161829 17403 161839
rect 1066 161297 6100 161307
rect 1066 160751 218906 161297
rect 1066 160741 9780 160751
rect 1066 160209 5811 160219
rect 1066 159663 218906 160209
rect 1066 159653 4155 159663
rect 1066 159121 17679 159131
rect 1066 158575 218906 159121
rect 1066 158565 33227 158575
rect 1066 158033 4628 158043
rect 1066 157487 218906 158033
rect 1066 157477 36447 157487
rect 1066 156945 69751 156955
rect 1066 156399 218906 156945
rect 1066 156389 43623 156399
rect 1066 155857 36460 155867
rect 1066 155311 218906 155857
rect 1066 155301 40219 155311
rect 1066 154769 67556 154779
rect 1066 154223 218906 154769
rect 1066 154213 70119 154223
rect 1066 153681 37735 153691
rect 1066 153135 218906 153681
rect 1066 153125 90543 153135
rect 1066 152593 161383 152603
rect 1066 152047 218906 152593
rect 1066 152037 114831 152047
rect 1066 151505 55123 151515
rect 1066 150959 218906 151505
rect 1066 150949 66531 150959
rect 1066 150417 49603 150427
rect 1066 149871 218906 150417
rect 1066 149861 9951 149871
rect 1066 149329 4996 149339
rect 1066 148783 218906 149329
rect 1066 148773 5088 148783
rect 1066 148241 21175 148251
rect 1066 147695 218906 148241
rect 1066 147685 62312 147695
rect 1066 147153 63587 147163
rect 1066 146607 218906 147153
rect 1066 146597 59079 146607
rect 1066 146065 13736 146075
rect 1066 145519 218906 146065
rect 1066 145509 5259 145519
rect 1066 144977 17955 144987
rect 1066 144431 218906 144977
rect 1066 144421 5548 144431
rect 1066 143889 11423 143899
rect 1066 143343 218906 143889
rect 1066 143333 25959 143343
rect 1066 142801 138199 142811
rect 1066 142255 218906 142801
rect 1066 142245 4904 142255
rect 1066 141713 23107 141723
rect 1066 141167 218906 141713
rect 1066 141157 5088 141167
rect 1066 140625 18047 140635
rect 1066 140079 218906 140625
rect 1066 140069 59644 140079
rect 1066 139537 6179 139547
rect 1066 138991 218906 139537
rect 1066 138981 70027 138991
rect 1066 138449 57068 138459
rect 1066 137903 218906 138449
rect 1066 137893 14275 137903
rect 1066 137361 55688 137371
rect 1066 136815 218906 137361
rect 1066 136805 4352 136815
rect 1066 136273 15116 136283
rect 1066 135727 218906 136273
rect 1066 135717 24763 135727
rect 1066 135185 21451 135195
rect 1066 134639 218906 135185
rect 1066 134629 5075 134639
rect 1066 134097 13092 134107
rect 1066 133551 218906 134097
rect 1066 133541 128000 133551
rect 1066 133009 145651 133019
rect 1066 132463 218906 133009
rect 1066 132453 70671 132463
rect 1066 131921 32399 131931
rect 1066 131375 218906 131921
rect 1066 131365 15103 131375
rect 1066 130833 61931 130843
rect 1066 130287 218906 130833
rect 1066 130277 50523 130287
rect 1066 129745 38944 129755
rect 1066 129199 218906 129745
rect 1066 129189 4168 129199
rect 1066 128657 15392 128667
rect 1066 128111 218906 128657
rect 1066 128101 4628 128111
rect 1066 127569 5259 127579
rect 1066 127023 218906 127569
rect 1066 127013 91923 127023
rect 1066 126481 4891 126491
rect 1066 125935 218906 126481
rect 1066 125925 5272 125935
rect 1066 125393 15116 125403
rect 1066 124847 218906 125393
rect 1066 124837 5640 124847
rect 1066 124305 5180 124315
rect 1066 123759 218906 124305
rect 1066 123749 86140 123759
rect 1066 123217 37840 123227
rect 1066 122671 218906 123217
rect 1066 122661 50983 122671
rect 1066 122129 86324 122139
rect 1066 121583 218906 122129
rect 1066 121573 99651 121583
rect 1066 121041 11331 121051
rect 1066 120495 218906 121041
rect 1066 120485 4996 120495
rect 1066 119953 26143 119963
rect 1066 119407 218906 119953
rect 1066 119397 17495 119407
rect 1066 118865 4812 118875
rect 1066 118319 218906 118865
rect 1066 118309 56319 118319
rect 1066 117777 86508 117787
rect 1066 117231 218906 117777
rect 1066 117221 5088 117231
rect 1066 116689 6455 116699
rect 1066 116143 218906 116689
rect 1066 116133 31295 116143
rect 1066 115601 9307 115611
rect 1066 115055 218906 115601
rect 1066 115045 28627 115055
rect 1066 114513 15195 114523
rect 1066 113967 218906 114513
rect 1066 113957 25867 113967
rect 1066 113425 59907 113435
rect 1066 112879 218906 113425
rect 1066 112869 4260 112879
rect 1066 112337 53099 112347
rect 1066 111791 218906 112337
rect 1066 111781 18139 111791
rect 1066 111249 15287 111259
rect 1066 110703 218906 111249
rect 1066 110693 9136 110703
rect 1066 110161 27339 110171
rect 1066 109615 218906 110161
rect 1066 109605 5259 109615
rect 1066 109073 5548 109083
rect 1066 108527 218906 109073
rect 1066 108517 86784 108527
rect 1066 107985 86508 107995
rect 1066 107439 218906 107985
rect 1066 107429 18704 107439
rect 1066 106897 7480 106907
rect 1066 106351 218906 106897
rect 1066 106341 3892 106351
rect 1066 105809 23475 105819
rect 1066 105263 218906 105809
rect 1066 105253 130747 105263
rect 1066 104721 36999 104731
rect 1066 104175 218906 104721
rect 1066 104165 38668 104175
rect 1066 103633 38011 103643
rect 1066 103087 218906 103633
rect 1066 103077 85851 103087
rect 1066 102545 38208 102555
rect 1066 101999 218906 102545
rect 1066 101989 85956 101999
rect 1066 101457 49156 101467
rect 1066 100911 218906 101457
rect 1066 100901 88887 100911
rect 1066 100369 63587 100379
rect 1066 99823 218906 100369
rect 1066 99813 48591 99823
rect 1066 99281 37932 99291
rect 1066 98735 218906 99281
rect 1066 98725 36723 98735
rect 1066 98193 86324 98203
rect 1066 97647 218906 98193
rect 1066 97637 85956 97647
rect 1066 97105 102227 97115
rect 1066 96559 218906 97105
rect 1066 96549 123019 96559
rect 1066 96017 12527 96027
rect 1066 95471 218906 96017
rect 1066 95461 4352 95471
rect 1066 94929 4707 94939
rect 1066 94383 218906 94929
rect 1066 94373 13907 94383
rect 1066 93841 4628 93851
rect 1066 93295 218906 93841
rect 1066 93285 120180 93295
rect 1066 92753 47868 92763
rect 1066 92207 218906 92753
rect 1066 92197 10411 92207
rect 1066 91665 21359 91675
rect 1066 91119 218906 91665
rect 1066 91109 4260 91119
rect 1066 90577 10779 90587
rect 1066 90031 218906 90577
rect 1066 90021 14643 90031
rect 1066 89489 11344 89499
rect 1066 88943 218906 89489
rect 1066 88933 18244 88943
rect 1066 88401 4628 88411
rect 1066 87855 218906 88401
rect 1066 87845 26800 87855
rect 1066 87313 48236 87323
rect 1066 86767 218906 87313
rect 1066 86757 13907 86767
rect 1066 86225 4720 86235
rect 1066 85679 218906 86225
rect 1066 85669 10700 85679
rect 1066 85137 28259 85147
rect 1066 84591 218906 85137
rect 1066 84581 7204 84591
rect 1066 84049 10595 84059
rect 1066 83503 218906 84049
rect 1066 83493 75376 83503
rect 1066 82961 93947 82971
rect 1066 82415 218906 82961
rect 1066 82405 5640 82415
rect 1066 81873 16943 81883
rect 1066 81327 218906 81873
rect 1066 81317 5259 81327
rect 1066 80785 28903 80795
rect 1066 80239 218906 80785
rect 1066 80229 10700 80239
rect 1066 79697 11068 79707
rect 1066 79151 218906 79697
rect 1066 79141 4628 79151
rect 1066 78609 23567 78619
rect 1066 78063 218906 78609
rect 1066 78053 97995 78063
rect 1066 77521 80252 77531
rect 1066 76975 218906 77521
rect 1066 76965 26800 76975
rect 1066 76433 10871 76443
rect 1066 75887 218906 76433
rect 1066 75877 18507 75887
rect 1066 75345 19795 75355
rect 1066 74799 218906 75345
rect 1066 74789 4260 74799
rect 1066 74257 14551 74267
rect 1066 73711 218906 74257
rect 1066 73701 4996 73711
rect 1066 73169 5088 73179
rect 1066 72623 218906 73169
rect 1066 72613 11068 72623
rect 1066 72081 20531 72091
rect 1066 71535 218906 72081
rect 1066 71525 4168 71535
rect 1066 70993 16943 71003
rect 1066 70447 218906 70993
rect 1066 70437 23015 70447
rect 1066 69905 49879 69915
rect 1066 69359 218906 69905
rect 1066 69349 40324 69359
rect 1066 68817 11344 68827
rect 1066 68271 218906 68817
rect 1066 68261 4076 68271
rect 1066 67729 10700 67739
rect 1066 67183 218906 67729
rect 1066 67173 190744 67183
rect 1066 66641 74364 66651
rect 1066 66095 218906 66641
rect 1066 66085 28443 66095
rect 1066 65553 4063 65563
rect 1066 65007 218906 65553
rect 1066 64997 4260 65007
rect 1066 64465 28719 64475
rect 1066 63919 218906 64465
rect 1066 63909 12803 63919
rect 1066 63377 13276 63387
rect 1066 62831 218906 63377
rect 1066 62821 4247 62831
rect 1066 62289 39956 62299
rect 1066 61743 218906 62289
rect 1066 61733 49892 61743
rect 1066 61201 13736 61211
rect 1066 60655 218906 61201
rect 1066 60645 4352 60655
rect 1066 60113 13092 60123
rect 1066 59567 218906 60113
rect 1066 59557 10884 59567
rect 1066 59025 54019 59035
rect 1066 58479 218906 59025
rect 1066 58469 40232 58479
rect 1066 57937 12724 57947
rect 1066 57391 218906 57937
rect 1066 57381 5259 57391
rect 1066 56849 4996 56859
rect 1066 56303 218906 56849
rect 1066 56293 13355 56303
rect 1066 55761 48959 55771
rect 1066 55215 218906 55761
rect 1066 55205 26235 55215
rect 1066 54673 29100 54683
rect 1066 54127 218906 54673
rect 1066 54117 5824 54127
rect 1066 53585 46580 53595
rect 1066 53039 218906 53585
rect 1066 53029 6915 53039
rect 1066 52497 18415 52507
rect 1066 51951 218906 52497
rect 1066 51941 3787 51951
rect 1066 50863 218906 51419
rect 1066 50853 3984 50863
rect 1066 50321 7927 50331
rect 1066 49775 218906 50321
rect 1066 49765 57239 49775
rect 1066 49233 50444 49243
rect 1066 48687 218906 49233
rect 1066 48677 40403 48687
rect 1066 48145 41336 48155
rect 1066 47599 218906 48145
rect 1066 47589 53927 47599
rect 1066 47057 106932 47067
rect 1066 46511 218906 47057
rect 1066 46501 190836 46511
rect 1066 45969 39956 45979
rect 1066 45423 218906 45969
rect 1066 45413 51732 45423
rect 1066 44881 39588 44891
rect 1066 44335 218906 44881
rect 1066 44325 46843 44335
rect 1066 43793 67175 43803
rect 1066 43247 218906 43793
rect 1066 43237 8032 43247
rect 1066 42705 13736 42715
rect 1066 42159 218906 42705
rect 1066 42149 7651 42159
rect 1066 41617 8216 41627
rect 1066 41071 218906 41617
rect 1066 41061 23291 41071
rect 1066 40529 8216 40539
rect 1066 39983 218906 40529
rect 1066 39973 42072 39983
rect 1066 39441 13171 39451
rect 1066 38895 218906 39441
rect 1066 38885 8032 38895
rect 1066 38353 7835 38363
rect 1066 37807 218906 38353
rect 1066 37797 7572 37807
rect 1066 37265 7927 37275
rect 1066 36719 218906 37265
rect 1066 36709 81172 36719
rect 1066 36177 8124 36187
rect 1066 35631 218906 36177
rect 1066 35621 27615 35631
rect 1066 35089 41520 35099
rect 1066 34543 218906 35089
rect 1066 34533 52376 34543
rect 1066 34001 49879 34011
rect 1066 33455 218906 34001
rect 1066 33445 77768 33455
rect 1066 32913 192847 32923
rect 1066 32367 218906 32913
rect 1066 32357 60919 32367
rect 1066 31825 43176 31835
rect 1066 31279 218906 31825
rect 1066 31269 41231 31279
rect 1066 30737 57147 30747
rect 1066 30191 218906 30737
rect 1066 30181 8308 30191
rect 1066 29649 7848 29659
rect 1066 29103 218906 29649
rect 1066 29093 20991 29103
rect 1066 28561 7467 28571
rect 1066 28015 218906 28561
rect 1066 28005 7375 28015
rect 1066 27473 12711 27483
rect 1066 26927 218906 27473
rect 1066 26917 7572 26927
rect 1066 26385 7756 26395
rect 1066 25839 218906 26385
rect 1066 25829 7572 25839
rect 1066 25297 25039 25307
rect 1066 24751 218906 25297
rect 1066 24741 7572 24751
rect 1066 24209 7835 24219
rect 1066 23663 218906 24209
rect 1066 23653 7572 23663
rect 1066 23121 8308 23131
rect 1066 22575 218906 23121
rect 1066 22565 12159 22575
rect 1066 22033 64875 22043
rect 1066 21487 218906 22033
rect 1066 21477 103436 21487
rect 1066 20945 117131 20955
rect 1066 20399 218906 20945
rect 1066 20389 55136 20399
rect 1066 19857 84747 19867
rect 1066 19311 218906 19857
rect 1066 19301 24027 19311
rect 1066 18769 28732 18779
rect 1066 18223 218906 18769
rect 1066 18213 61760 18223
rect 1066 17681 14827 17691
rect 1066 17135 218906 17681
rect 1066 17125 7283 17135
rect 1066 16593 7940 16603
rect 1066 16047 218906 16593
rect 1066 16037 10503 16047
rect 1066 15505 8032 15515
rect 1066 14959 218906 15505
rect 1066 14949 14275 14959
rect 1066 14417 7559 14427
rect 1066 13871 218906 14417
rect 1066 13861 7848 13871
rect 1066 13329 10871 13339
rect 1066 12783 218906 13329
rect 1066 12773 14827 12783
rect 1066 12241 8032 12251
rect 1066 11695 218906 12241
rect 1066 11685 10503 11695
rect 1066 11153 7848 11163
rect 1066 10607 218906 11153
rect 1066 10597 39943 10607
rect 1066 10065 7375 10075
rect 1066 9519 218906 10065
rect 1066 9509 20715 9519
rect 1066 8977 22476 8987
rect 1066 8431 218906 8977
rect 1066 8421 7664 8431
rect 1066 7889 7388 7899
rect 1066 7343 218906 7889
rect 1066 7333 7835 7343
rect 1066 6801 8032 6811
rect 1066 6255 218906 6801
rect 1066 6245 15944 6255
rect 1066 5713 165720 5723
rect 1066 5167 218906 5713
rect 1066 5157 180611 5167
rect 1066 4069 218906 4635
rect 1066 2981 218906 3547
rect 1066 2138 218906 2459
<< obsli1 >>
rect 1104 2159 219023 277457
<< obsm1 >>
rect 1104 1708 219035 277568
<< metal2 >>
rect 1306 279200 1362 280000
rect 3974 279200 4030 280000
rect 6734 279200 6790 280000
rect 9494 279200 9550 280000
rect 12254 279200 12310 280000
rect 15014 279200 15070 280000
rect 17774 279200 17830 280000
rect 20534 279200 20590 280000
rect 23294 279200 23350 280000
rect 25962 279200 26018 280000
rect 28722 279200 28778 280000
rect 31482 279200 31538 280000
rect 34242 279200 34298 280000
rect 37002 279200 37058 280000
rect 39762 279200 39818 280000
rect 42522 279200 42578 280000
rect 45282 279200 45338 280000
rect 48042 279200 48098 280000
rect 50710 279200 50766 280000
rect 53470 279200 53526 280000
rect 56230 279200 56286 280000
rect 58990 279200 59046 280000
rect 61750 279200 61806 280000
rect 64510 279200 64566 280000
rect 67270 279200 67326 280000
rect 70030 279200 70086 280000
rect 72790 279200 72846 280000
rect 75458 279200 75514 280000
rect 78218 279200 78274 280000
rect 80978 279200 81034 280000
rect 83738 279200 83794 280000
rect 86498 279200 86554 280000
rect 89258 279200 89314 280000
rect 92018 279200 92074 280000
rect 94778 279200 94834 280000
rect 97538 279200 97594 280000
rect 100206 279200 100262 280000
rect 102966 279200 103022 280000
rect 105726 279200 105782 280000
rect 108486 279200 108542 280000
rect 111246 279200 111302 280000
rect 114006 279200 114062 280000
rect 116766 279200 116822 280000
rect 119526 279200 119582 280000
rect 122286 279200 122342 280000
rect 124954 279200 125010 280000
rect 127714 279200 127770 280000
rect 130474 279200 130530 280000
rect 133234 279200 133290 280000
rect 135994 279200 136050 280000
rect 138754 279200 138810 280000
rect 141514 279200 141570 280000
rect 144274 279200 144330 280000
rect 147034 279200 147090 280000
rect 149702 279200 149758 280000
rect 152462 279200 152518 280000
rect 155222 279200 155278 280000
rect 157982 279200 158038 280000
rect 160742 279200 160798 280000
rect 163502 279200 163558 280000
rect 166262 279200 166318 280000
rect 169022 279200 169078 280000
rect 171782 279200 171838 280000
rect 174450 279200 174506 280000
rect 177210 279200 177266 280000
rect 179970 279200 180026 280000
rect 182730 279200 182786 280000
rect 185490 279200 185546 280000
rect 188250 279200 188306 280000
rect 191010 279200 191066 280000
rect 193770 279200 193826 280000
rect 196530 279200 196586 280000
rect 199198 279200 199254 280000
rect 201958 279200 202014 280000
rect 204718 279200 204774 280000
rect 207478 279200 207534 280000
rect 210238 279200 210294 280000
rect 212998 279200 213054 280000
rect 215758 279200 215814 280000
rect 218518 279200 218574 280000
<< obsm2 >>
rect 1418 279144 3918 279200
rect 4086 279144 6678 279200
rect 6846 279144 9438 279200
rect 9606 279144 12198 279200
rect 12366 279144 14958 279200
rect 15126 279144 17718 279200
rect 17886 279144 20478 279200
rect 20646 279144 23238 279200
rect 23406 279144 25906 279200
rect 26074 279144 28666 279200
rect 28834 279144 31426 279200
rect 31594 279144 34186 279200
rect 34354 279144 36946 279200
rect 37114 279144 39706 279200
rect 39874 279144 42466 279200
rect 42634 279144 45226 279200
rect 45394 279144 47986 279200
rect 48154 279144 50654 279200
rect 50822 279144 53414 279200
rect 53582 279144 56174 279200
rect 56342 279144 58934 279200
rect 59102 279144 61694 279200
rect 61862 279144 64454 279200
rect 64622 279144 67214 279200
rect 67382 279144 69974 279200
rect 70142 279144 72734 279200
rect 72902 279144 75402 279200
rect 75570 279144 78162 279200
rect 78330 279144 80922 279200
rect 81090 279144 83682 279200
rect 83850 279144 86442 279200
rect 86610 279144 89202 279200
rect 89370 279144 91962 279200
rect 92130 279144 94722 279200
rect 94890 279144 97482 279200
rect 97650 279144 100150 279200
rect 100318 279144 102910 279200
rect 103078 279144 105670 279200
rect 105838 279144 108430 279200
rect 108598 279144 111190 279200
rect 111358 279144 113950 279200
rect 114118 279144 116710 279200
rect 116878 279144 119470 279200
rect 119638 279144 122230 279200
rect 122398 279144 124898 279200
rect 125066 279144 127658 279200
rect 127826 279144 130418 279200
rect 130586 279144 133178 279200
rect 133346 279144 135938 279200
rect 136106 279144 138698 279200
rect 138866 279144 141458 279200
rect 141626 279144 144218 279200
rect 144386 279144 146978 279200
rect 147146 279144 149646 279200
rect 149814 279144 152406 279200
rect 152574 279144 155166 279200
rect 155334 279144 157926 279200
rect 158094 279144 160686 279200
rect 160854 279144 163446 279200
rect 163614 279144 166206 279200
rect 166374 279144 168966 279200
rect 169134 279144 171726 279200
rect 171894 279144 174394 279200
rect 174562 279144 177154 279200
rect 177322 279144 179914 279200
rect 180082 279144 182674 279200
rect 182842 279144 185434 279200
rect 185602 279144 188194 279200
rect 188362 279144 190954 279200
rect 191122 279144 193714 279200
rect 193882 279144 196474 279200
rect 196642 279144 199142 279200
rect 199310 279144 201902 279200
rect 202070 279144 204662 279200
rect 204830 279144 207422 279200
rect 207590 279144 210182 279200
rect 210350 279144 212942 279200
rect 213110 279144 215702 279200
rect 215870 279144 218462 279200
rect 218630 279144 218848 279200
rect 1308 1702 218848 279144
<< obsm3 >>
rect 1761 2143 218763 277473
<< metal4 >>
rect 4208 2128 4528 277488
rect 19568 2128 19888 277488
rect 34928 2128 35248 277488
rect 50288 2128 50608 277488
rect 65648 2128 65968 277488
rect 81008 2128 81328 277488
rect 96368 2128 96688 277488
rect 111728 2128 112048 277488
rect 127088 2128 127408 277488
rect 142448 2128 142768 277488
rect 157808 2128 158128 277488
rect 173168 2128 173488 277488
rect 188528 2128 188848 277488
rect 203888 2128 204208 277488
<< obsm4 >>
rect 9443 3979 19488 277133
rect 19968 3979 34848 277133
rect 35328 3979 50208 277133
rect 50688 3979 65568 277133
rect 66048 3979 80928 277133
rect 81408 3979 96288 277133
rect 96768 3979 111648 277133
rect 112128 3979 127008 277133
rect 127488 3979 142368 277133
rect 142848 3979 157728 277133
rect 158208 3979 173088 277133
rect 173568 3979 188448 277133
rect 188928 3979 203808 277133
rect 204288 3979 217981 277133
<< labels >>
rlabel metal2 s 89258 279200 89314 280000 6 A[0]
port 1 nsew signal input
rlabel metal2 s 92018 279200 92074 280000 6 A[1]
port 2 nsew signal input
rlabel metal2 s 94778 279200 94834 280000 6 A[2]
port 3 nsew signal input
rlabel metal2 s 97538 279200 97594 280000 6 A[3]
port 4 nsew signal input
rlabel metal2 s 100206 279200 100262 280000 6 A[4]
port 5 nsew signal input
rlabel metal2 s 102966 279200 103022 280000 6 A[5]
port 6 nsew signal input
rlabel metal2 s 105726 279200 105782 280000 6 A[6]
port 7 nsew signal input
rlabel metal2 s 108486 279200 108542 280000 6 A[7]
port 8 nsew signal input
rlabel metal2 s 111246 279200 111302 280000 6 A[8]
port 9 nsew signal input
rlabel metal2 s 114006 279200 114062 280000 6 A[9]
port 10 nsew signal input
rlabel metal2 s 116766 279200 116822 280000 6 CLK
port 11 nsew signal input
rlabel metal2 s 133234 279200 133290 280000 6 Di[0]
port 12 nsew signal input
rlabel metal2 s 160742 279200 160798 280000 6 Di[10]
port 13 nsew signal input
rlabel metal2 s 163502 279200 163558 280000 6 Di[11]
port 14 nsew signal input
rlabel metal2 s 166262 279200 166318 280000 6 Di[12]
port 15 nsew signal input
rlabel metal2 s 169022 279200 169078 280000 6 Di[13]
port 16 nsew signal input
rlabel metal2 s 171782 279200 171838 280000 6 Di[14]
port 17 nsew signal input
rlabel metal2 s 174450 279200 174506 280000 6 Di[15]
port 18 nsew signal input
rlabel metal2 s 177210 279200 177266 280000 6 Di[16]
port 19 nsew signal input
rlabel metal2 s 179970 279200 180026 280000 6 Di[17]
port 20 nsew signal input
rlabel metal2 s 182730 279200 182786 280000 6 Di[18]
port 21 nsew signal input
rlabel metal2 s 185490 279200 185546 280000 6 Di[19]
port 22 nsew signal input
rlabel metal2 s 135994 279200 136050 280000 6 Di[1]
port 23 nsew signal input
rlabel metal2 s 188250 279200 188306 280000 6 Di[20]
port 24 nsew signal input
rlabel metal2 s 191010 279200 191066 280000 6 Di[21]
port 25 nsew signal input
rlabel metal2 s 193770 279200 193826 280000 6 Di[22]
port 26 nsew signal input
rlabel metal2 s 196530 279200 196586 280000 6 Di[23]
port 27 nsew signal input
rlabel metal2 s 199198 279200 199254 280000 6 Di[24]
port 28 nsew signal input
rlabel metal2 s 201958 279200 202014 280000 6 Di[25]
port 29 nsew signal input
rlabel metal2 s 204718 279200 204774 280000 6 Di[26]
port 30 nsew signal input
rlabel metal2 s 207478 279200 207534 280000 6 Di[27]
port 31 nsew signal input
rlabel metal2 s 210238 279200 210294 280000 6 Di[28]
port 32 nsew signal input
rlabel metal2 s 212998 279200 213054 280000 6 Di[29]
port 33 nsew signal input
rlabel metal2 s 138754 279200 138810 280000 6 Di[2]
port 34 nsew signal input
rlabel metal2 s 215758 279200 215814 280000 6 Di[30]
port 35 nsew signal input
rlabel metal2 s 218518 279200 218574 280000 6 Di[31]
port 36 nsew signal input
rlabel metal2 s 141514 279200 141570 280000 6 Di[3]
port 37 nsew signal input
rlabel metal2 s 144274 279200 144330 280000 6 Di[4]
port 38 nsew signal input
rlabel metal2 s 147034 279200 147090 280000 6 Di[5]
port 39 nsew signal input
rlabel metal2 s 149702 279200 149758 280000 6 Di[6]
port 40 nsew signal input
rlabel metal2 s 152462 279200 152518 280000 6 Di[7]
port 41 nsew signal input
rlabel metal2 s 155222 279200 155278 280000 6 Di[8]
port 42 nsew signal input
rlabel metal2 s 157982 279200 158038 280000 6 Di[9]
port 43 nsew signal input
rlabel metal2 s 1306 279200 1362 280000 6 Do[0]
port 44 nsew signal output
rlabel metal2 s 28722 279200 28778 280000 6 Do[10]
port 45 nsew signal output
rlabel metal2 s 31482 279200 31538 280000 6 Do[11]
port 46 nsew signal output
rlabel metal2 s 34242 279200 34298 280000 6 Do[12]
port 47 nsew signal output
rlabel metal2 s 37002 279200 37058 280000 6 Do[13]
port 48 nsew signal output
rlabel metal2 s 39762 279200 39818 280000 6 Do[14]
port 49 nsew signal output
rlabel metal2 s 42522 279200 42578 280000 6 Do[15]
port 50 nsew signal output
rlabel metal2 s 45282 279200 45338 280000 6 Do[16]
port 51 nsew signal output
rlabel metal2 s 48042 279200 48098 280000 6 Do[17]
port 52 nsew signal output
rlabel metal2 s 50710 279200 50766 280000 6 Do[18]
port 53 nsew signal output
rlabel metal2 s 53470 279200 53526 280000 6 Do[19]
port 54 nsew signal output
rlabel metal2 s 3974 279200 4030 280000 6 Do[1]
port 55 nsew signal output
rlabel metal2 s 56230 279200 56286 280000 6 Do[20]
port 56 nsew signal output
rlabel metal2 s 58990 279200 59046 280000 6 Do[21]
port 57 nsew signal output
rlabel metal2 s 61750 279200 61806 280000 6 Do[22]
port 58 nsew signal output
rlabel metal2 s 64510 279200 64566 280000 6 Do[23]
port 59 nsew signal output
rlabel metal2 s 67270 279200 67326 280000 6 Do[24]
port 60 nsew signal output
rlabel metal2 s 70030 279200 70086 280000 6 Do[25]
port 61 nsew signal output
rlabel metal2 s 72790 279200 72846 280000 6 Do[26]
port 62 nsew signal output
rlabel metal2 s 75458 279200 75514 280000 6 Do[27]
port 63 nsew signal output
rlabel metal2 s 78218 279200 78274 280000 6 Do[28]
port 64 nsew signal output
rlabel metal2 s 80978 279200 81034 280000 6 Do[29]
port 65 nsew signal output
rlabel metal2 s 6734 279200 6790 280000 6 Do[2]
port 66 nsew signal output
rlabel metal2 s 83738 279200 83794 280000 6 Do[30]
port 67 nsew signal output
rlabel metal2 s 86498 279200 86554 280000 6 Do[31]
port 68 nsew signal output
rlabel metal2 s 9494 279200 9550 280000 6 Do[3]
port 69 nsew signal output
rlabel metal2 s 12254 279200 12310 280000 6 Do[4]
port 70 nsew signal output
rlabel metal2 s 15014 279200 15070 280000 6 Do[5]
port 71 nsew signal output
rlabel metal2 s 17774 279200 17830 280000 6 Do[6]
port 72 nsew signal output
rlabel metal2 s 20534 279200 20590 280000 6 Do[7]
port 73 nsew signal output
rlabel metal2 s 23294 279200 23350 280000 6 Do[8]
port 74 nsew signal output
rlabel metal2 s 25962 279200 26018 280000 6 Do[9]
port 75 nsew signal output
rlabel metal2 s 130474 279200 130530 280000 6 EN
port 76 nsew signal input
rlabel metal2 s 119526 279200 119582 280000 6 WE[0]
port 77 nsew signal input
rlabel metal2 s 122286 279200 122342 280000 6 WE[1]
port 78 nsew signal input
rlabel metal2 s 124954 279200 125010 280000 6 WE[2]
port 79 nsew signal input
rlabel metal2 s 127714 279200 127770 280000 6 WE[3]
port 80 nsew signal input
rlabel metal4 s 188528 2128 188848 277488 6 vccd1
port 81 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 277488 6 vccd1
port 82 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 277488 6 vccd1
port 83 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 277488 6 vccd1
port 84 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 277488 6 vccd1
port 85 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 277488 6 vccd1
port 86 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 277488 6 vccd1
port 87 nsew power bidirectional
rlabel metal4 s 203888 2128 204208 277488 6 vssd1
port 88 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 277488 6 vssd1
port 89 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 277488 6 vssd1
port 90 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 277488 6 vssd1
port 91 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 277488 6 vssd1
port 92 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 277488 6 vssd1
port 93 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 277488 6 vssd1
port 94 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 220000 280000
string LEFview TRUE
string GDS_FILE /project/openlane/DFFRAM_1Kx32/runs/DFFRAM_1Kx32/results/magic/DFFRAM_1Kx32.gds
string GDS_END 238362704
string GDS_START 181870
<< end >>

