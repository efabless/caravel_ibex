* NGSPICE file created from apb_sys_0.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd1_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_1 abstract view
.subckt sky130_fd_sc_hd__clkinv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_1 abstract view
.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_16 abstract view
.subckt sky130_fd_sc_hd__inv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_2 abstract view
.subckt sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_2 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4bb_2 abstract view
.subckt sky130_fd_sc_hd__nand4bb_2 A_N B_N C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_16 abstract view
.subckt sky130_fd_sc_hd__clkinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4bb_4 abstract view
.subckt sky130_fd_sc_hd__nand4bb_4 A_N B_N C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

.subckt apb_sys_0 HADDR[0] HADDR[10] HADDR[11] HADDR[12] HADDR[13] HADDR[14] HADDR[15]
+ HADDR[16] HADDR[17] HADDR[18] HADDR[19] HADDR[1] HADDR[20] HADDR[21] HADDR[22] HADDR[23]
+ HADDR[24] HADDR[25] HADDR[26] HADDR[27] HADDR[28] HADDR[29] HADDR[2] HADDR[30] HADDR[31]
+ HADDR[3] HADDR[4] HADDR[5] HADDR[6] HADDR[7] HADDR[8] HADDR[9] HCLK HRDATA[0] HRDATA[10]
+ HRDATA[11] HRDATA[12] HRDATA[13] HRDATA[14] HRDATA[15] HRDATA[16] HRDATA[17] HRDATA[18]
+ HRDATA[19] HRDATA[1] HRDATA[20] HRDATA[21] HRDATA[22] HRDATA[23] HRDATA[24] HRDATA[25]
+ HRDATA[26] HRDATA[27] HRDATA[28] HRDATA[29] HRDATA[2] HRDATA[30] HRDATA[31] HRDATA[3]
+ HRDATA[4] HRDATA[5] HRDATA[6] HRDATA[7] HRDATA[8] HRDATA[9] HREADY HREADYOUT HRESETn
+ HSEL HTRANS[0] HTRANS[1] HWDATA[0] HWDATA[10] HWDATA[11] HWDATA[12] HWDATA[13] HWDATA[14]
+ HWDATA[15] HWDATA[16] HWDATA[17] HWDATA[18] HWDATA[19] HWDATA[1] HWDATA[20] HWDATA[21]
+ HWDATA[22] HWDATA[23] HWDATA[24] HWDATA[25] HWDATA[26] HWDATA[27] HWDATA[28] HWDATA[29]
+ HWDATA[2] HWDATA[30] HWDATA[31] HWDATA[3] HWDATA[4] HWDATA[5] HWDATA[6] HWDATA[7]
+ HWDATA[8] HWDATA[9] HWRITE IRQ[0] IRQ[10] IRQ[11] IRQ[12] IRQ[13] IRQ[14] IRQ[15]
+ IRQ[1] IRQ[2] IRQ[3] IRQ[4] IRQ[5] IRQ[6] IRQ[7] IRQ[8] IRQ[9] MSI_S2 MSI_S3 MSO_S2
+ MSO_S3 RsRx_S0 RsRx_S1 RsTx_S0 RsTx_S1 SCLK_S2 SCLK_S3 SSn_S2 SSn_S3 pwm_S6 pwm_S7
+ scl_i_S4 scl_i_S5 scl_o_S4 scl_o_S5 scl_oen_o_S4 scl_oen_o_S5 sda_i_S4 sda_i_S5
+ sda_o_S4 sda_o_S5 sda_oen_o_S4 sda_oen_o_S5 vccd1 vssd1
XFILLER_228_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09671_ _19428_/Q vssd1 vssd1 vccd1 vccd1 _09671_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15057__B1 _15020_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18869_ _18869_/CLK _18869_/D repeater195/X vssd1 vssd1 vccd1 vccd1 _18869_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_94_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_242_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17521__S _17539_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15830__A _15830_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16557__B1 _17108_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16645__B _16647_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19175__RESET_B repeater212/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09105_ _12238_/A vssd1 vssd1 vccd1 vccd1 _09105_/X sky130_fd_sc_hd__buf_4
XFILLER_108_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09036_ _20115_/Q _09029_/X hold305/X _09031_/X vssd1 vssd1 vccd1 vccd1 _20115_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_190_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold340 hold360/X vssd1 vssd1 vccd1 vccd1 hold359/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_123_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold351 hold351/A vssd1 vssd1 vccd1 vccd1 hold351/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold362 hold362/A vssd1 vssd1 vccd1 vccd1 hold362/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17904__S0 _19633_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold373 hold373/A vssd1 vssd1 vccd1 vccd1 hold373/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09938_ _19339_/Q vssd1 vssd1 vccd1 vccd1 _16472_/A sky130_fd_sc_hd__inv_2
XFILLER_219_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20058_ _20058_/CLK _20058_/D repeater194/X vssd1 vssd1 vccd1 vccd1 _20058_/Q sky130_fd_sc_hd__dfrtp_1
X_09869_ _09869_/A _09869_/B vssd1 vssd1 vccd1 vccd1 _09963_/A sky130_fd_sc_hd__or2_1
XFILLER_219_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11900_ _19417_/Q _11898_/X hold276/X _11899_/X vssd1 vssd1 vccd1 vccd1 _19417_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16796__A0 _15963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12880_ _12965_/A _12988_/A vssd1 vssd1 vccd1 vccd1 _12881_/B sky130_fd_sc_hd__or2_1
XFILLER_18_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater190 repeater191/X vssd1 vssd1 vccd1 vccd1 repeater190/X sky130_fd_sc_hd__buf_6
XFILLER_93_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11831_ _12371_/A _16234_/A vssd1 vssd1 vccd1 vccd1 _12558_/B sky130_fd_sc_hd__or2_4
XPHY_4344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19945__RESET_B repeater244/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17431__S _17566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14550_ _18312_/Q _14546_/X _14535_/X _14548_/X vssd1 vssd1 vccd1 vccd1 _18312_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11762_ hold162/X _11757_/X _19482_/Q _11758_/X vssd1 vssd1 vccd1 vccd1 hold164/A
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12282__B1 _12104_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13501_ _18764_/Q vssd1 vssd1 vccd1 vccd1 _14629_/B sky130_fd_sc_hd__buf_1
XFILLER_199_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10713_ _15404_/A _10704_/B _15753_/A _10712_/Y _10716_/S vssd1 vssd1 vccd1 vccd1
+ _10714_/A sky130_fd_sc_hd__o32a_1
XPHY_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14481_ _18353_/Q _14478_/X _12714_/X _14480_/X vssd1 vssd1 vccd1 vccd1 _18353_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11693_ _19528_/Q _11690_/X _10877_/X _11692_/X vssd1 vssd1 vccd1 vccd1 _19528_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10884__A hold245/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16220_ _19689_/Q vssd1 vssd1 vccd1 vccd1 _16220_/Y sky130_fd_sc_hd__inv_2
XPHY_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13432_ _19260_/Q _13445_/A vssd1 vssd1 vccd1 vccd1 _13432_/X sky130_fd_sc_hd__or2_1
XPHY_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10644_ _19784_/Q _10644_/B vssd1 vssd1 vccd1 vccd1 _10645_/B sky130_fd_sc_hd__or2_1
XPHY_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11388__A2 _19143_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16151_ _15846_/X _16131_/X _15859_/X _16140_/X _16150_/X vssd1 vssd1 vccd1 vccd1
+ _16151_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_6_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10575_ _10575_/A _10574_/X vssd1 vssd1 vccd1 vccd1 _10614_/A sky130_fd_sc_hd__or2b_1
X_13363_ _20116_/Q _13433_/A _13362_/Y _18862_/Q vssd1 vssd1 vccd1 vccd1 _13363_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_139_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrebuffer7 _13077_/B vssd1 vssd1 vccd1 vccd1 _13188_/B1 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_182_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15102_ _17989_/Q _15095_/X _14812_/A _15097_/X vssd1 vssd1 vccd1 vccd1 _17989_/D
+ sky130_fd_sc_hd__a22o_1
X_12314_ _15774_/A _12316_/B vssd1 vssd1 vccd1 vccd1 _12315_/S sky130_fd_sc_hd__or2_1
X_16082_ _17989_/Q vssd1 vssd1 vccd1 vccd1 _16082_/Y sky130_fd_sc_hd__inv_2
X_13294_ _14366_/B _13291_/Y _13293_/X vssd1 vssd1 vccd1 vccd1 _13294_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_181_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18898__RESET_B repeater188/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19910_ _20006_/CLK _19910_/D repeater191/X vssd1 vssd1 vccd1 vccd1 _19910_/Q sky130_fd_sc_hd__dfrtp_1
X_15033_ _18034_/Q _15024_/A _15020_/X _15025_/A vssd1 vssd1 vccd1 vccd1 _18034_/D
+ sky130_fd_sc_hd__a22o_1
X_12245_ _15232_/A _15232_/B _12247_/A vssd1 vssd1 vccd1 vccd1 _12245_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__18827__RESET_B repeater217/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19841_ _19841_/CLK _19841_/D repeater270/X vssd1 vssd1 vccd1 vccd1 _19841_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_111_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12176_ _19265_/Q _12171_/X _11920_/X _12172_/X vssd1 vssd1 vccd1 vccd1 _19265_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_1_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11127_ _11127_/A _11127_/B vssd1 vssd1 vccd1 vccd1 _19633_/D sky130_fd_sc_hd__nor2_1
X_19772_ _19772_/CLK _19772_/D repeater189/X vssd1 vssd1 vccd1 vccd1 _19772_/Q sky130_fd_sc_hd__dfstp_2
X_16984_ _17824_/X _19902_/Q _16986_/S vssd1 vssd1 vccd1 vccd1 _16984_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11058_ _11056_/A _14316_/B _11056_/Y vssd1 vssd1 vccd1 vccd1 _19641_/D sky130_fd_sc_hd__a21oi_1
X_15935_ _19843_/Q vssd1 vssd1 vccd1 vccd1 _15935_/Y sky130_fd_sc_hd__inv_2
X_18723_ _18727_/CLK _18723_/D repeater253/X vssd1 vssd1 vccd1 vccd1 _18723_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15039__B1 _14996_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10009_ _10009_/A _10009_/B vssd1 vssd1 vccd1 vccd1 _10048_/A sky130_fd_sc_hd__or2_1
X_18654_ _20048_/CLK _18654_/D repeater209/X vssd1 vssd1 vccd1 vccd1 _18654_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_237_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15866_ _15866_/A vssd1 vssd1 vccd1 vccd1 _15867_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__16787__A0 _17473_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14817_ _18163_/Q _14803_/A _14816_/X _14804_/A vssd1 vssd1 vccd1 vccd1 _18163_/D
+ sky130_fd_sc_hd__a22o_1
X_17605_ _13285_/B _13283_/C _17605_/S vssd1 vssd1 vccd1 vccd1 _17605_/X sky130_fd_sc_hd__mux2_1
X_18585_ _19470_/CLK _18585_/D repeater272/X vssd1 vssd1 vccd1 vccd1 _18585_/Q sky130_fd_sc_hd__dfrtp_1
X_15797_ _18042_/Q vssd1 vssd1 vccd1 vccd1 _15797_/Y sky130_fd_sc_hd__inv_2
XFILLER_240_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17341__S _17568_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17536_ _17535_/X _13528_/A _17536_/S vssd1 vssd1 vccd1 vccd1 _17536_/X sky130_fd_sc_hd__mux2_4
XFILLER_205_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12273__B1 _12088_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14748_ _18201_/Q _14744_/X _14745_/X _14747_/X vssd1 vssd1 vccd1 vccd1 _18201_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16539__B1 _17166_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17467_ _17466_/X _17889_/X _17568_/S vssd1 vssd1 vccd1 vccd1 _17467_/X sky130_fd_sc_hd__mux2_2
XFILLER_220_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14679_ _18234_/Q _14670_/A _14626_/X _14671_/A vssd1 vssd1 vccd1 vccd1 _18234_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_32_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16418_ _18097_/Q vssd1 vssd1 vccd1 vccd1 _16418_/Y sky130_fd_sc_hd__inv_2
X_19206_ _19585_/CLK _19206_/D hold365/X vssd1 vssd1 vccd1 vccd1 _19206_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12025__B1 hold276/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17398_ _17397_/X _16200_/X _17567_/S vssd1 vssd1 vccd1 vccd1 _17398_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19137_ _19137_/CLK _19137_/D hold348/X vssd1 vssd1 vccd1 vccd1 _19137_/Q sky130_fd_sc_hd__dfrtp_4
X_16349_ _17951_/Q vssd1 vssd1 vccd1 vccd1 _16349_/Y sky130_fd_sc_hd__inv_2
X_19068_ _19109_/CLK _19068_/D hold361/X vssd1 vssd1 vccd1 vccd1 _19068_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_218_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10018__B _10039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18019_ _18142_/CLK _18019_/D vssd1 vssd1 vccd1 vccd1 _18019_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13525__B1 _18761_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09807__B _09807_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18568__RESET_B repeater272/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15825__A _19685_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17516__S _17539_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09723_ _19414_/Q vssd1 vssd1 vccd1 vccd1 _09723_/Y sky130_fd_sc_hd__inv_2
XANTENNA__10969__A _12053_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09654_ _09749_/A _09748_/A _09741_/A _09740_/A vssd1 vssd1 vccd1 vccd1 _09660_/C
+ sky130_fd_sc_hd__or4_4
XFILLER_67_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16242__A2 _16638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_242_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09585_ _09585_/A vssd1 vssd1 vccd1 vccd1 _09585_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_82_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17251__S _17529_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12264__B1 _12069_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19356__RESET_B hold371/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14176__A _19113_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14556__A2 _14547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10360_ _10360_/A vssd1 vssd1 vccd1 vccd1 _19861_/D sky130_fd_sc_hd__inv_2
XFILLER_12_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09019_ _09043_/A vssd1 vssd1 vccd1 vccd1 _09019_/X sky130_fd_sc_hd__buf_1
XFILLER_191_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10291_ _18643_/Q _10291_/B vssd1 vssd1 vccd1 vccd1 _10291_/X sky130_fd_sc_hd__and2_1
XFILLER_2_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17258__A1 _19210_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12030_ _12030_/A vssd1 vssd1 vccd1 vccd1 _12030_/X sky130_fd_sc_hd__buf_4
Xhold170 hold170/A vssd1 vssd1 vccd1 vccd1 hold170/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 HADDR[8] vssd1 vssd1 vccd1 vccd1 input31/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 hold192/A vssd1 vssd1 vccd1 vccd1 hold192/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17426__S _17548_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10750__B1 _10425_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13981_ _18693_/Q vssd1 vssd1 vccd1 vccd1 _14023_/A sky130_fd_sc_hd__inv_2
XFILLER_18_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13255__A _18752_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15720_ _15727_/B vssd1 vssd1 vccd1 vccd1 _15725_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__16769__A0 _15768_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12932_ _12929_/Y _18947_/Q _12930_/Y _18923_/Q _12931_/Y vssd1 vssd1 vccd1 vccd1
+ _12941_/B sky130_fd_sc_hd__o221a_1
XFILLER_37_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15651_ _18605_/Q _15649_/C _18606_/Q vssd1 vssd1 vccd1 vccd1 _15651_/X sky130_fd_sc_hd__o21a_1
XFILLER_234_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12863_ _18919_/Q vssd1 vssd1 vccd1 vccd1 _12864_/A sky130_fd_sc_hd__inv_2
XPHY_4141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17161__S _17482_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14602_ _14602_/A vssd1 vssd1 vccd1 vccd1 _14602_/X sky130_fd_sc_hd__clkbuf_2
XPHY_4163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18370_ _19515_/CLK _18370_/D vssd1 vssd1 vccd1 vccd1 _18370_/Q sky130_fd_sc_hd__dfxtp_1
X_11814_ _11821_/A vssd1 vssd1 vccd1 vccd1 _11814_/X sky130_fd_sc_hd__clkbuf_2
XPHY_4174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15582_ _15584_/A _15581_/X _15702_/A vssd1 vssd1 vccd1 vccd1 _15582_/Y sky130_fd_sc_hd__a21oi_1
XPHY_4185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12794_ _19250_/Q _13550_/A _12793_/Y _18816_/Q vssd1 vssd1 vccd1 vccd1 _12794_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15992__B2 _15915_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17321_ _17486_/A0 _09908_/Y _17543_/S vssd1 vssd1 vccd1 vccd1 _17321_/X sky130_fd_sc_hd__mux2_1
XFILLER_202_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14533_ _14533_/A vssd1 vssd1 vccd1 vccd1 _14533_/X sky130_fd_sc_hd__clkbuf_2
XPHY_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11745_ _19495_/Q _11730_/A _16927_/X _11731_/A vssd1 vssd1 vccd1 vccd1 hold262/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17194__A0 _15768_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_230_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17252_ _17251_/X _20021_/Q _17482_/S vssd1 vssd1 vccd1 vccd1 _17252_/X sky130_fd_sc_hd__mux2_2
XANTENNA__12007__B1 _09025_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_230_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14464_ _14464_/A vssd1 vssd1 vccd1 vccd1 _14465_/A sky130_fd_sc_hd__inv_2
XPHY_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11676_ _10732_/B _11674_/X _10493_/A _11675_/X vssd1 vssd1 vccd1 vccd1 _19541_/D
+ sky130_fd_sc_hd__o22ai_1
XPHY_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16203_ _17941_/Q _16344_/B vssd1 vssd1 vccd1 vccd1 _16203_/Y sky130_fd_sc_hd__nand2_1
XFILLER_128_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13415_ _20114_/Q _13431_/C _13414_/Y _18860_/Q vssd1 vssd1 vccd1 vccd1 _13415_/X
+ sky130_fd_sc_hd__o22a_1
X_10627_ _10627_/A vssd1 vssd1 vccd1 vccd1 _19806_/D sky130_fd_sc_hd__inv_2
XFILLER_186_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17183_ _17182_/X _14077_/Y _17490_/S vssd1 vssd1 vccd1 vccd1 _17183_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14395_ _14395_/A vssd1 vssd1 vccd1 vccd1 _14396_/A sky130_fd_sc_hd__inv_2
XANTENNA_repeater244_A repeater245/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16134_ _19759_/Q vssd1 vssd1 vccd1 vccd1 _16134_/Y sky130_fd_sc_hd__inv_2
X_13346_ _13431_/D _13346_/B vssd1 vssd1 vccd1 vccd1 _13442_/A sky130_fd_sc_hd__or2_1
XFILLER_127_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10558_ _19806_/Q _10558_/B _10581_/C vssd1 vssd1 vccd1 vccd1 _10614_/C sky130_fd_sc_hd__nor3_4
XFILLER_142_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16065_ _15390_/Y _16049_/X _16059_/Y _15836_/X _16064_/X vssd1 vssd1 vccd1 vccd1
+ _16065_/X sky130_fd_sc_hd__o221a_2
X_13277_ _18750_/Q _13276_/Y _18750_/Q _13276_/Y vssd1 vssd1 vccd1 vccd1 _13299_/A
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__12334__A _12334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10489_ _10501_/C _10517_/A vssd1 vssd1 vccd1 vccd1 _11654_/A sky130_fd_sc_hd__or2_1
X_15016_ _18046_/Q _15010_/X _15000_/X _15012_/X vssd1 vssd1 vccd1 vccd1 _18046_/D
+ sky130_fd_sc_hd__a22o_1
X_12228_ _12228_/A vssd1 vssd1 vccd1 vccd1 _12228_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_97_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12053__B _12053_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17336__S _17546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19824_ _19825_/CLK _19824_/D repeater229/X vssd1 vssd1 vccd1 vccd1 _19824_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_151_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12159_ _19278_/Q _12157_/X _12107_/X _12158_/X vssd1 vssd1 vccd1 vccd1 _19278_/D
+ sky130_fd_sc_hd__a22o_1
X_19755_ _19825_/CLK _19755_/D repeater229/X vssd1 vssd1 vccd1 vccd1 _19755_/Q sky130_fd_sc_hd__dfrtp_1
X_16967_ _16671_/Y _19425_/Q _17459_/S vssd1 vssd1 vccd1 vccd1 _16967_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18706_ _19224_/CLK _18706_/D repeater186/X vssd1 vssd1 vccd1 vccd1 _18706_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12494__B1 _12380_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15918_ _15918_/A _15918_/B _15918_/C _15918_/D vssd1 vssd1 vccd1 vccd1 _15918_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_204_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19686_ _20049_/CLK _19686_/D repeater202/X vssd1 vssd1 vccd1 vccd1 _19686_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_76_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16898_ _16897_/X _16708_/Y _17512_/S vssd1 vssd1 vccd1 vccd1 _16898_/X sky130_fd_sc_hd__mux2_1
XFILLER_237_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18637_ _19813_/CLK _18637_/D repeater224/X vssd1 vssd1 vccd1 vccd1 _18637_/Q sky130_fd_sc_hd__dfrtp_2
X_15849_ _19756_/Q vssd1 vssd1 vccd1 vccd1 _15849_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17071__S _17493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09370_ _20007_/Q vssd1 vssd1 vccd1 vccd1 _09468_/A sky130_fd_sc_hd__inv_2
XFILLER_212_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18568_ _19841_/CLK _18568_/D repeater272/X vssd1 vssd1 vccd1 vccd1 _18568_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_220_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17185__A0 _15768_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17519_ _15875_/Y _09807_/B _17537_/S vssd1 vssd1 vccd1 vccd1 _17519_/X sky130_fd_sc_hd__mux2_1
X_18499_ _19794_/CLK _18499_/D repeater219/X vssd1 vssd1 vccd1 vccd1 _18499_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_220_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17246__S _17487_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16463__A2 _16148_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_157_HCLK_A clkbuf_4_0_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09706_ _09788_/A _19405_/Q _09629_/A _19429_/Q vssd1 vssd1 vccd1 vccd1 _09706_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12485__B1 _12238_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09637_ _19978_/Q vssd1 vssd1 vccd1 vccd1 _09790_/A sky130_fd_sc_hd__inv_2
XFILLER_216_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12237__B1 _12236_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09568_ _20035_/Q _09495_/Y _09496_/Y _09495_/A _09567_/X vssd1 vssd1 vccd1 vccd1
+ _20035_/D sky130_fd_sc_hd__o221a_1
XANTENNA__19190__RESET_B repeater244/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold337_A HWDATA[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09102__B1 _09101_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17176__A0 _17486_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09499_ _09496_/Y _19325_/Q _20013_/Q _09497_/Y _09498_/X vssd1 vssd1 vccd1 vccd1
+ _09512_/A sky130_fd_sc_hd__o221a_1
XPHY_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11530_ _11468_/B _11530_/A2 _19587_/Q _11529_/Y _11490_/X vssd1 vssd1 vccd1 vccd1
+ _19587_/D sky130_fd_sc_hd__o221a_1
XPHY_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11461_ _11461_/A _11461_/B vssd1 vssd1 vccd1 vccd1 _11538_/A sky130_fd_sc_hd__or2_1
XPHY_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13200_ _13200_/A vssd1 vssd1 vccd1 vccd1 _13200_/Y sky130_fd_sc_hd__clkinv_1
X_10412_ _14681_/A _15197_/A vssd1 vssd1 vccd1 vccd1 _10413_/S sky130_fd_sc_hd__or2_1
XFILLER_137_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14180_ _19118_/Q vssd1 vssd1 vccd1 vccd1 _14180_/Y sky130_fd_sc_hd__inv_2
X_11392_ _19555_/Q vssd1 vssd1 vccd1 vccd1 _11625_/A sky130_fd_sc_hd__inv_2
XFILLER_180_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13131_ _19163_/Q vssd1 vssd1 vccd1 vccd1 _13131_/Y sky130_fd_sc_hd__inv_2
XFILLER_164_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10343_ _10343_/A vssd1 vssd1 vccd1 vccd1 _10344_/B sky130_fd_sc_hd__inv_2
XANTENNA__09708__A2 _19421_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10274_ _19643_/Q vssd1 vssd1 vccd1 vccd1 _14317_/B sky130_fd_sc_hd__buf_1
X_13062_ _13062_/A _13062_/B vssd1 vssd1 vccd1 vccd1 _13210_/A sky130_fd_sc_hd__or2_1
XANTENNA__17156__S _17534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12013_ _19355_/Q _12009_/X hold305/X _12010_/X vssd1 vssd1 vccd1 vccd1 _19355_/D
+ sky130_fd_sc_hd__a22o_1
X_17870_ _16152_/Y _16153_/Y _16154_/Y _16155_/Y _17913_/S0 _19632_/Q vssd1 vssd1
+ vccd1 vccd1 _17870_/X sky130_fd_sc_hd__mux4_2
XFILLER_105_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10723__B1 _10446_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_238_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16821_ _16820_/X _13078_/A _17542_/S vssd1 vssd1 vccd1 vccd1 _16821_/X sky130_fd_sc_hd__mux2_2
XFILLER_65_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16995__S _17545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19540_ _19540_/CLK _19540_/D repeater221/X vssd1 vssd1 vccd1 vccd1 _19540_/Q sky130_fd_sc_hd__dfrtp_4
X_16752_ _20058_/Q _19741_/Q vssd1 vssd1 vccd1 vccd1 _16752_/X sky130_fd_sc_hd__and2_2
XFILLER_19_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11279__B2 _19018_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12476__B1 _12225_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13964_ _13964_/A _13964_/B _13964_/C vssd1 vssd1 vccd1 vccd1 _13967_/A sky130_fd_sc_hd__or3_4
XFILLER_246_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09341__A0 _09339_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15703_ _18619_/Q vssd1 vssd1 vccd1 vccd1 _15703_/Y sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_16_HCLK_A clkbuf_4_3_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12915_ _19270_/Q _18927_/Q _19270_/Q _18927_/Q vssd1 vssd1 vccd1 vccd1 _12915_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_206_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19471_ _19515_/CLK hold195/X repeater260/X vssd1 vssd1 vccd1 vccd1 _19471_/Q sky130_fd_sc_hd__dfrtp_1
X_16683_ _16683_/A vssd1 vssd1 vccd1 vccd1 _16683_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__14217__A1 _19110_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13895_ _19208_/Q _13911_/A _13894_/Y _18735_/Q vssd1 vssd1 vccd1 vccd1 _13895_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA_clkbuf_leaf_79_HCLK_A clkbuf_4_13_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16611__C1 _16610_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18422_ _18441_/CLK _18422_/D vssd1 vssd1 vccd1 vccd1 _18422_/Q sky130_fd_sc_hd__dfxtp_1
X_15634_ _15666_/A _15634_/B vssd1 vssd1 vccd1 vccd1 _15634_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_4_HCLK_A clkbuf_4_0_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12846_ _18938_/Q vssd1 vssd1 vccd1 vccd1 _12965_/A sky130_fd_sc_hd__inv_4
XFILLER_234_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18353_ _18959_/CLK _18353_/D vssd1 vssd1 vccd1 vccd1 _18353_/Q sky130_fd_sc_hd__dfxtp_1
X_15565_ _18585_/Q vssd1 vssd1 vccd1 vccd1 _15565_/Y sky130_fd_sc_hd__inv_2
X_12777_ _19245_/Q vssd1 vssd1 vccd1 vccd1 _12777_/Y sky130_fd_sc_hd__inv_2
XPHY_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17304_ _17303_/X _09857_/A _17518_/S vssd1 vssd1 vccd1 vccd1 _17304_/X sky130_fd_sc_hd__mux2_1
XPHY_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14516_ _18330_/Q _14504_/A _14474_/X _14505_/A vssd1 vssd1 vccd1 vccd1 _18330_/D
+ sky130_fd_sc_hd__a22o_1
X_18284_ _18435_/CLK _18284_/D vssd1 vssd1 vccd1 vccd1 _18284_/Q sky130_fd_sc_hd__dfxtp_1
X_11728_ _19507_/Q _11723_/X _16939_/X _11724_/X vssd1 vssd1 vccd1 vccd1 hold218/A
+ sky130_fd_sc_hd__a22o_1
X_15496_ _15535_/A _15496_/B vssd1 vssd1 vccd1 vccd1 _15496_/Y sky130_fd_sc_hd__nor2_1
XFILLER_230_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16743__B _16743_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17235_ _17234_/X _12917_/Y _17541_/S vssd1 vssd1 vccd1 vccd1 _17235_/X sky130_fd_sc_hd__mux2_1
XPHY_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14447_ _18372_/Q _14438_/A _14419_/X _14439_/A vssd1 vssd1 vccd1 vccd1 _18372_/D
+ sky130_fd_sc_hd__a22o_1
X_11659_ _11659_/A vssd1 vssd1 vccd1 vccd1 _19545_/D sky130_fd_sc_hd__inv_2
XANTENNA__18842__RESET_B repeater233/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17166_ _17165_/X _13540_/A _17536_/S vssd1 vssd1 vccd1 vccd1 _17166_/X sky130_fd_sc_hd__mux2_2
X_14378_ _19849_/Q _14378_/B _15318_/B vssd1 vssd1 vccd1 vccd1 _15058_/C sky130_fd_sc_hd__or3_4
XFILLER_127_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16117_ _20062_/Q _16204_/A vssd1 vssd1 vccd1 vccd1 _16117_/X sky130_fd_sc_hd__and2_1
X_13329_ _18846_/Q vssd1 vssd1 vccd1 vccd1 _13469_/A sky130_fd_sc_hd__inv_1
XANTENNA__09698__A2_N _19409_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17097_ _17096_/X _09700_/Y _17523_/S vssd1 vssd1 vccd1 vccd1 _17097_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12064__A _15774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16048_ _19027_/Q vssd1 vssd1 vccd1 vccd1 _16048_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17066__S _17474_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19807_ _19813_/CLK _19807_/D repeater224/X vssd1 vssd1 vccd1 vccd1 _19807_/Q sky130_fd_sc_hd__dfrtp_1
X_17999_ _18412_/CLK _17999_/D vssd1 vssd1 vccd1 vccd1 _17999_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12467__B1 _12344_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19738_ _20051_/CLK _19738_/D repeater206/X vssd1 vssd1 vccd1 vccd1 _19738_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__19630__RESET_B repeater257/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19669_ _19867_/CLK hold150/X repeater262/X vssd1 vssd1 vccd1 vccd1 _19669_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__14208__A1 _19119_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_225_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09422_ _19912_/Q _09381_/Y _19933_/Q _09418_/Y _09421_/X vssd1 vssd1 vccd1 vccd1
+ _09440_/A sky130_fd_sc_hd__o221a_1
XFILLER_241_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09353_ _20024_/Q vssd1 vssd1 vccd1 vccd1 _09484_/A sky130_fd_sc_hd__inv_2
X_09284_ _15749_/C _14245_/A _11742_/A _09340_/B vssd1 vssd1 vccd1 vccd1 _09293_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_193_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18583__RESET_B repeater274/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11745__A2 _11730_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17330__A0 _17486_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19789__RESET_B repeater203/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold287_A HWDATA[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08999_ _15890_/A _11936_/A vssd1 vssd1 vccd1 vccd1 _12187_/A sky130_fd_sc_hd__or2_4
XFILLER_87_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19371__RESET_B repeater241/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10961_ _10996_/A _10996_/B vssd1 vssd1 vccd1 vccd1 _10992_/A sky130_fd_sc_hd__or2_1
XFILLER_90_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12700_ _18966_/Q _12698_/X _12599_/X _12699_/X vssd1 vssd1 vccd1 vccd1 _18966_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_43_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13680_ hold335/X vssd1 vssd1 vccd1 vccd1 _13680_/X sky130_fd_sc_hd__buf_2
XFILLER_216_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10892_ _15826_/A _14245_/D vssd1 vssd1 vccd1 vccd1 _10894_/A sky130_fd_sc_hd__or2_2
XFILLER_203_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12631_ _19013_/Q _12629_/X _12401_/X _12630_/X vssd1 vssd1 vccd1 vccd1 _19013_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15350_ _15358_/A _17594_/X vssd1 vssd1 vccd1 vccd1 _18496_/D sky130_fd_sc_hd__and2_1
XFILLER_169_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12562_ _12600_/A vssd1 vssd1 vccd1 vccd1 _12577_/A sky130_fd_sc_hd__clkbuf_2
XPHY_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14301_ _15296_/B _14301_/B vssd1 vssd1 vccd1 vccd1 _14557_/C sky130_fd_sc_hd__or2_2
XPHY_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17795__S1 _19646_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11513_ _11476_/A _11476_/B _11506_/X _11511_/Y vssd1 vssd1 vccd1 vccd1 _19596_/D
+ sky130_fd_sc_hd__a211oi_2
XPHY_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11988__A _12309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15281_ _15205_/Y _15334_/B _15386_/A _10638_/Y _15277_/Y vssd1 vssd1 vccd1 vccd1
+ _15282_/A sky130_fd_sc_hd__o32a_1
XPHY_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10892__A _15826_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12493_ _19092_/Q _12489_/X _12375_/X _12492_/X vssd1 vssd1 vccd1 vccd1 _19092_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17020_ _17019_/X _09374_/Y _17413_/S vssd1 vssd1 vccd1 vccd1 _17020_/X sky130_fd_sc_hd__mux2_1
XPHY_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14232_ _18502_/Q _14232_/B vssd1 vssd1 vccd1 vccd1 _14233_/B sky130_fd_sc_hd__or2_1
XFILLER_8_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11444_ _19128_/Q vssd1 vssd1 vccd1 vccd1 _11444_/Y sky130_fd_sc_hd__inv_2
XFILLER_109_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_161_HCLK clkbuf_4_0_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19513_/CLK sky130_fd_sc_hd__clkbuf_16
X_14163_ _19115_/Q vssd1 vssd1 vccd1 vccd1 _16644_/A sky130_fd_sc_hd__inv_2
XANTENNA__17321__A0 _17486_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10944__A0 _19671_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11375_ _19569_/Q vssd1 vssd1 vccd1 vccd1 _11582_/A sky130_fd_sc_hd__inv_2
XFILLER_152_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13114_ _19188_/Q vssd1 vssd1 vccd1 vccd1 _13114_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10326_ _10361_/A _10361_/B vssd1 vssd1 vccd1 vccd1 _10357_/A sky130_fd_sc_hd__or2_1
XANTENNA__19754__CLK _19900_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14094_ _14094_/A _14094_/B _14080_/X _14093_/X vssd1 vssd1 vccd1 vccd1 _14116_/A
+ sky130_fd_sc_hd__or4bb_4
X_18971_ _19591_/CLK _18971_/D hold363/X vssd1 vssd1 vccd1 vccd1 _18971_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_106_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15195__A _15195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17922_ _18329_/Q _18009_/Q _18313_/Q _18305_/Q _17923_/S0 _19646_/Q vssd1 vssd1
+ vccd1 vccd1 _17922_/X sky130_fd_sc_hd__mux4_2
XFILLER_59_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13045_ _18901_/Q vssd1 vssd1 vccd1 vccd1 _13073_/A sky130_fd_sc_hd__inv_2
XANTENNA__13708__A _18761_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10257_ _14300_/A vssd1 vssd1 vccd1 vccd1 _11027_/B sky130_fd_sc_hd__inv_2
XANTENNA__12697__B1 _12596_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_repeater207_A repeater208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12612__A _12650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19459__RESET_B repeater272/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17853_ _16340_/Y _16341_/Y _16342_/Y _16343_/Y _17913_/S0 _19632_/Q vssd1 vssd1
+ vccd1 vccd1 _17853_/X sky130_fd_sc_hd__mux4_2
X_10188_ _10147_/X _19874_/Q _10188_/S vssd1 vssd1 vccd1 vccd1 _19874_/D sky130_fd_sc_hd__mux2_1
XFILLER_120_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17614__S _17614_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16804_ _17486_/A0 _13101_/Y _17543_/S vssd1 vssd1 vccd1 vccd1 _16804_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12449__B1 _12386_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17784_ _17780_/X _17781_/X _17782_/X _17783_/X _19647_/Q _19648_/Q vssd1 vssd1 vccd1
+ vccd1 _17784_/X sky130_fd_sc_hd__mux4_2
X_14996_ _18958_/Q vssd1 vssd1 vccd1 vccd1 _14996_/X sky130_fd_sc_hd__buf_2
XFILLER_208_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_140_HCLK_A clkbuf_4_3_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19523_ _20049_/CLK _19523_/D repeater190/X vssd1 vssd1 vccd1 vccd1 _19523_/Q sky130_fd_sc_hd__dfstp_1
X_16735_ _16682_/X _16735_/B _16735_/C vssd1 vssd1 vccd1 vccd1 _16735_/Y sky130_fd_sc_hd__nand3b_4
X_13947_ _13947_/A _13947_/B vssd1 vssd1 vccd1 vccd1 _13957_/A sky130_fd_sc_hd__or2_1
XFILLER_35_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16666_ _16666_/A _16668_/B vssd1 vssd1 vccd1 vccd1 _16666_/Y sky130_fd_sc_hd__nor2_1
X_19454_ _19462_/CLK _19454_/D repeater272/X vssd1 vssd1 vccd1 vccd1 _19454_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_179_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13878_ _19210_/Q vssd1 vssd1 vccd1 vccd1 _13878_/Y sky130_fd_sc_hd__inv_2
X_15617_ _15617_/A vssd1 vssd1 vccd1 vccd1 _15622_/B sky130_fd_sc_hd__inv_2
X_18405_ _18959_/CLK _18405_/D vssd1 vssd1 vccd1 vccd1 _18405_/Q sky130_fd_sc_hd__dfxtp_1
X_12829_ _18835_/Q vssd1 vssd1 vccd1 vccd1 _12829_/Y sky130_fd_sc_hd__inv_2
X_19385_ _19927_/CLK _19385_/D repeater234/X vssd1 vssd1 vccd1 vccd1 _19385_/Q sky130_fd_sc_hd__dfrtp_1
X_16597_ _16597_/A vssd1 vssd1 vccd1 vccd1 _16597_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_188_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15548_ _15552_/B _15547_/X _15512_/X vssd1 vssd1 vccd1 vccd1 _15548_/X sky130_fd_sc_hd__o21a_1
X_18336_ _19849_/CLK _18336_/D vssd1 vssd1 vccd1 vccd1 _18336_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12621__B1 _12386_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16473__B _17517_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17786__S1 _19646_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18267_ _18268_/CLK _18267_/D vssd1 vssd1 vccd1 vccd1 _18267_/Q sky130_fd_sc_hd__dfxtp_1
X_15479_ _15479_/A _15479_/B vssd1 vssd1 vccd1 vccd1 _15479_/Y sky130_fd_sc_hd__nor2_1
XFILLER_147_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14374__B1 _14326_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17218_ _17217_/X _13069_/B _17542_/S vssd1 vssd1 vccd1 vccd1 _17218_/X sky130_fd_sc_hd__mux2_1
X_18198_ _18198_/CLK _18198_/D vssd1 vssd1 vccd1 vccd1 _18198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17149_ _17148_/X _09859_/A _17414_/S vssd1 vssd1 vccd1 vccd1 _17149_/X sky130_fd_sc_hd__mux2_1
X_09971_ _09867_/A _09867_/B _09967_/Y _09970_/X vssd1 vssd1 vccd1 vccd1 _19959_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_226_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08922_ _18785_/Q vssd1 vssd1 vccd1 vccd1 _08922_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13618__A _15195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20091_ _20091_/CLK _20091_/D repeater234/X vssd1 vssd1 vccd1 vccd1 _20091_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__19811__RESET_B repeater222/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12688__B1 _12028_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19129__RESET_B repeater274/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_245_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17524__S _17524_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_42_HCLK clkbuf_opt_2_HCLK/A vssd1 vssd1 vccd1 vccd1 _19812_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_37_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_241_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_62_HCLK_A clkbuf_opt_3_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_225_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09405_ _19925_/Q _09401_/Y _10041_/A _19385_/Q _09404_/X vssd1 vssd1 vccd1 vccd1
+ _09417_/C sky130_fd_sc_hd__o221a_1
XFILLER_52_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18764__RESET_B repeater196/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_241_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09336_ _10791_/A _15727_/B vssd1 vssd1 vccd1 vccd1 _10786_/B sky130_fd_sc_hd__and2_1
XFILLER_187_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17777__S1 _19646_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09267_ _19499_/Q _15749_/A _11842_/B vssd1 vssd1 vccd1 vccd1 _12436_/C sky130_fd_sc_hd__or3_4
XFILLER_194_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14365__B1 _14314_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19777__CLK _19780_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09198_ _09198_/A _09205_/B vssd1 vssd1 vccd1 vccd1 _09198_/X sky130_fd_sc_hd__or2_1
XFILLER_106_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11160_ _19615_/Q _11160_/B vssd1 vssd1 vccd1 vccd1 _11161_/B sky130_fd_sc_hd__or2_1
XFILLER_122_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10111_ _18557_/Q _18556_/Q vssd1 vssd1 vccd1 vccd1 _15453_/A sky130_fd_sc_hd__or2_2
X_11091_ _11106_/A vssd1 vssd1 vccd1 vccd1 _11091_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__12679__B1 hold315/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19552__RESET_B hold348/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10042_ _10042_/A _10042_/B vssd1 vssd1 vccd1 vccd1 _10065_/A sky130_fd_sc_hd__or2_1
XFILLER_248_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17434__S _17564_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14850_ _18143_/Q _14845_/X _14808_/X _14847_/X vssd1 vssd1 vccd1 vccd1 _18143_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_29_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13801_ _18705_/Q vssd1 vssd1 vccd1 vccd1 _13964_/C sky130_fd_sc_hd__inv_2
XFILLER_91_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input18_A HADDR[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14781_ _18179_/Q _14772_/A _14780_/X _14773_/A vssd1 vssd1 vccd1 vccd1 _18179_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18476__D _18476_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11993_ _11991_/X _19364_/Q _11993_/S vssd1 vssd1 vccd1 vccd1 _19364_/D sky130_fd_sc_hd__mux2_1
X_16520_ _17275_/X _15904_/X _17287_/X _16509_/X vssd1 vssd1 vccd1 vccd1 _16520_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_205_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13732_ _13733_/A _13293_/X _13731_/X vssd1 vssd1 vccd1 vccd1 _18755_/D sky130_fd_sc_hd__o21ba_1
X_10944_ _19671_/Q _10943_/X _17751_/X vssd1 vssd1 vccd1 vccd1 _19671_/D sky130_fd_sc_hd__mux2_1
XFILLER_17_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16451_ _16449_/Y _15867_/B _16450_/Y _16049_/X vssd1 vssd1 vccd1 vccd1 _16451_/X
+ sky130_fd_sc_hd__o22a_1
X_13663_ _18783_/Q _13656_/X hold239/X _13658_/X vssd1 vssd1 vccd1 vccd1 _18783_/D
+ sky130_fd_sc_hd__a22o_1
X_10875_ _10878_/A vssd1 vssd1 vccd1 vccd1 _10875_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_43_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16593__A1 _17252_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16574__A _16684_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_231_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15402_ _15402_/A _17579_/X vssd1 vssd1 vccd1 vccd1 _18533_/D sky130_fd_sc_hd__and2_1
XPHY_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12614_ _12650_/A vssd1 vssd1 vccd1 vccd1 _12651_/A sky130_fd_sc_hd__inv_2
X_19170_ _19208_/CLK _19170_/D hold370/X vssd1 vssd1 vccd1 vccd1 _19170_/Q sky130_fd_sc_hd__dfrtp_2
X_16382_ _18521_/Q vssd1 vssd1 vccd1 vccd1 _16382_/Y sky130_fd_sc_hd__inv_2
XPHY_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12603__B1 _12602_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13594_ _13594_/A vssd1 vssd1 vccd1 vccd1 _13597_/B sky130_fd_sc_hd__inv_2
XFILLER_185_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18121_ _18145_/CLK _18121_/D vssd1 vssd1 vccd1 vccd1 _18121_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15333_ _15333_/A _15850_/A vssd1 vssd1 vccd1 vccd1 _18514_/D sky130_fd_sc_hd__nor2_1
XANTENNA__17768__S1 _19646_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12545_ _12545_/A vssd1 vssd1 vccd1 vccd1 _12545_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_repeater157_A _17459_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10090__B1 _10079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18052_ _19851_/CLK _18052_/D vssd1 vssd1 vccd1 vccd1 _18052_/Q sky130_fd_sc_hd__dfxtp_1
X_15264_ _19780_/Q _18551_/Q _15256_/A _15304_/A _15259_/B vssd1 vssd1 vccd1 vccd1
+ _15264_/X sky130_fd_sc_hd__o32a_1
X_12476_ _19101_/Q _12471_/X _12225_/X _12472_/X vssd1 vssd1 vccd1 vccd1 _19101_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_177_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17003_ _17473_/A0 _16609_/Y _17547_/S vssd1 vssd1 vccd1 vccd1 _17003_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14215_ _19117_/Q vssd1 vssd1 vccd1 vccd1 _16666_/A sky130_fd_sc_hd__inv_2
XFILLER_144_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11427_ _19572_/Q _11423_/Y _11620_/A _19130_/Q _11426_/X vssd1 vssd1 vccd1 vccd1
+ _11433_/C sky130_fd_sc_hd__o221a_1
X_15195_ _15195_/A _15195_/B vssd1 vssd1 vccd1 vccd1 _15195_/Y sky130_fd_sc_hd__nor2_1
XFILLER_6_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output86_A _16581_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14146_ _18675_/Q _14145_/Y _14112_/A _14146_/C1 vssd1 vssd1 vccd1 vccd1 _18675_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_141_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11358_ _18991_/Q vssd1 vssd1 vccd1 vccd1 _11358_/Y sky130_fd_sc_hd__inv_2
XFILLER_193_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10309_ _15640_/B _10309_/B vssd1 vssd1 vccd1 vccd1 _15678_/B sky130_fd_sc_hd__or2_1
X_14077_ _19076_/Q vssd1 vssd1 vccd1 vccd1 _14077_/Y sky130_fd_sc_hd__inv_2
X_18954_ _18954_/CLK _18954_/D repeater257/X vssd1 vssd1 vccd1 vccd1 _18954_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_113_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11289_ _19600_/Q vssd1 vssd1 vccd1 vccd1 _11480_/A sky130_fd_sc_hd__inv_2
XFILLER_79_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17905_ _15802_/Y _15803_/Y _15804_/Y _15805_/Y _17908_/S0 _18759_/Q vssd1 vssd1
+ vccd1 vccd1 _17905_/X sky130_fd_sc_hd__mux4_2
X_13028_ _13021_/A _13021_/B _18919_/Q _12969_/D _12962_/X vssd1 vssd1 vccd1 vccd1
+ _18919_/D sky130_fd_sc_hd__o221a_1
Xclkbuf_leaf_65_HCLK clkbuf_opt_4_HCLK/A vssd1 vssd1 vccd1 vccd1 _20122_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_79_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18885_ _18886_/CLK _18885_/D repeater220/X vssd1 vssd1 vccd1 vccd1 _18885_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_66_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17344__S _17568_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11893__A1 _19422_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17836_ _16421_/Y _16422_/Y _16423_/Y _16424_/Y _17908_/S0 _18759_/Q vssd1 vssd1
+ vccd1 vccd1 _17836_/X sky130_fd_sc_hd__mux4_2
XFILLER_227_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16468__B _16469_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrebuffer17 _13071_/B vssd1 vssd1 vccd1 vccd1 _13195_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_26_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17767_ _18322_/Q _18002_/Q _18306_/Q _18298_/Q _17923_/S0 _19646_/Q vssd1 vssd1
+ vccd1 vccd1 _17767_/X sky130_fd_sc_hd__mux4_2
Xrebuffer28 _14011_/B vssd1 vssd1 vccd1 vccd1 _14140_/C1 sky130_fd_sc_hd__dlygate4sd1_1
X_14979_ _14979_/A vssd1 vssd1 vccd1 vccd1 _14979_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_81_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrebuffer39 _19286_/Q vssd1 vssd1 vccd1 vccd1 _17055_/A1 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_19_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19506_ _19506_/CLK hold228/X repeater256/X vssd1 vssd1 vccd1 vccd1 _19506_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_235_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16718_ _16718_/A _16718_/B vssd1 vssd1 vccd1 vccd1 _16718_/Y sky130_fd_sc_hd__nor2_1
XFILLER_212_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17698_ _19820_/Q _19762_/Q _18548_/Q vssd1 vssd1 vccd1 vccd1 _17698_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19437_ _19437_/CLK _19437_/D repeater269/X vssd1 vssd1 vccd1 vccd1 _19437_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_90_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16649_ _16649_/A _16668_/B vssd1 vssd1 vccd1 vccd1 _16649_/Y sky130_fd_sc_hd__nor2_1
XFILLER_34_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_4_13_0_HCLK_A clkbuf_3_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14595__B1 _14582_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19368_ _19971_/CLK _19368_/D repeater241/X vssd1 vssd1 vccd1 vccd1 _19368_/Q sky130_fd_sc_hd__dfrtp_1
X_09121_ _20083_/Q vssd1 vssd1 vccd1 vccd1 _09154_/A sky130_fd_sc_hd__inv_2
X_18319_ _18431_/CLK _18319_/D vssd1 vssd1 vccd1 vccd1 _18319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrebuffer107 _13079_/B vssd1 vssd1 vccd1 vccd1 _13185_/C1 sky130_fd_sc_hd__dlygate4sd1_1
X_19299_ _20013_/CLK _19299_/D repeater241/X vssd1 vssd1 vccd1 vccd1 _19299_/Q sky130_fd_sc_hd__dfrtp_1
Xrebuffer118 _11472_/B vssd1 vssd1 vccd1 vccd1 _11522_/C1 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_176_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09052_ _20108_/Q _09041_/X _09051_/X _09043_/X vssd1 vssd1 vccd1 vccd1 _20108_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_108_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17519__S _17537_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20007__CLK _20013_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09954_ _09954_/A vssd1 vssd1 vccd1 vccd1 _09954_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20074_ _20076_/CLK _20074_/D repeater196/X vssd1 vssd1 vccd1 vccd1 _20074_/Q sky130_fd_sc_hd__dfrtp_4
X_09885_ _19958_/Q _09884_/Y _09861_/A _19345_/Q vssd1 vssd1 vccd1 vccd1 _09885_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_85_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17254__S _17513_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold152_A HSEL vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16394__A _16633_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16575__B2 _15898_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13389__A1 _20101_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10660_ _10660_/A _18508_/D vssd1 vssd1 vccd1 vccd1 _10676_/A sky130_fd_sc_hd__or2_4
XFILLER_201_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09319_ _15721_/A _09317_/X _18656_/Q _09318_/Y vssd1 vssd1 vccd1 vccd1 _15723_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_178_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16327__A1 _15846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10591_ _10593_/B _19799_/Q _19800_/Q vssd1 vssd1 vccd1 vccd1 _10594_/A sky130_fd_sc_hd__nor3b_2
XFILLER_21_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16327__B2 _16319_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12330_ _19183_/Q _12327_/X _12086_/X _12328_/X vssd1 vssd1 vccd1 vccd1 _19183_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_127_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17429__S _17564_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12261_ _12298_/A vssd1 vssd1 vccd1 vccd1 _12300_/A sky130_fd_sc_hd__inv_2
XANTENNA__19733__RESET_B repeater208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14000_ _18674_/Q vssd1 vssd1 vccd1 vccd1 _14005_/A sky130_fd_sc_hd__inv_2
X_11212_ _19601_/Q vssd1 vssd1 vccd1 vccd1 _11481_/A sky130_fd_sc_hd__inv_2
XFILLER_107_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12192_ _12206_/A vssd1 vssd1 vccd1 vccd1 _12192_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_88_HCLK clkbuf_4_12_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20035_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__17922__S1 _19646_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11143_ _19628_/Q vssd1 vssd1 vccd1 vccd1 _11144_/A sky130_fd_sc_hd__inv_2
Xoutput86 _16581_/Y vssd1 vssd1 vccd1 vccd1 HRDATA[16] sky130_fd_sc_hd__clkbuf_2
Xoutput97 _16698_/Y vssd1 vssd1 vccd1 vccd1 HRDATA[26] sky130_fd_sc_hd__clkbuf_2
XANTENNA__14510__B1 _14509_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11074_ _19849_/Q _14489_/B _14476_/A vssd1 vssd1 vccd1 vccd1 _11074_/Y sky130_fd_sc_hd__o21ai_1
X_15951_ _17978_/Q vssd1 vssd1 vccd1 vccd1 _15951_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17164__S _17534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10025_ _10025_/A vssd1 vssd1 vccd1 vccd1 _10026_/A sky130_fd_sc_hd__clkbuf_2
X_14902_ _18110_/Q _14896_/X _14707_/X _14898_/X vssd1 vssd1 vccd1 vccd1 _18110_/D
+ sky130_fd_sc_hd__a22o_1
X_18670_ _19812_/CLK _18670_/D repeater222/X vssd1 vssd1 vccd1 vccd1 _18670_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_76_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15882_ _17558_/X vssd1 vssd1 vccd1 vccd1 _15882_/Y sky130_fd_sc_hd__inv_2
XFILLER_237_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17621_ _20051_/Q _19725_/Q _17621_/S vssd1 vssd1 vccd1 vccd1 _17621_/X sky130_fd_sc_hd__mux2_1
X_14833_ _14833_/A vssd1 vssd1 vccd1 vccd1 _14834_/A sky130_fd_sc_hd__inv_2
XANTENNA_output124_A _15775_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18686__RESET_B hold359/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_245_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14764_ _18191_/Q _14759_/X _14751_/X _14761_/X vssd1 vssd1 vccd1 vccd1 _18191_/D
+ sky130_fd_sc_hd__a22o_1
X_17552_ _17551_/X _20040_/Q _19498_/Q vssd1 vssd1 vccd1 vccd1 _17552_/X sky130_fd_sc_hd__mux2_1
X_11976_ _19373_/Q _11969_/X _11975_/X _11970_/X vssd1 vssd1 vccd1 vccd1 _19373_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10410__A _10410_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18615__RESET_B repeater267/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19942__CLK _20013_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16503_ _19035_/Q vssd1 vssd1 vccd1 vccd1 _16503_/Y sky130_fd_sc_hd__inv_2
X_13715_ _17762_/X vssd1 vssd1 vccd1 vccd1 _13715_/Y sky130_fd_sc_hd__inv_2
XFILLER_205_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17483_ _15963_/X _12827_/Y _17534_/S vssd1 vssd1 vccd1 vccd1 _17483_/X sky130_fd_sc_hd__mux2_1
X_10927_ _17723_/X _10923_/X _19678_/Q _10924_/X vssd1 vssd1 vccd1 vccd1 _19678_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_60_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14695_ _14695_/A vssd1 vssd1 vccd1 vccd1 _15145_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA_repeater274_A hold348/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16566__B2 _16003_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19222_ _19222_/CLK _19222_/D repeater186/X vssd1 vssd1 vccd1 vccd1 _19222_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_31_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13646_ _13646_/A vssd1 vssd1 vccd1 vccd1 _13646_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16434_ _17313_/X _16434_/B vssd1 vssd1 vccd1 vccd1 _16434_/X sky130_fd_sc_hd__and2_1
X_10858_ _19708_/Q _10855_/X _10446_/X _10857_/X vssd1 vssd1 vccd1 vccd1 _19708_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19153_ _19576_/CLK _19153_/D repeater268/X vssd1 vssd1 vccd1 vccd1 _19153_/Q sky130_fd_sc_hd__dfrtp_4
X_16365_ _17342_/X _16435_/B vssd1 vssd1 vccd1 vccd1 _16365_/Y sky130_fd_sc_hd__nand2_1
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13577_ _13577_/A vssd1 vssd1 vccd1 vccd1 _13577_/Y sky130_fd_sc_hd__inv_2
XFILLER_158_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10789_ _10805_/A _19739_/Q vssd1 vssd1 vccd1 vccd1 _10789_/Y sky130_fd_sc_hd__nor2_1
XFILLER_9_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15316_ _15315_/Y _15307_/X _15242_/Y _15245_/X vssd1 vssd1 vccd1 vccd1 _15316_/X
+ sky130_fd_sc_hd__o22a_1
X_18104_ _18137_/CLK _18104_/D vssd1 vssd1 vccd1 vccd1 _18104_/Q sky130_fd_sc_hd__dfxtp_1
X_12528_ _12528_/A vssd1 vssd1 vccd1 vccd1 _12528_/X sky130_fd_sc_hd__clkbuf_2
X_19084_ _19119_/CLK _19084_/D hold351/X vssd1 vssd1 vccd1 vccd1 _19084_/Q sky130_fd_sc_hd__dfrtp_2
X_16296_ _17374_/X _16415_/B vssd1 vssd1 vccd1 vccd1 _16296_/Y sky130_fd_sc_hd__nand2_1
X_15247_ _15389_/B _15285_/A _15436_/A _15246_/Y vssd1 vssd1 vccd1 vccd1 _18631_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_8_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18035_ _19851_/CLK _18035_/D vssd1 vssd1 vccd1 vccd1 _18035_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17339__S _19498_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12459_ _19114_/Q _12457_/X _12401_/X _12458_/X vssd1 vssd1 vccd1 vccd1 _19114_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_126_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15178_ _17939_/Q _15171_/A _10423_/A _15172_/A vssd1 vssd1 vccd1 vccd1 _17939_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_153_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14129_ _14129_/A vssd1 vssd1 vccd1 vccd1 _14129_/Y sky130_fd_sc_hd__clkinv_1
XANTENNA__17913__S1 _19632_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19986_ _19992_/CLK _19986_/D repeater193/X vssd1 vssd1 vccd1 vccd1 _19986_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_98_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18937_ _19325_/CLK _18937_/D repeater215/X vssd1 vssd1 vccd1 vccd1 _18937_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_239_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17074__S _17386_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09670_ _20003_/Q vssd1 vssd1 vccd1 vccd1 _09670_/Y sky130_fd_sc_hd__inv_2
X_18868_ _20122_/CLK _18868_/D repeater217/X vssd1 vssd1 vccd1 vccd1 _18868_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_95_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17819_ _17815_/X _17816_/X _17817_/X _17818_/X _18751_/Q _18752_/Q vssd1 vssd1 vccd1
+ vccd1 _17819_/X sky130_fd_sc_hd__mux4_2
XFILLER_54_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16629__D _16629_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18799_ _19435_/CLK _18799_/D repeater258/X vssd1 vssd1 vccd1 vccd1 _18799_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_235_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14568__B1 _14567_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09104_ _14780_/A vssd1 vssd1 vccd1 vccd1 _12238_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_175_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09035_ hold306/X vssd1 vssd1 vccd1 vccd1 hold305/A sky130_fd_sc_hd__buf_4
XANTENNA__17249__S _17541_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09556__A _19319_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold330 hold330/A vssd1 vssd1 vccd1 vccd1 hold330/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold341 input71/X vssd1 vssd1 vccd1 vccd1 hold341/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold352 input34/X vssd1 vssd1 vccd1 vccd1 hold352/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17904__S1 _19634_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold363 hold363/A vssd1 vssd1 vccd1 vccd1 hold363/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20049__RESET_B repeater208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09937_ _09868_/A _19352_/Q _09857_/B _19340_/Q _09936_/X vssd1 vssd1 vccd1 vccd1
+ _09947_/B sky130_fd_sc_hd__o221a_1
XFILLER_131_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20057_ _20057_/CLK _20057_/D repeater204/X vssd1 vssd1 vccd1 vccd1 _20057_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_218_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09868_ _09868_/A _09967_/A vssd1 vssd1 vccd1 vccd1 _09869_/B sky130_fd_sc_hd__or2_2
XFILLER_219_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09799_ _09792_/A _09792_/B _09797_/Y _09813_/C vssd1 vssd1 vccd1 vccd1 _19980_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_234_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater180 _17530_/S vssd1 vssd1 vccd1 vccd1 _17414_/S sky130_fd_sc_hd__buf_8
XPHY_4312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17712__S _18546_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater191 repeater210/X vssd1 vssd1 vccd1 vccd1 repeater191/X sky130_fd_sc_hd__buf_8
XPHY_4323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11830_ _11830_/A _11830_/B _13279_/C vssd1 vssd1 vccd1 vccd1 _16234_/A sky130_fd_sc_hd__or3_4
XPHY_4334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10230__A _19832_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09278__A2 _09270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11761_ hold174/X _11757_/X _19483_/Q _11758_/X vssd1 vssd1 vccd1 vccd1 hold176/A
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12282__A1 _19210_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13500_ _18760_/Q vssd1 vssd1 vccd1 vccd1 _13500_/Y sky130_fd_sc_hd__inv_2
XPHY_3666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10712_ hold322/X vssd1 vssd1 vccd1 vccd1 _10712_/Y sky130_fd_sc_hd__inv_2
XPHY_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10832__A2 _10831_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17840__S0 _17913_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14480_ _14480_/A vssd1 vssd1 vccd1 vccd1 _14480_/X sky130_fd_sc_hd__clkbuf_2
XPHY_3688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11692_ _11692_/A vssd1 vssd1 vccd1 vccd1 _11692_/X sky130_fd_sc_hd__clkbuf_2
XPHY_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19985__RESET_B repeater193/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13431_ _13431_/A _13431_/B _13431_/C _13431_/D vssd1 vssd1 vccd1 vccd1 _13433_/C
+ sky130_fd_sc_hd__or4_4
XFILLER_42_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10643_ _19783_/Q _10643_/B vssd1 vssd1 vccd1 vccd1 _10644_/B sky130_fd_sc_hd__or2_1
XPHY_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11061__A _19633_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16150_ _15749_/B _16143_/X _16145_/X _16147_/X _16149_/X vssd1 vssd1 vccd1 vccd1
+ _16150_/X sky130_fd_sc_hd__o2111a_1
X_13362_ _20116_/Q vssd1 vssd1 vccd1 vccd1 _13362_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10574_ _10574_/A _19807_/Q _19808_/Q vssd1 vssd1 vccd1 vccd1 _10574_/X sky130_fd_sc_hd__or3b_1
XFILLER_167_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15101_ _17990_/Q _15095_/X _14810_/A _15097_/X vssd1 vssd1 vccd1 vccd1 _17990_/D
+ sky130_fd_sc_hd__a22o_1
Xrebuffer8 _13077_/B vssd1 vssd1 vccd1 vccd1 _13186_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_139_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17159__S _17534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11996__A _11996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12313_ _12313_/A vssd1 vssd1 vccd1 vccd1 _12313_/X sky130_fd_sc_hd__buf_4
X_16081_ _18117_/Q vssd1 vssd1 vccd1 vccd1 _16081_/Y sky130_fd_sc_hd__inv_2
XFILLER_155_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13293_ _13729_/A _13293_/B vssd1 vssd1 vccd1 vccd1 _13293_/X sky130_fd_sc_hd__or2_2
X_15032_ _18035_/Q _15024_/A _15006_/X _15025_/A vssd1 vssd1 vccd1 vccd1 _18035_/D
+ sky130_fd_sc_hd__a22o_1
X_12244_ _19226_/Q _15232_/B vssd1 vssd1 vccd1 vccd1 _12247_/A sky130_fd_sc_hd__nor2_1
XANTENNA__16998__S _17385_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19840_ _19846_/CLK _19840_/D repeater272/X vssd1 vssd1 vccd1 vccd1 _19840_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_107_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12175_ _19266_/Q _12171_/X _11918_/X _12172_/X vssd1 vssd1 vccd1 vccd1 _19266_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_3_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11126_ _17747_/X _11066_/B _11061_/X vssd1 vssd1 vccd1 vccd1 _11127_/B sky130_fd_sc_hd__a21oi_1
X_19771_ _19771_/CLK _19771_/D repeater228/X vssd1 vssd1 vccd1 vccd1 _19771_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_95_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16983_ _17819_/X _19901_/Q _16986_/S vssd1 vssd1 vccd1 vccd1 _16983_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13298__B1 _18752_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18722_ _19224_/CLK _18722_/D repeater253/X vssd1 vssd1 vccd1 vccd1 _18722_/Q sky130_fd_sc_hd__dfrtp_1
X_11057_ _19642_/Q _11056_/Y _11049_/A vssd1 vssd1 vccd1 vccd1 _19642_/D sky130_fd_sc_hd__o21a_1
X_15934_ _18043_/Q vssd1 vssd1 vccd1 vccd1 _15934_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10008_ _19932_/Q vssd1 vssd1 vccd1 vccd1 _10047_/C sky130_fd_sc_hd__inv_2
X_18653_ _20050_/CLK _18653_/D repeater206/X vssd1 vssd1 vccd1 vccd1 _18653_/Q sky130_fd_sc_hd__dfrtp_2
X_15865_ _18736_/Q vssd1 vssd1 vccd1 vccd1 _15865_/Y sky130_fd_sc_hd__inv_2
X_17604_ _15319_/X _15319_/A _17605_/S vssd1 vssd1 vccd1 vccd1 _17604_/X sky130_fd_sc_hd__mux2_1
X_14816_ _14816_/A vssd1 vssd1 vccd1 vccd1 _14816_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_91_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14798__B1 _14782_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18584_ _19470_/CLK _18584_/D repeater274/X vssd1 vssd1 vccd1 vccd1 _18584_/Q sky130_fd_sc_hd__dfrtp_4
X_15796_ _18466_/Q vssd1 vssd1 vccd1 vccd1 _15796_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17535_ _17534_/X _13365_/Y _17535_/S vssd1 vssd1 vccd1 vccd1 _17535_/X sky130_fd_sc_hd__mux2_1
X_11959_ _19385_/Q _11955_/X hold317/X _11956_/X vssd1 vssd1 vccd1 vccd1 _19385_/D
+ sky130_fd_sc_hd__a22o_1
X_14747_ _14747_/A vssd1 vssd1 vccd1 vccd1 _14747_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__14547__A _14547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_199_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17831__S0 _17918_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17466_ _17465_/X _13491_/Y _17567_/S vssd1 vssd1 vccd1 vccd1 _17466_/X sky130_fd_sc_hd__mux2_1
X_14678_ _18235_/Q _14670_/A _09185_/X _14671_/A vssd1 vssd1 vccd1 vccd1 _18235_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_149_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19205_ _19208_/CLK _19205_/D hold367/X vssd1 vssd1 vccd1 vccd1 _19205_/Q sky130_fd_sc_hd__dfrtp_1
X_16417_ _18129_/Q vssd1 vssd1 vccd1 vccd1 _16417_/Y sky130_fd_sc_hd__inv_2
X_13629_ _11861_/B _15233_/A _17614_/S _12058_/B vssd1 vssd1 vccd1 vccd1 _13630_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_177_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12067__A _12121_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17397_ _17396_/X _08959_/Y _17566_/S vssd1 vssd1 vccd1 vccd1 _17397_/X sky130_fd_sc_hd__mux2_1
X_19136_ _19137_/CLK _19136_/D hold348/X vssd1 vssd1 vccd1 vccd1 _19136_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_192_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16348_ _18096_/Q vssd1 vssd1 vccd1 vccd1 _16348_/Y sky130_fd_sc_hd__inv_2
XFILLER_146_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16481__B _16481_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17069__S _17413_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19067_ _19585_/CLK _19067_/D hold363/X vssd1 vssd1 vccd1 vccd1 _19067_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_118_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16279_ _18271_/Q vssd1 vssd1 vccd1 vccd1 _16279_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16711__A1 _16798_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16711__B2 _16512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18018_ _18142_/CLK _18018_/D vssd1 vssd1 vccd1 vccd1 _18018_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14722__B1 _14606_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_218_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17898__S0 _17908_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18862__CLK _18866_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19988__CLK _19992_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19969_ _19970_/CLK _19969_/D repeater274/X vssd1 vssd1 vccd1 vccd1 _19969_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_234_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09722_ _09745_/A _09722_/A2 _09749_/A _19422_/Q _09721_/X vssd1 vssd1 vccd1 vccd1
+ _09727_/C sky130_fd_sc_hd__o221a_1
XFILLER_234_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09653_ _19984_/Q vssd1 vssd1 vccd1 vccd1 _09740_/A sky130_fd_sc_hd__inv_2
XFILLER_28_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17532__S _17548_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14789__B1 _14749_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09584_ _09584_/A vssd1 vssd1 vccd1 vccd1 _09584_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16656__B _16656_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18242__CLK _19847_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17822__S0 _17918_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_117_HCLK_A clkbuf_opt_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09018_ _09087_/A vssd1 vssd1 vccd1 vccd1 _09043_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_88_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10290_ _19869_/Q _10290_/B vssd1 vssd1 vccd1 vccd1 _10291_/B sky130_fd_sc_hd__nand2_1
XFILLER_151_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09196__A1 _18870_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17707__S _18546_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold160 HADDR[16] vssd1 vssd1 vccd1 vccd1 input8/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09196__B2 _17605_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold171 input11/X vssd1 vssd1 vccd1 vccd1 hold171/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17889__S0 _18760_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold182 hold182/A vssd1 vssd1 vccd1 vccd1 hold182/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 input1/X vssd1 vssd1 vccd1 vccd1 hold193/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15735__B _15735_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10750__A1 _19757_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20109_ _20122_/CLK _20109_/D repeater217/X vssd1 vssd1 vccd1 vccd1 _20109_/Q sky130_fd_sc_hd__dfrtp_4
X_13980_ _18694_/Q vssd1 vssd1 vccd1 vccd1 _14024_/A sky130_fd_sc_hd__inv_2
XANTENNA__12440__A _12478_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09499__A2 _19325_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_118_HCLK clkbuf_opt_0_HCLK/A vssd1 vssd1 vccd1 vccd1 _19610_/CLK sky130_fd_sc_hd__clkbuf_16
X_12931_ _19272_/Q _13008_/A _19284_/Q _12967_/B vssd1 vssd1 vccd1 vccd1 _12931_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_18_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17442__S _17518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15650_ _15654_/B vssd1 vssd1 vccd1 vccd1 _15657_/B sky130_fd_sc_hd__inv_2
X_12862_ _18924_/Q vssd1 vssd1 vccd1 vccd1 _13003_/A sky130_fd_sc_hd__inv_2
XPHY_4120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14601_ _14601_/A vssd1 vssd1 vccd1 vccd1 _14602_/A sky130_fd_sc_hd__inv_2
X_11813_ _19451_/Q _11807_/X _09067_/X _11808_/X vssd1 vssd1 vccd1 vccd1 _19451_/D
+ sky130_fd_sc_hd__a22o_1
X_15581_ _15581_/A _15581_/B vssd1 vssd1 vccd1 vccd1 _15581_/X sky130_fd_sc_hd__or2_1
XPHY_4164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12793_ _19239_/Q vssd1 vssd1 vccd1 vccd1 _12793_/Y sky130_fd_sc_hd__inv_2
XPHY_4175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14367__A _14368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14532_ _14532_/A vssd1 vssd1 vccd1 vccd1 _14533_/A sky130_fd_sc_hd__inv_2
X_17320_ _17319_/X _15471_/A _17524_/S vssd1 vssd1 vccd1 vccd1 _17320_/X sky130_fd_sc_hd__mux2_1
XPHY_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11744_ _19496_/Q _11737_/X _16928_/X _11738_/X vssd1 vssd1 vccd1 vccd1 hold253/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_53_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17813__S0 _17918_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17251_ _16587_/Y _19383_/Q _17529_/S vssd1 vssd1 vccd1 vccd1 _17251_/X sky130_fd_sc_hd__mux2_1
X_14463_ _14464_/A vssd1 vssd1 vccd1 vccd1 _14463_/X sky130_fd_sc_hd__clkbuf_2
XPHY_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11675_ _11675_/A vssd1 vssd1 vccd1 vccd1 _11675_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_14_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13414_ _20114_/Q vssd1 vssd1 vccd1 vccd1 _13414_/Y sky130_fd_sc_hd__inv_2
XFILLER_186_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16202_ _17965_/Q vssd1 vssd1 vccd1 vccd1 _16202_/Y sky130_fd_sc_hd__inv_2
XPHY_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10626_ _10625_/Y _10598_/A _10617_/X _10581_/A _10618_/A vssd1 vssd1 vccd1 vccd1
+ _10627_/A sky130_fd_sc_hd__o32a_1
X_17182_ _15768_/Y _14203_/Y _17546_/S vssd1 vssd1 vccd1 vccd1 _17182_/X sky130_fd_sc_hd__mux2_1
X_14394_ _14395_/A vssd1 vssd1 vccd1 vccd1 _14394_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_139_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16133_ _19768_/Q vssd1 vssd1 vccd1 vccd1 _16133_/Y sky130_fd_sc_hd__inv_2
X_13345_ _13428_/A _13447_/A vssd1 vssd1 vccd1 vccd1 _13346_/B sky130_fd_sc_hd__or2_2
X_10557_ _10595_/A _10559_/C _10557_/C vssd1 vssd1 vccd1 vccd1 _10581_/C sky130_fd_sc_hd__or3_4
XANTENNA_repeater237_A repeater239/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12615__A _12651_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_39_HCLK_A clkbuf_opt_1_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16064_ _16060_/Y _15828_/A _10701_/Y _15854_/X _16063_/X vssd1 vssd1 vccd1 vccd1
+ _16064_/X sky130_fd_sc_hd__o221a_1
XFILLER_182_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13276_ _18754_/Q _14270_/B _14392_/A vssd1 vssd1 vccd1 vccd1 _13276_/Y sky130_fd_sc_hd__o21ai_1
X_10488_ _19542_/Q _19541_/Q _10514_/C _10511_/A vssd1 vssd1 vccd1 vccd1 _10517_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_185_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15015_ _18047_/Q _15010_/X _14998_/X _15012_/X vssd1 vssd1 vccd1 vccd1 _18047_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_170_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12227_ _19234_/Q _12219_/X _11975_/X _12220_/X vssd1 vssd1 vccd1 vccd1 _19234_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_97_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19823_ _19825_/CLK _19823_/D repeater229/X vssd1 vssd1 vccd1 vccd1 _19823_/Q sky130_fd_sc_hd__dfrtp_1
X_12158_ _12172_/A vssd1 vssd1 vccd1 vccd1 _12158_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_229_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_229_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11109_ _11105_/Y _17754_/S _11108_/Y vssd1 vssd1 vccd1 vccd1 _11116_/A sky130_fd_sc_hd__o21ai_1
X_19754_ _19900_/CLK _19754_/D repeater196/X vssd1 vssd1 vccd1 vccd1 _19754_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_238_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12089_ _19318_/Q _12082_/X _12088_/X _12084_/X vssd1 vssd1 vccd1 vccd1 _19318_/D
+ sky130_fd_sc_hd__a22o_1
X_16966_ _16650_/Y _15536_/Y _17474_/S vssd1 vssd1 vccd1 vccd1 _16966_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18705_ _19224_/CLK _18705_/D repeater253/X vssd1 vssd1 vccd1 vccd1 _18705_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_237_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15917_ _17513_/X _15908_/X _17563_/X _16505_/A _15916_/X vssd1 vssd1 vccd1 vccd1
+ _15918_/D sky130_fd_sc_hd__o221a_2
X_19685_ _20049_/CLK _19685_/D repeater202/X vssd1 vssd1 vccd1 vccd1 _19685_/Q sky130_fd_sc_hd__dfrtp_2
X_16897_ _17473_/A0 _09905_/Y _17522_/S vssd1 vssd1 vccd1 vccd1 _16897_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13691__B1 _13682_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17352__S _17517_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_237_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18636_ _19780_/CLK _18636_/D repeater227/X vssd1 vssd1 vccd1 vccd1 _18636_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_64_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15848_ _19521_/Q vssd1 vssd1 vccd1 vccd1 _15848_/Y sky130_fd_sc_hd__inv_2
XFILLER_224_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19510__CLK _19510_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_224_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18567_ _19841_/CLK _18567_/D repeater271/X vssd1 vssd1 vccd1 vccd1 _18567_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_80_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14277__A _14277_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15779_ _19938_/Q _19365_/Q vssd1 vssd1 vccd1 vccd1 _15779_/X sky130_fd_sc_hd__and2_2
XANTENNA__19836__RESET_B repeater271/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17518_ _17517_/X _15450_/B _17518_/S vssd1 vssd1 vccd1 vccd1 _17518_/X sky130_fd_sc_hd__mux2_1
XFILLER_220_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17804__S0 _18751_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18498_ _19794_/CLK _18498_/D repeater203/X vssd1 vssd1 vccd1 vccd1 _18498_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17449_ _15963_/X _12760_/Y _17534_/S vssd1 vssd1 vccd1 vccd1 _17449_/X sky130_fd_sc_hd__mux2_1
XFILLER_178_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19119_ _19119_/CLK _19119_/D hold353/X vssd1 vssd1 vccd1 vccd1 _19119_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__16145__C1 _16144_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12525__A hold260/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18789__RESET_B repeater260/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17527__S _17539_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09178__B2 _09165_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18718__RESET_B repeater253/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09705_ _19978_/Q _09672_/Y _09635_/A _19404_/Q _09704_/X vssd1 vssd1 vccd1 vccd1
+ _09705_/X sky130_fd_sc_hd__a221o_1
XFILLER_55_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12485__B2 _12458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_243_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17262__S _17523_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15571__A _15571_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09636_ _19979_/Q vssd1 vssd1 vccd1 vccd1 _09791_/A sky130_fd_sc_hd__inv_2
XFILLER_82_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12237__A1 _19229_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09567_ _09585_/A vssd1 vssd1 vccd1 vccd1 _09567_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_15_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18758__CLK _20123_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_231_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09498_ _09473_/A _19302_/Q _09481_/A _19311_/Q vssd1 vssd1 vccd1 vccd1 _09498_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15187__B1 _10698_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16923__A1 _09420_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11460_ _11460_/A _11541_/A vssd1 vssd1 vccd1 vccd1 _11461_/B sky130_fd_sc_hd__or2_2
XPHY_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10411_ _10842_/A _14680_/A vssd1 vssd1 vccd1 vccd1 _15197_/A sky130_fd_sc_hd__or2_4
X_11391_ _19139_/Q vssd1 vssd1 vccd1 vccd1 _11391_/Y sky130_fd_sc_hd__inv_2
XFILLER_136_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10420__B1 _10418_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13130_ _19179_/Q _13080_/A _19175_/Q _13076_/A _13129_/X vssd1 vssd1 vccd1 vccd1
+ _13144_/A sky130_fd_sc_hd__o221a_1
XFILLER_125_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10342_ _10332_/B _10335_/B _10341_/X _10319_/A _19865_/Q vssd1 vssd1 vccd1 vccd1
+ _19865_/D sky130_fd_sc_hd__a32o_1
XFILLER_180_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09169__B2 _09165_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17437__S _17567_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13061_ _13061_/A _13061_/B vssd1 vssd1 vccd1 vccd1 _13062_/B sky130_fd_sc_hd__or2_2
XFILLER_140_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10273_ _11150_/B _17746_/X vssd1 vssd1 vccd1 vccd1 _10281_/B sky130_fd_sc_hd__or2b_1
XANTENNA__12173__B1 _11978_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12012_ _19356_/Q _12009_/X _09033_/X _12010_/X vssd1 vssd1 vccd1 vccd1 _19356_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_133_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10723__A1 _19772_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16820_ _16819_/X _12911_/Y _17541_/S vssd1 vssd1 vccd1 vccd1 _16820_/X sky130_fd_sc_hd__mux2_1
XFILLER_238_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16751_ _19896_/Q _19868_/Q vssd1 vssd1 vccd1 vccd1 _16751_/X sky130_fd_sc_hd__and2_4
XFILLER_46_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13963_ _18708_/Q _13966_/A _13960_/A _13901_/X vssd1 vssd1 vccd1 vccd1 _18708_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__16577__A _16687_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13673__B1 _12602_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17172__S _17536_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15702_ _15702_/A _15702_/B vssd1 vssd1 vccd1 vccd1 _15702_/Y sky130_fd_sc_hd__nor2_1
XFILLER_246_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19470_ _19470_/CLK _19470_/D repeater274/X vssd1 vssd1 vccd1 vccd1 _19470_/Q sky130_fd_sc_hd__dfrtp_1
X_12914_ _19269_/Q _18926_/Q _12913_/Y _13005_/A vssd1 vssd1 vccd1 vccd1 _12916_/C
+ sky130_fd_sc_hd__o22a_1
X_16682_ _16682_/A vssd1 vssd1 vccd1 vccd1 _16682_/X sky130_fd_sc_hd__buf_1
X_13894_ _19224_/Q vssd1 vssd1 vccd1 vccd1 _13894_/Y sky130_fd_sc_hd__inv_2
XFILLER_206_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18421_ _18441_/CLK _18421_/D vssd1 vssd1 vccd1 vccd1 _18421_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12845_ _18939_/Q vssd1 vssd1 vccd1 vccd1 _12964_/B sky130_fd_sc_hd__inv_2
X_15633_ _18602_/Q _15629_/A _15632_/Y _15629_/Y vssd1 vssd1 vccd1 vccd1 _15634_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_206_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_repeater187_A repeater188/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10239__B1 _19836_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_221_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18352_ _18959_/CLK _18352_/D vssd1 vssd1 vccd1 vccd1 _18352_/Q sky130_fd_sc_hd__dfxtp_1
X_12776_ _19227_/Q _13528_/A _12772_/Y _18823_/Q _12775_/X vssd1 vssd1 vccd1 vccd1
+ _12783_/C sky130_fd_sc_hd__o221a_1
X_15564_ _15571_/A _15564_/B vssd1 vssd1 vccd1 vccd1 _15564_/Y sky130_fd_sc_hd__nor2_1
XPHY_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11987__B1 _11926_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17303_ _17302_/X _09685_/Y _17523_/S vssd1 vssd1 vccd1 vccd1 _17303_/X sky130_fd_sc_hd__mux2_1
XPHY_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11727_ _19508_/Q _11723_/X _16940_/X _11724_/X vssd1 vssd1 vccd1 vccd1 hold214/A
+ sky130_fd_sc_hd__a22o_1
X_14515_ _18331_/Q _14504_/A hold334/X _14505_/A vssd1 vssd1 vccd1 vccd1 _18331_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_159_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18283_ _18435_/CLK _18283_/D vssd1 vssd1 vccd1 vccd1 _18283_/Q sky130_fd_sc_hd__dfxtp_1
X_15495_ _18568_/Q _15490_/A _15493_/Y _15490_/Y vssd1 vssd1 vccd1 vccd1 _15496_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_187_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17234_ _17486_/A0 _13122_/Y _17543_/S vssd1 vssd1 vccd1 vccd1 _17234_/X sky130_fd_sc_hd__mux2_1
XPHY_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11658_ _11647_/Y _15311_/A _10531_/X _10519_/D _11661_/A vssd1 vssd1 vccd1 vccd1
+ _11659_/A sky130_fd_sc_hd__o32a_1
XFILLER_30_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14446_ _18373_/Q _14436_/X _14417_/X _14439_/X vssd1 vssd1 vccd1 vccd1 _18373_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_174_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11739__B1 _16932_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10609_ _10609_/A vssd1 vssd1 vccd1 vccd1 _10609_/X sky130_fd_sc_hd__clkbuf_2
XPHY_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17165_ _17164_/X _13413_/Y _17535_/S vssd1 vssd1 vccd1 vccd1 _17165_/X sky130_fd_sc_hd__mux2_1
X_14377_ _18410_/Q _14368_/A _14314_/X _14369_/A vssd1 vssd1 vccd1 vccd1 _18410_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_100_HCLK_A clkbuf_4_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11589_ _19575_/Q _11586_/Y _11560_/C _11586_/A _11588_/X vssd1 vssd1 vccd1 vccd1
+ _19575_/D sky130_fd_sc_hd__o221a_1
XFILLER_127_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13328_ _13467_/A _13466_/A _13465_/A _13483_/B vssd1 vssd1 vccd1 vccd1 _13334_/C
+ sky130_fd_sc_hd__or4_4
XANTENNA_clkbuf_leaf_163_HCLK_A clkbuf_4_0_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16116_ _17940_/Q _16433_/B vssd1 vssd1 vccd1 vccd1 _16116_/Y sky130_fd_sc_hd__nor2_1
XFILLER_182_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17096_ _17486_/A0 _09892_/Y _17543_/S vssd1 vssd1 vccd1 vccd1 _17096_/X sky130_fd_sc_hd__mux2_1
XANTENNA__17347__S _17473_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13259_ _13259_/A _13259_/B vssd1 vssd1 vccd1 vccd1 _13262_/B sky130_fd_sc_hd__nor2_4
X_16047_ _19441_/Q vssd1 vssd1 vccd1 vccd1 _16047_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20040__CLK _20051_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19806_ _19810_/CLK _19806_/D repeater224/X vssd1 vssd1 vccd1 vccd1 _19806_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_69_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12080__A hold286/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17998_ _18416_/CLK _17998_/D vssd1 vssd1 vccd1 vccd1 _17998_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_245_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16850__A0 _16849_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19737_ _20051_/CLK _19737_/D repeater207/X vssd1 vssd1 vccd1 vccd1 _19737_/Q sky130_fd_sc_hd__dfrtp_1
X_16949_ _19493_/Q hold136/X _16950_/S vssd1 vssd1 vccd1 vccd1 _16949_/X sky130_fd_sc_hd__mux2_2
XFILLER_238_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17082__S _17473_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19668_ _19668_/CLK _19668_/D repeater270/X vssd1 vssd1 vccd1 vccd1 _19668_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_65_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09421_ _10047_/A _19391_/Q _19931_/Q _09420_/Y vssd1 vssd1 vccd1 vccd1 _09421_/X
+ sky130_fd_sc_hd__o22a_1
X_18619_ _19561_/CLK _18619_/D repeater269/X vssd1 vssd1 vccd1 vccd1 _18619_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_198_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19599_ _19600_/CLK _19599_/D hold273/X vssd1 vssd1 vccd1 vccd1 _19599_/Q sky130_fd_sc_hd__dfrtp_4
X_09352_ _20025_/Q vssd1 vssd1 vccd1 vccd1 _09485_/A sky130_fd_sc_hd__inv_2
XFILLER_100_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11442__A2 _19129_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09283_ _11842_/B vssd1 vssd1 vccd1 vccd1 _11742_/A sky130_fd_sc_hd__buf_2
XFILLER_221_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13719__A1 _18760_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19406__CLK _19984_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_opt_0_HCLK clkbuf_opt_0_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_opt_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_106_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17257__S _17490_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_22_HCLK_A clkbuf_4_3_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12155__B1 _12102_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_85_HCLK_A clkbuf_4_13_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09020__B1 _09016_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11902__B1 _09061_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08998_ _13280_/A vssd1 vssd1 vccd1 vccd1 _11936_/A sky130_fd_sc_hd__buf_2
XFILLER_85_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10960_ _19660_/Q _10999_/B vssd1 vssd1 vccd1 vccd1 _10996_/B sky130_fd_sc_hd__nand2_1
XANTENNA__17397__A1 _08959_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09619_ _20005_/Q _09618_/Y _09467_/B _09581_/X vssd1 vssd1 vccd1 vccd1 _20005_/D
+ sky130_fd_sc_hd__o211a_1
X_10891_ _19693_/Q _10878_/A _10870_/X _10879_/A vssd1 vssd1 vccd1 vccd1 _19693_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_204_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17720__S _18546_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12630_ _12630_/A vssd1 vssd1 vccd1 vccd1 _12630_/X sky130_fd_sc_hd__clkbuf_2
XPHY_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12561_ _12598_/A vssd1 vssd1 vccd1 vccd1 _12600_/A sky130_fd_sc_hd__inv_2
XPHY_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11512_ _19597_/Q _11511_/Y _11504_/X _11478_/B vssd1 vssd1 vccd1 vccd1 _19597_/D
+ sky130_fd_sc_hd__o211a_1
X_14300_ _14300_/A vssd1 vssd1 vccd1 vccd1 _15296_/B sky130_fd_sc_hd__buf_1
XPHY_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15280_ _10631_/Y _15277_/Y _15326_/A vssd1 vssd1 vccd1 vccd1 _18554_/D sky130_fd_sc_hd__o21ai_1
XPHY_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12492_ _12506_/A vssd1 vssd1 vccd1 vccd1 _12492_/X sky130_fd_sc_hd__clkbuf_2
XPHY_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10892__B _14245_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14231_ _18501_/Q _14231_/B vssd1 vssd1 vccd1 vccd1 _14232_/B sky130_fd_sc_hd__or2_1
XPHY_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11443_ _11584_/A _19151_/Q _19564_/Q _11439_/Y _11442_/X vssd1 vssd1 vccd1 vccd1
+ _11456_/B sky130_fd_sc_hd__o221a_1
XPHY_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14162_ _19107_/Q _14016_/A _16543_/A _18686_/Q _14161_/X vssd1 vssd1 vccd1 vccd1
+ _14166_/C sky130_fd_sc_hd__o221a_1
X_11374_ _19547_/Q vssd1 vssd1 vccd1 vccd1 _11639_/C sky130_fd_sc_hd__inv_2
XFILLER_4_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13113_ _19160_/Q _13062_/A _13110_/Y _18889_/Q _13112_/X vssd1 vssd1 vccd1 vccd1
+ _13113_/X sky130_fd_sc_hd__a221o_1
X_10325_ _19859_/Q _10364_/B vssd1 vssd1 vccd1 vccd1 _10361_/B sky130_fd_sc_hd__nand2_1
XANTENNA__17167__S _17566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14093_ _14093_/A _14093_/B _14093_/C _14093_/D vssd1 vssd1 vccd1 vccd1 _14093_/X
+ sky130_fd_sc_hd__and4_1
X_18970_ _19582_/CLK _18970_/D hold348/A vssd1 vssd1 vccd1 vccd1 _18970_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_180_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12146__B1 _12086_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17921_ _18393_/Q _18385_/Q _18377_/Q _18369_/Q _17923_/S0 _19646_/Q vssd1 vssd1
+ vccd1 vccd1 _17921_/X sky130_fd_sc_hd__mux4_2
X_13044_ _18902_/Q vssd1 vssd1 vccd1 vccd1 _13074_/A sky130_fd_sc_hd__inv_2
X_10256_ _19627_/Q _10409_/A _15190_/A vssd1 vssd1 vccd1 vccd1 _14300_/A sky130_fd_sc_hd__or3_4
XFILLER_239_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17852_ _16336_/Y _16337_/Y _16338_/Y _16339_/Y _17913_/S0 _19632_/Q vssd1 vssd1
+ vccd1 vccd1 _17852_/X sky130_fd_sc_hd__mux4_1
XFILLER_94_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10187_ _09339_/X _19875_/Q _10188_/S vssd1 vssd1 vccd1 vccd1 _19875_/D sky130_fd_sc_hd__mux2_1
XFILLER_79_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16832__A0 _15963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16803_ _16802_/X _09492_/A _17482_/S vssd1 vssd1 vccd1 vccd1 _16803_/X sky130_fd_sc_hd__mux2_1
XFILLER_66_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17783_ _18293_/Q _18285_/Q _18277_/Q _18445_/Q _17923_/S0 _19646_/Q vssd1 vssd1
+ vccd1 vccd1 _17783_/X sky130_fd_sc_hd__mux4_2
X_14995_ _18057_/Q _14991_/X _14992_/X _14994_/X vssd1 vssd1 vccd1 vccd1 _18057_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19522_ _20049_/CLK _19522_/D repeater190/X vssd1 vssd1 vccd1 vccd1 _19522_/Q sky130_fd_sc_hd__dfstp_1
X_16734_ _16771_/X _16687_/X _16788_/X _16688_/X _16733_/X vssd1 vssd1 vccd1 vccd1
+ _16735_/C sky130_fd_sc_hd__o221a_1
XFILLER_235_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13946_ _13946_/A _13960_/A vssd1 vssd1 vccd1 vccd1 _13947_/B sky130_fd_sc_hd__or2_2
XFILLER_62_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19453_ _19462_/CLK _19453_/D repeater272/X vssd1 vssd1 vccd1 vccd1 _19453_/Q sky130_fd_sc_hd__dfrtp_1
X_16665_ _16665_/A _16668_/B vssd1 vssd1 vccd1 vccd1 _16665_/Y sky130_fd_sc_hd__nor2_1
XFILLER_90_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13877_ _13875_/Y _18711_/Q _19200_/Q _13948_/A _13876_/X vssd1 vssd1 vccd1 vccd1
+ _13882_/C sky130_fd_sc_hd__o221a_1
XFILLER_62_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18404_ _18954_/CLK _18404_/D vssd1 vssd1 vccd1 vccd1 _18404_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10880__B1 _10877_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15616_ _18598_/Q vssd1 vssd1 vccd1 vccd1 _15618_/A sky130_fd_sc_hd__inv_2
XFILLER_201_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12828_ _18820_/Q vssd1 vssd1 vccd1 vccd1 _13543_/A sky130_fd_sc_hd__inv_2
XANTENNA__09078__B1 _09077_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19384_ _19927_/CLK _19384_/D repeater235/X vssd1 vssd1 vccd1 vccd1 _19384_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16596_ _17260_/X _16594_/X _17258_/X _16595_/X vssd1 vssd1 vccd1 vccd1 _16600_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_188_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18335_ _19849_/CLK _18335_/D vssd1 vssd1 vccd1 vccd1 _18335_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15547_ _18580_/Q _15547_/B vssd1 vssd1 vccd1 vccd1 _15547_/X sky130_fd_sc_hd__and2_1
X_12759_ _18806_/Q vssd1 vssd1 vccd1 vccd1 _13530_/A sky130_fd_sc_hd__inv_2
XFILLER_187_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18266_ _18268_/CLK _18266_/D vssd1 vssd1 vccd1 vccd1 _18266_/Q sky130_fd_sc_hd__dfxtp_1
X_15478_ _18564_/Q _15474_/A _15477_/Y _15474_/Y vssd1 vssd1 vccd1 vccd1 _15479_/B
+ sky130_fd_sc_hd__o22a_1
X_17217_ _17216_/X _12919_/Y _17487_/S vssd1 vssd1 vccd1 vccd1 _17217_/X sky130_fd_sc_hd__mux2_1
X_14429_ _18383_/Q _14424_/X _14359_/X _14426_/X vssd1 vssd1 vccd1 vccd1 _18383_/D
+ sky130_fd_sc_hd__a22o_1
X_18197_ _18216_/CLK _18197_/D vssd1 vssd1 vccd1 vccd1 _18197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12385__B1 _12384_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17148_ _17147_/X _09717_/Y _17517_/S vssd1 vssd1 vccd1 vccd1 _17148_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17312__A1 _18779_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17077__S _17543_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09970_ _09990_/A vssd1 vssd1 vccd1 vccd1 _09970_/X sky130_fd_sc_hd__buf_2
X_17079_ _17078_/X _13085_/A _17542_/S vssd1 vssd1 vccd1 vccd1 _17079_/X sky130_fd_sc_hd__mux2_2
XFILLER_115_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12803__A _19231_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08921_ _10321_/A vssd1 vssd1 vccd1 vccd1 _08921_/X sky130_fd_sc_hd__clkbuf_2
X_20090_ _20090_/CLK _20090_/D repeater204/X vssd1 vssd1 vccd1 vccd1 _20090_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12688__A1 _18974_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10163__A2 _10155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19851__RESET_B repeater258/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09404_ _10086_/A _19374_/Q _10086_/A _19374_/Q vssd1 vssd1 vccd1 vccd1 _09404_/X
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__17540__S _17543_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10871__B1 _10870_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16664__B _16664_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09335_ _13766_/D vssd1 vssd1 vccd1 vccd1 _15727_/B sky130_fd_sc_hd__inv_2
Xclkbuf_2_3_0_HCLK clkbuf_2_3_0_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__17000__A0 _15768_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09266_ _19497_/Q vssd1 vssd1 vccd1 vccd1 _11842_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__17551__A1 _19741_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09197_ _17605_/X _09197_/B vssd1 vssd1 vccd1 vccd1 _09205_/B sky130_fd_sc_hd__or2_2
XFILLER_119_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17926__D _19814_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15296__A _15296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12128__B1 _11924_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10110_ _18581_/Q _18580_/Q vssd1 vssd1 vccd1 vccd1 _10126_/C sky130_fd_sc_hd__or2_1
XFILLER_20_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12679__A1 _18981_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11090_ _15318_/A _15295_/B vssd1 vssd1 vccd1 vccd1 _11106_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19939__RESET_B hold371/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10041_ _10041_/A _10068_/A vssd1 vssd1 vccd1 vccd1 _10042_/B sky130_fd_sc_hd__or2_2
XANTENNA__17715__S _18546_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17970__CLK _20123_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19592__RESET_B hold346/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13800_ _18706_/Q vssd1 vssd1 vccd1 vccd1 _13802_/B sky130_fd_sc_hd__inv_2
XFILLER_152_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14780_ _14780_/A vssd1 vssd1 vccd1 vccd1 _14780_/X sky130_fd_sc_hd__buf_2
X_11992_ _15776_/A _11998_/A vssd1 vssd1 vccd1 vccd1 _11993_/S sky130_fd_sc_hd__or2_1
XFILLER_205_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10943_ _18512_/Q _15298_/D _15213_/A _15298_/C vssd1 vssd1 vccd1 vccd1 _10943_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_72_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13731_ _13725_/A _14392_/A _14758_/B vssd1 vssd1 vccd1 vccd1 _13731_/X sky130_fd_sc_hd__o21a_1
XFILLER_90_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17450__S _17535_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16450_ _19528_/Q vssd1 vssd1 vccd1 vccd1 _16450_/Y sky130_fd_sc_hd__inv_2
XANTENNA__10862__B1 _10861_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10874_ _15973_/A _14245_/D vssd1 vssd1 vccd1 vccd1 _10878_/A sky130_fd_sc_hd__or2_2
X_13662_ _18784_/Q _13656_/X _12032_/A _13658_/X vssd1 vssd1 vccd1 vccd1 _18784_/D
+ sky130_fd_sc_hd__a22o_1
X_15401_ _18533_/Q _13220_/B _13221_/B vssd1 vssd1 vccd1 vccd1 _15401_/X sky130_fd_sc_hd__a21bo_1
XPHY_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12613_ _12629_/A vssd1 vssd1 vccd1 vccd1 _12613_/X sky130_fd_sc_hd__buf_1
XFILLER_231_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13593_ _13539_/A _13593_/A2 _13588_/X _13590_/Y vssd1 vssd1 vccd1 vccd1 _18816_/D
+ sky130_fd_sc_hd__a211oi_2
X_16381_ _19527_/Q vssd1 vssd1 vccd1 vccd1 _16381_/Y sky130_fd_sc_hd__inv_2
XPHY_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18120_ _18169_/CLK _18120_/D vssd1 vssd1 vccd1 vccd1 _18120_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_185_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15332_ _18518_/Q vssd1 vssd1 vccd1 vccd1 _15850_/A sky130_fd_sc_hd__inv_2
X_12544_ _19061_/Q _12505_/A _12543_/X _12506_/A vssd1 vssd1 vccd1 vccd1 _19061_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_184_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18051_ _18142_/CLK _18051_/D vssd1 vssd1 vccd1 vccd1 _18051_/Q sky130_fd_sc_hd__dfxtp_1
X_15263_ _15263_/A vssd1 vssd1 vccd1 vccd1 _15263_/Y sky130_fd_sc_hd__inv_2
X_12475_ _19102_/Q _12471_/X _12223_/X _12472_/X vssd1 vssd1 vccd1 vccd1 _19102_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12367__B1 _12236_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17002_ _17001_/X _11423_/Y _17548_/S vssd1 vssd1 vccd1 vccd1 _17002_/X sky130_fd_sc_hd__mux2_1
X_11426_ _11561_/A _11425_/Y _19576_/Q _19156_/Q vssd1 vssd1 vccd1 vccd1 _11426_/X
+ sky130_fd_sc_hd__a22o_1
X_14214_ _19097_/Q _14007_/A _16209_/A _18676_/Q _14213_/X vssd1 vssd1 vccd1 vccd1
+ _14218_/C sky130_fd_sc_hd__o221a_1
XFILLER_126_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15194_ _18757_/Q vssd1 vssd1 vccd1 vccd1 _15194_/Y sky130_fd_sc_hd__inv_2
X_14145_ _14145_/A vssd1 vssd1 vccd1 vccd1 _14145_/Y sky130_fd_sc_hd__clkinv_1
X_11357_ _19590_/Q _11354_/Y _19598_/Q _11355_/Y _11356_/X vssd1 vssd1 vccd1 vccd1
+ _11361_/C sky130_fd_sc_hd__o221a_1
XANTENNA__19871__CLK _20070_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12119__B1 _11911_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10308_ _18605_/Q _18606_/Q _10308_/C _15668_/A vssd1 vssd1 vccd1 vccd1 _10309_/B
+ sky130_fd_sc_hd__or4_1
XANTENNA_output79_A _15918_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14076_ _19087_/Q _14028_/A _14072_/Y _18672_/Q _14075_/X vssd1 vssd1 vccd1 vccd1
+ _14080_/C sky130_fd_sc_hd__o221a_1
X_18953_ _18959_/CLK _18953_/D repeater257/X vssd1 vssd1 vccd1 vccd1 _18953_/Q sky130_fd_sc_hd__dfrtp_1
X_11288_ _19593_/Q vssd1 vssd1 vccd1 vccd1 _11473_/A sky130_fd_sc_hd__inv_2
XFILLER_193_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17904_ _17900_/X _17901_/X _17902_/X _17903_/X _19633_/Q _19634_/Q vssd1 vssd1 vccd1
+ vccd1 _17904_/X sky130_fd_sc_hd__mux4_2
X_13027_ _13027_/A _13027_/B _13027_/C vssd1 vssd1 vccd1 vccd1 _18920_/D sky130_fd_sc_hd__nor3_1
XFILLER_239_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10239_ _10234_/Y _19666_/Q _19836_/Q _10963_/A _10238_/X vssd1 vssd1 vccd1 vccd1
+ _10246_/C sky130_fd_sc_hd__o221a_1
X_18884_ _18886_/CLK _18884_/D repeater220/X vssd1 vssd1 vccd1 vccd1 _18884_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__19609__RESET_B hold359/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17835_ _16417_/Y _16418_/Y _16419_/Y _16420_/Y _17908_/S0 _18759_/Q vssd1 vssd1
+ vccd1 vccd1 _17835_/X sky130_fd_sc_hd__mux4_2
XFILLER_48_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrebuffer18 _14024_/B vssd1 vssd1 vccd1 vccd1 _14117_/C1 sky130_fd_sc_hd__dlygate4sd1_1
X_17766_ _18386_/Q _18378_/Q _18370_/Q _18362_/Q _17923_/S0 _19646_/Q vssd1 vssd1
+ vccd1 vccd1 _17766_/X sky130_fd_sc_hd__mux4_2
XANTENNA__09299__B1 _09108_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrebuffer29 _14011_/B vssd1 vssd1 vccd1 vccd1 _14138_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XANTENNA__14292__B1 _14277_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14978_ _14978_/A vssd1 vssd1 vccd1 vccd1 _14979_/A sky130_fd_sc_hd__inv_2
XANTENNA__19262__RESET_B repeater212/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19505_ _19506_/CLK hold221/X repeater256/X vssd1 vssd1 vccd1 vccd1 _19505_/Q sky130_fd_sc_hd__dfrtp_1
X_16717_ _16717_/A _16718_/B vssd1 vssd1 vccd1 vccd1 _16717_/Y sky130_fd_sc_hd__nor2_1
X_13929_ _13929_/A vssd1 vssd1 vccd1 vccd1 _13929_/Y sky130_fd_sc_hd__inv_2
X_17697_ _19821_/Q _19763_/Q _18548_/Q vssd1 vssd1 vccd1 vccd1 _17697_/X sky130_fd_sc_hd__mux2_1
XFILLER_235_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17360__S _17543_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10853__B1 _10427_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19436_ _19905_/CLK _19436_/D repeater210/X vssd1 vssd1 vccd1 vccd1 _19436_/Q sky130_fd_sc_hd__dfrtp_1
X_16648_ _16669_/A vssd1 vssd1 vccd1 vccd1 _16668_/B sky130_fd_sc_hd__buf_4
XFILLER_90_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19367_ _20091_/CLK _19367_/D repeater236/X vssd1 vssd1 vccd1 vccd1 _19367_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_176_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16579_ _17263_/X _15889_/X _17254_/X _15887_/X vssd1 vssd1 vccd1 vccd1 _16579_/X
+ sky130_fd_sc_hd__o22a_1
X_09120_ _09120_/A vssd1 vssd1 vccd1 vccd1 _15319_/A sky130_fd_sc_hd__buf_1
X_18318_ _19637_/CLK _18318_/D vssd1 vssd1 vccd1 vccd1 _18318_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19298_ _20013_/CLK _19298_/D repeater242/X vssd1 vssd1 vccd1 vccd1 _19298_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_31_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrebuffer108 _13079_/B vssd1 vssd1 vccd1 vccd1 _13183_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_30_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrebuffer119 _11472_/B vssd1 vssd1 vccd1 vccd1 _11519_/A2 sky130_fd_sc_hd__dlygate4sd1_1
X_09051_ hold294/X vssd1 vssd1 vccd1 vccd1 _09051_/X sky130_fd_sc_hd__buf_4
X_18249_ _18465_/CLK _18249_/D vssd1 vssd1 vccd1 vccd1 _18249_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12358__B1 _12223_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17297__A0 _17486_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12533__A hold325/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17993__CLK _18169_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09953_ _09877_/A _09877_/B _09878_/Y _09987_/B vssd1 vssd1 vccd1 vccd1 _19969_/D
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__17049__A0 _15768_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17535__S _17535_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20073_ _20124_/CLK _20073_/D repeater196/X vssd1 vssd1 vccd1 vccd1 _20073_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_58_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09884_ _19350_/Q vssd1 vssd1 vccd1 vccd1 _09884_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12530__B1 _12299_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14283__B1 _13678_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_151_HCLK clkbuf_4_1_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19873_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_66_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17270__S _17522_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16575__A2 _16394_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19744__CLK _20070_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_213_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12597__B1 _12596_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18914__RESET_B repeater188/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09318_ _18654_/Q _09317_/X _18656_/Q vssd1 vssd1 vccd1 vccd1 _09318_/Y sky130_fd_sc_hd__a21oi_1
X_10590_ _19798_/Q _19797_/Q _19813_/Q _10590_/D vssd1 vssd1 vccd1 vccd1 _10593_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_22_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16327__A2 _16310_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09249_ _20062_/Q _20063_/Q _09250_/S vssd1 vssd1 vccd1 vccd1 _20063_/D sky130_fd_sc_hd__mux2_1
XFILLER_139_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16732__C1 _16731_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12349__B1 hold256/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12260_ _12276_/A vssd1 vssd1 vccd1 vccd1 _12260_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_108_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17288__A0 _15963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11211_ _19015_/Q vssd1 vssd1 vccd1 vccd1 _11211_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12191_ _12229_/A vssd1 vssd1 vccd1 vccd1 _12206_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_123_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11142_ _12253_/A _11133_/Y _11139_/Y _19630_/Q _11141_/X vssd1 vssd1 vccd1 vccd1
+ _19630_/D sky130_fd_sc_hd__a32o_1
Xoutput87 _16600_/X vssd1 vssd1 vccd1 vccd1 HRDATA[17] sky130_fd_sc_hd__clkbuf_2
XANTENNA__17445__S _17518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11073_ _14477_/B _11072_/Y _14477_/B _11072_/Y vssd1 vssd1 vccd1 vccd1 _11076_/C
+ sky130_fd_sc_hd__a2bb2o_1
X_15950_ _18259_/Q vssd1 vssd1 vccd1 vccd1 _15950_/Y sky130_fd_sc_hd__inv_2
Xoutput98 _16705_/Y vssd1 vssd1 vccd1 vccd1 HRDATA[27] sky130_fd_sc_hd__clkbuf_2
XANTENNA__12521__B1 _12353_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10024_ _10024_/A vssd1 vssd1 vccd1 vccd1 _10032_/B sky130_fd_sc_hd__inv_2
X_14901_ _18111_/Q _14896_/X _14705_/X _14898_/X vssd1 vssd1 vccd1 vccd1 _18111_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_48_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15881_ _19438_/Q _15881_/B vssd1 vssd1 vccd1 vccd1 _15881_/Y sky130_fd_sc_hd__nor2_1
X_17620_ _20052_/Q _19726_/Q _17621_/S vssd1 vssd1 vccd1 vccd1 _17620_/X sky130_fd_sc_hd__mux2_1
X_14832_ _14833_/A vssd1 vssd1 vccd1 vccd1 _14832_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_56_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17551_ _18737_/Q _19741_/Q _19499_/Q vssd1 vssd1 vccd1 vccd1 _17551_/X sky130_fd_sc_hd__mux2_1
X_14763_ _18192_/Q _14759_/X _14749_/X _14761_/X vssd1 vssd1 vccd1 vccd1 _18192_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_245_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11975_ _14273_/A vssd1 vssd1 vccd1 vccd1 _11975_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_44_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17212__A0 _17473_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16502_ _19449_/Q vssd1 vssd1 vccd1 vccd1 _16502_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17180__S _17541_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13714_ _13706_/A _13704_/B _17761_/X _17908_/S0 vssd1 vssd1 vccd1 vccd1 _18758_/D
+ sky130_fd_sc_hd__o22a_1
X_10926_ _17722_/X _10923_/X _19679_/Q _10924_/X vssd1 vssd1 vccd1 vccd1 _19679_/D
+ sky130_fd_sc_hd__a22o_1
X_17482_ _17481_/X _09466_/A _17482_/S vssd1 vssd1 vccd1 vccd1 _17482_/X sky130_fd_sc_hd__mux2_2
XFILLER_189_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14694_ _18226_/Q _14683_/A _14693_/X _14684_/A vssd1 vssd1 vccd1 vccd1 _18226_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16566__A2 _16684_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19221_ _19221_/CLK _19221_/D repeater186/X vssd1 vssd1 vccd1 vccd1 _19221_/Q sky130_fd_sc_hd__dfrtp_1
X_16433_ _17944_/Q _16433_/B vssd1 vssd1 vccd1 vccd1 _16433_/X sky130_fd_sc_hd__or2_1
XFILLER_220_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10857_ _10857_/A vssd1 vssd1 vccd1 vccd1 _10857_/X sky130_fd_sc_hd__clkbuf_2
X_13645_ _17924_/X _15201_/B _13646_/A _18795_/Q _13644_/X vssd1 vssd1 vccd1 vccd1
+ _18795_/D sky130_fd_sc_hd__a32o_1
XANTENNA__12588__B1 hold256/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18655__RESET_B repeater210/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19152_ _19597_/CLK _19152_/D repeater281/X vssd1 vssd1 vccd1 vccd1 _19152_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16364_ _17343_/X _16415_/B vssd1 vssd1 vccd1 vccd1 _16364_/X sky130_fd_sc_hd__and2_1
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13576_ _13549_/A _13576_/A2 _13571_/X _13573_/Y vssd1 vssd1 vccd1 vccd1 _18826_/D
+ sky130_fd_sc_hd__a211oi_2
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10788_ _18653_/Q vssd1 vssd1 vccd1 vccd1 _10788_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18103_ _18137_/CLK _18103_/D vssd1 vssd1 vccd1 vccd1 _18103_/Q sky130_fd_sc_hd__dfxtp_1
X_15315_ _18626_/Q vssd1 vssd1 vccd1 vccd1 _15315_/Y sky130_fd_sc_hd__inv_2
X_19083_ _19119_/CLK _19083_/D hold355/X vssd1 vssd1 vccd1 vccd1 _19083_/Q sky130_fd_sc_hd__dfrtp_1
X_12527_ _19068_/Q _12519_/X _12296_/X _12520_/X vssd1 vssd1 vccd1 vccd1 _19068_/D
+ sky130_fd_sc_hd__a22o_1
X_16295_ _17942_/Q _16433_/B vssd1 vssd1 vccd1 vccd1 _16295_/X sky130_fd_sc_hd__or2_1
XFILLER_200_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18034_ _19851_/CLK _18034_/D vssd1 vssd1 vccd1 vccd1 _18034_/Q sky130_fd_sc_hd__dfxtp_1
X_15246_ _15242_/Y _15243_/Y _15245_/X vssd1 vssd1 vccd1 vccd1 _15246_/Y sky130_fd_sc_hd__a21oi_1
X_12458_ _12458_/A vssd1 vssd1 vccd1 vccd1 _12458_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_32_HCLK _18641_/CLK vssd1 vssd1 vccd1 vccd1 _20124_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_172_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11409_ _19149_/Q vssd1 vssd1 vccd1 vccd1 _11409_/Y sky130_fd_sc_hd__inv_2
X_12389_ hold303/X vssd1 vssd1 vccd1 vccd1 _12389_/X sky130_fd_sc_hd__buf_2
X_15177_ _17940_/Q _15170_/X _10715_/X _15172_/X vssd1 vssd1 vccd1 vccd1 _17940_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_181_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14128_ _14016_/A _14128_/A2 _14126_/Y _14118_/X vssd1 vssd1 vccd1 vccd1 _18686_/D
+ sky130_fd_sc_hd__a211oi_2
X_19985_ _19992_/CLK _19985_/D repeater193/X vssd1 vssd1 vccd1 vccd1 _19985_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_113_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17355__S _17413_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18936_ _19315_/CLK _18936_/D repeater213/X vssd1 vssd1 vccd1 vccd1 _18936_/Q sky130_fd_sc_hd__dfrtp_1
X_14059_ _19061_/Q _14003_/A _14039_/Y _18691_/Q _14058_/X vssd1 vssd1 vccd1 vccd1
+ _14059_/X sky130_fd_sc_hd__o221a_1
XFILLER_141_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18867_ _20122_/CLK _18867_/D repeater234/X vssd1 vssd1 vccd1 vccd1 _18867_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_227_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17818_ _17931_/Q _18453_/Q _18461_/Q _18061_/Q _17918_/S0 _18750_/Q vssd1 vssd1
+ vccd1 vccd1 _17818_/X sky130_fd_sc_hd__mux4_2
XFILLER_94_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18641__CLK _18641_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18798_ _19435_/CLK _18798_/D repeater258/X vssd1 vssd1 vccd1 vccd1 _18798_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_242_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17749_ _15753_/B _18879_/Q _17749_/S vssd1 vssd1 vccd1 vccd1 _17749_/X sky130_fd_sc_hd__mux2_2
XANTENNA__17203__A0 _15963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17090__S _17543_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17754__A1 _11093_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16557__A2 _16597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19419_ _19997_/CLK _19419_/D repeater192/X vssd1 vssd1 vccd1 vccd1 _19419_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_168_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12528__A _12528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12579__B1 _12404_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09103_ hold336/X vssd1 vssd1 vccd1 vccd1 _14780_/A sky130_fd_sc_hd__buf_2
XFILLER_248_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15839__A _15839_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16714__C1 _16713_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09034_ _20116_/Q _09029_/X _09033_/X _09031_/X vssd1 vssd1 vccd1 vccd1 _20116_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_175_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold320 hold320/A vssd1 vssd1 vccd1 vccd1 hold320/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold331 hold331/A vssd1 vssd1 vccd1 vccd1 hold331/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold342 MSI_S2 vssd1 vssd1 vccd1 vccd1 input71/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold353 hold353/A vssd1 vssd1 vccd1 vccd1 hold353/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold364 hold364/A vssd1 vssd1 vccd1 vccd1 hold364/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__19297__CLK _20013_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17265__S _17413_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09936_ _19940_/Q _09934_/Y _19966_/Q _09935_/Y vssd1 vssd1 vccd1 vccd1 _09936_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_131_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11306__B2 _18974_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12503__B1 _12396_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20056_ _20057_/CLK _20056_/D repeater204/X vssd1 vssd1 vccd1 vccd1 _20056_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_97_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09867_ _09867_/A _09867_/B vssd1 vssd1 vccd1 vccd1 _09967_/A sky130_fd_sc_hd__or2_1
XANTENNA__20089__RESET_B repeater204/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09798_ _19981_/Q _09797_/Y _09794_/B _09731_/X vssd1 vssd1 vccd1 vccd1 _19981_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_4302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater170 _17386_/S vssd1 vssd1 vccd1 vccd1 _17536_/S sky130_fd_sc_hd__buf_8
Xrepeater181 _19645_/Q vssd1 vssd1 vccd1 vccd1 _17923_/S0 sky130_fd_sc_hd__clkbuf_16
XPHY_4313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater192 repeater193/X vssd1 vssd1 vccd1 vccd1 repeater192/X sky130_fd_sc_hd__buf_8
XPHY_4324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11760_ hold165/X _11757_/X _19484_/Q _11758_/X vssd1 vssd1 vccd1 vccd1 hold167/A
+ sky130_fd_sc_hd__o22a_1
XPHY_4368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10711_ _19774_/Q vssd1 vssd1 vccd1 vccd1 _15753_/A sky130_fd_sc_hd__inv_2
XPHY_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11691_ _11691_/A vssd1 vssd1 vccd1 vccd1 _11692_/A sky130_fd_sc_hd__inv_2
XPHY_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17840__S1 _19632_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13430_ _13430_/A _13430_/B _13430_/C _13430_/D vssd1 vssd1 vccd1 vccd1 _13431_/B
+ sky130_fd_sc_hd__or4_4
X_10642_ _19782_/Q _19781_/Q vssd1 vssd1 vccd1 vccd1 _10643_/B sky130_fd_sc_hd__or2_1
XPHY_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_55_HCLK clkbuf_opt_3_HCLK/A vssd1 vssd1 vccd1 vccd1 _19771_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13361_ _18864_/Q vssd1 vssd1 vccd1 vccd1 _13361_/Y sky130_fd_sc_hd__inv_2
XFILLER_158_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10573_ _19808_/Q _10573_/B _10574_/A vssd1 vssd1 vccd1 vccd1 _10575_/A sky130_fd_sc_hd__nor3_4
XFILLER_182_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15100_ _17991_/Q _15095_/X _14808_/A _15097_/X vssd1 vssd1 vccd1 vccd1 _17991_/D
+ sky130_fd_sc_hd__a22o_1
Xrebuffer9 _13075_/B vssd1 vssd1 vccd1 vccd1 _13191_/C1 sky130_fd_sc_hd__dlygate4sd1_1
X_12312_ _12180_/X _19191_/Q _12312_/S vssd1 vssd1 vccd1 vccd1 _19191_/D sky130_fd_sc_hd__mux2_1
X_16080_ _18029_/Q vssd1 vssd1 vccd1 vccd1 _16080_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13292_ _18755_/Q vssd1 vssd1 vccd1 vccd1 _13729_/A sky130_fd_sc_hd__inv_2
XANTENNA__11996__B _16053_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19954__RESET_B repeater245/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15031_ _18036_/Q _15024_/A _15004_/X _15025_/A vssd1 vssd1 vccd1 vccd1 _18036_/D
+ sky130_fd_sc_hd__a22o_1
X_12243_ _12708_/B vssd1 vssd1 vccd1 vccd1 _15232_/B sky130_fd_sc_hd__buf_1
XFILLER_170_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12174_ _19267_/Q _12171_/X _11981_/X _12172_/X vssd1 vssd1 vccd1 vccd1 _19267_/D
+ sky130_fd_sc_hd__a22o_1
X_11125_ _19634_/Q _11127_/A _11060_/Y _11124_/A vssd1 vssd1 vccd1 vccd1 _19634_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_122_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17175__S _17542_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19770_ _19771_/CLK _19770_/D repeater228/X vssd1 vssd1 vccd1 vccd1 _19770_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_3_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16982_ _17814_/X _19900_/Q _16986_/S vssd1 vssd1 vccd1 vccd1 _16982_/X sky130_fd_sc_hd__mux2_1
XFILLER_123_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18721_ _18727_/CLK _18721_/D repeater253/X vssd1 vssd1 vccd1 vccd1 _18721_/Q sky130_fd_sc_hd__dfrtp_1
X_11056_ _11056_/A _14316_/B vssd1 vssd1 vccd1 vccd1 _11056_/Y sky130_fd_sc_hd__nor2_1
X_15933_ _18467_/Q vssd1 vssd1 vccd1 vccd1 _15933_/Y sky130_fd_sc_hd__inv_2
XFILLER_236_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10007_ _10081_/B vssd1 vssd1 vccd1 vccd1 _10101_/B sky130_fd_sc_hd__clkbuf_2
X_18652_ _20124_/CLK hold341/X repeater205/X vssd1 vssd1 vccd1 vccd1 _18652_/Q sky130_fd_sc_hd__dfrtp_1
X_15864_ _15867_/A _15864_/B vssd1 vssd1 vccd1 vccd1 _17530_/S sky130_fd_sc_hd__nor2_8
XFILLER_236_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17603_ _15320_/Y _13495_/B _17605_/S vssd1 vssd1 vccd1 vccd1 _17603_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14815_ _18164_/Q _14803_/A _14814_/X _14804_/A vssd1 vssd1 vccd1 vccd1 _18164_/D
+ sky130_fd_sc_hd__a22o_1
X_18583_ _19970_/CLK _18583_/D repeater274/X vssd1 vssd1 vccd1 vccd1 _18583_/Q sky130_fd_sc_hd__dfrtp_1
X_15795_ _18402_/Q vssd1 vssd1 vccd1 vccd1 _15795_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18836__RESET_B repeater196/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17534_ _17533_/X _12797_/Y _17534_/S vssd1 vssd1 vccd1 vccd1 _17534_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14746_ _14746_/A vssd1 vssd1 vccd1 vccd1 _14747_/A sky130_fd_sc_hd__inv_2
X_11958_ _19386_/Q _11955_/X hold300/X _11956_/X vssd1 vssd1 vccd1 vccd1 _19386_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16539__A2 _16684_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10909_ _10909_/A vssd1 vssd1 vccd1 vccd1 _15384_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_199_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17465_ _17464_/X _08941_/Y _17566_/S vssd1 vssd1 vccd1 vccd1 _17465_/X sky130_fd_sc_hd__mux2_1
XANTENNA__17831__S1 _18750_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14677_ _18236_/Q _14670_/A _09183_/X _14671_/A vssd1 vssd1 vccd1 vccd1 _18236_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_60_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11889_ _19424_/Q _11884_/X _09037_/X _11885_/X vssd1 vssd1 vccd1 vccd1 _19424_/D
+ sky130_fd_sc_hd__a22o_1
X_19204_ _19585_/CLK _19204_/D hold365/X vssd1 vssd1 vccd1 vccd1 _19204_/Q sky130_fd_sc_hd__dfrtp_4
X_16416_ _17315_/X _16435_/B vssd1 vssd1 vccd1 vccd1 _16416_/Y sky130_fd_sc_hd__nand2_1
X_13628_ _18800_/Q _13620_/Y _18800_/Q _13620_/Y vssd1 vssd1 vccd1 vccd1 _18800_/D
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_220_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17396_ _17395_/X _16201_/Y _17565_/S vssd1 vssd1 vccd1 vccd1 _17396_/X sky130_fd_sc_hd__mux2_1
XFILLER_186_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19135_ _19137_/CLK _19135_/D repeater249/X vssd1 vssd1 vccd1 vccd1 _19135_/Q sky130_fd_sc_hd__dfrtp_1
X_16347_ _18128_/Q vssd1 vssd1 vccd1 vccd1 _16347_/Y sky130_fd_sc_hd__inv_2
X_13559_ _13588_/A vssd1 vssd1 vccd1 vccd1 _13591_/A sky130_fd_sc_hd__inv_2
XFILLER_173_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19066_ _19585_/CLK _19066_/D hold361/X vssd1 vssd1 vccd1 vccd1 _19066_/Q sky130_fd_sc_hd__dfrtp_1
X_16278_ _17974_/Q vssd1 vssd1 vccd1 vccd1 _16278_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16711__A2 _16493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19695__RESET_B repeater208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18017_ _18959_/CLK _18017_/D vssd1 vssd1 vccd1 vccd1 _18017_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15229_ _15278_/B _15229_/B vssd1 vssd1 vccd1 vccd1 _15386_/A sky130_fd_sc_hd__or2_2
XANTENNA__12083__A hold303/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17898__S1 _18759_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17085__S _17544_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16475__A1 _08962_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16475__B2 _16506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19968_ _19968_/CLK _19968_/D repeater185/X vssd1 vssd1 vccd1 vccd1 _19968_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_234_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09721_ _19987_/Q _09720_/Y _09743_/A _19416_/Q vssd1 vssd1 vccd1 vccd1 _09721_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_228_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18919_ _18947_/CLK _18919_/D repeater211/X vssd1 vssd1 vccd1 vccd1 _18919_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_110_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17424__A0 _15768_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19899_ _19900_/CLK _19899_/D repeater195/X vssd1 vssd1 vccd1 vccd1 _19899_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_67_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09652_ _19985_/Q vssd1 vssd1 vccd1 vccd1 _09741_/A sky130_fd_sc_hd__inv_2
XFILLER_216_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20111__RESET_B repeater217/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09583_ _09486_/A _09486_/B _09580_/Y _09604_/B vssd1 vssd1 vccd1 vccd1 _20026_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_82_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17727__A1 _19686_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18506__RESET_B repeater233/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_78_HCLK clkbuf_4_13_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19324_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17822__S1 _18750_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12258__A _12372_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16672__B _16673_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11775__A1 hold199/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09017_ _09084_/A vssd1 vssd1 vccd1 vccd1 _09087_/A sky130_fd_sc_hd__inv_2
XFILLER_12_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19365__RESET_B repeater210/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold150 hold150/A vssd1 vssd1 vccd1 vccd1 hold150/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold161 hold161/A vssd1 vssd1 vccd1 vccd1 hold161/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17889__S1 _18761_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold172 HADDR[19] vssd1 vssd1 vccd1 vccd1 input11/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 input28/X vssd1 vssd1 vccd1 vccd1 hold183/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 HADDR[0] vssd1 vssd1 vccd1 vccd1 input1/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15674__C1 _15673_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20108_ _20120_/CLK _20108_/D repeater217/X vssd1 vssd1 vccd1 vccd1 _20108_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_144_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09919_ _19962_/Q _09918_/Y _09859_/A _19343_/Q vssd1 vssd1 vccd1 vccd1 _09919_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_59_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17415__A0 _15963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20039_ _20051_/CLK _20039_/D repeater206/X vssd1 vssd1 vccd1 vccd1 _20039_/Q sky130_fd_sc_hd__dfrtp_1
X_12930_ _19266_/Q vssd1 vssd1 vccd1 vccd1 _12930_/Y sky130_fd_sc_hd__inv_2
XFILLER_219_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12861_ _18925_/Q vssd1 vssd1 vccd1 vccd1 _13004_/A sky130_fd_sc_hd__inv_2
XFILLER_234_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14600_ _14745_/A vssd1 vssd1 vccd1 vccd1 _14600_/X sky130_fd_sc_hd__buf_2
XPHY_4143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11812_ _19452_/Q _11807_/X _09064_/X _11808_/X vssd1 vssd1 vccd1 vccd1 _19452_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15580_ _18588_/Q vssd1 vssd1 vccd1 vccd1 _15581_/B sky130_fd_sc_hd__inv_2
XFILLER_61_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12792_ _18827_/Q vssd1 vssd1 vccd1 vccd1 _13550_/A sky130_fd_sc_hd__inv_2
XPHY_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14531_ _14745_/A vssd1 vssd1 vccd1 vccd1 _14531_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_242_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11743_ _15749_/B _11737_/X _16929_/X _11738_/X vssd1 vssd1 vccd1 vccd1 _19497_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17813__S1 _18750_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17250_ _17249_/X _18904_/Q _17542_/S vssd1 vssd1 vccd1 vccd1 _17250_/X sky130_fd_sc_hd__mux2_1
XPHY_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14462_ _15082_/A _14731_/B _14758_/C vssd1 vssd1 vccd1 vccd1 _14464_/A sky130_fd_sc_hd__or3_4
X_11674_ _11674_/A vssd1 vssd1 vccd1 vccd1 _11674_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_230_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14401__B1 _14326_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16582__B _16583_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16201_ _18771_/Q vssd1 vssd1 vccd1 vccd1 _16201_/Y sky130_fd_sc_hd__inv_2
XPHY_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13413_ _20104_/Q vssd1 vssd1 vccd1 vccd1 _13413_/Y sky130_fd_sc_hd__inv_4
XFILLER_174_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10625_ _18552_/Q vssd1 vssd1 vccd1 vccd1 _10625_/Y sky130_fd_sc_hd__inv_2
XFILLER_155_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15479__A _15479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17181_ _17180_/X _13071_/A _17542_/S vssd1 vssd1 vccd1 vccd1 _17181_/X sky130_fd_sc_hd__mux2_1
X_14393_ _15082_/A _14731_/B _14975_/C vssd1 vssd1 vccd1 vccd1 _14395_/A sky130_fd_sc_hd__or3_4
XFILLER_128_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16132_ _19524_/Q vssd1 vssd1 vccd1 vccd1 _16132_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11800__A _11800_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10556_ _19810_/Q _19809_/Q _10939_/C vssd1 vssd1 vccd1 vccd1 _10559_/C sky130_fd_sc_hd__or3_1
X_13344_ _13428_/B _13344_/B vssd1 vssd1 vccd1 vccd1 _13447_/A sky130_fd_sc_hd__or2_1
XFILLER_185_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14165__C1 _14164_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16063_ _16061_/Y _16053_/X _16062_/Y _16055_/X vssd1 vssd1 vccd1 vccd1 _16063_/X
+ sky130_fd_sc_hd__o22a_1
X_10487_ _19536_/Q _19535_/Q _19534_/Q _19533_/Q vssd1 vssd1 vccd1 vccd1 _10511_/A
+ sky130_fd_sc_hd__or4_4
XANTENNA__16802__S _17385_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13275_ _13293_/B vssd1 vssd1 vccd1 vccd1 _14392_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__14704__B2 _14701_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15014_ _18048_/Q _15010_/X _14996_/X _15012_/X vssd1 vssd1 vccd1 vccd1 _18048_/D
+ sky130_fd_sc_hd__a22o_1
X_12226_ _19235_/Q _12219_/X _12225_/X _12220_/X vssd1 vssd1 vccd1 vccd1 _19235_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_151_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19035__RESET_B repeater267/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19822_ _19822_/CLK _19822_/D repeater227/X vssd1 vssd1 vccd1 vccd1 _19822_/Q sky130_fd_sc_hd__dfrtp_4
X_12157_ _12171_/A vssd1 vssd1 vccd1 vccd1 _12157_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11108_ _19635_/Q _11119_/B vssd1 vssd1 vccd1 vccd1 _11108_/Y sky130_fd_sc_hd__nand2_1
XFILLER_111_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16965_ _16672_/Y _15544_/Y _17474_/S vssd1 vssd1 vccd1 vccd1 _16965_/X sky130_fd_sc_hd__mux2_1
X_12088_ hold306/X vssd1 vssd1 vccd1 vccd1 _12088_/X sky130_fd_sc_hd__clkbuf_4
X_19753_ _19900_/CLK _19753_/D repeater196/X vssd1 vssd1 vccd1 vccd1 _19753_/Q sky130_fd_sc_hd__dfrtp_1
X_11039_ _11039_/A _11039_/B vssd1 vssd1 vccd1 vccd1 _11040_/A sky130_fd_sc_hd__or2_1
X_18704_ _19224_/CLK _18704_/D repeater253/X vssd1 vssd1 vccd1 vccd1 _18704_/Q sky130_fd_sc_hd__dfrtp_4
X_15916_ _17545_/X _16683_/A _15913_/Y _15915_/X vssd1 vssd1 vccd1 vccd1 _15916_/X
+ sky130_fd_sc_hd__o22a_1
X_19684_ _19780_/CLK _19684_/D repeater227/X vssd1 vssd1 vccd1 vccd1 _19684_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_37_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16896_ _16895_/X _15692_/Y _17474_/S vssd1 vssd1 vccd1 vccd1 _16896_/X sky130_fd_sc_hd__mux2_1
X_18635_ _19780_/CLK _18635_/D repeater227/X vssd1 vssd1 vccd1 vccd1 _18635_/Q sky130_fd_sc_hd__dfstp_2
X_15847_ _15833_/X _15844_/X _15846_/X vssd1 vssd1 vccd1 vccd1 _15847_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA_clkbuf_leaf_123_HCLK_A clkbuf_4_4_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18566_ _19841_/CLK _18566_/D repeater271/X vssd1 vssd1 vccd1 vccd1 _18566_/Q sky130_fd_sc_hd__dfrtp_1
X_15778_ _19971_/Q _19328_/Q vssd1 vssd1 vccd1 vccd1 _15778_/X sky130_fd_sc_hd__and2_2
XFILLER_91_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17517_ _17516_/X _15876_/Y _17517_/S vssd1 vssd1 vccd1 vccd1 _17517_/X sky130_fd_sc_hd__mux2_1
X_14729_ _18211_/Q _14718_/A _14691_/X _14719_/A vssd1 vssd1 vccd1 vccd1 _18211_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_178_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18497_ _19794_/CLK _18497_/D repeater203/X vssd1 vssd1 vccd1 vccd1 _18497_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17804__S1 _18752_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12078__A hold279/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17448_ _17447_/X _09467_/A _17530_/S vssd1 vssd1 vccd1 vccd1 _17448_/X sky130_fd_sc_hd__mux2_2
XFILLER_33_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_7_HCLK clkbuf_4_2_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _18959_/CLK sky130_fd_sc_hd__clkbuf_16
X_17379_ _16217_/Y _15594_/A _17474_/S vssd1 vssd1 vccd1 vccd1 _17379_/X sky130_fd_sc_hd__mux2_2
XFILLER_20_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19118_ _19119_/CLK _19118_/D hold353/X vssd1 vssd1 vccd1 vccd1 _19118_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_192_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16696__A1 _16971_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19049_ _19576_/CLK _19049_/D repeater255/X vssd1 vssd1 vccd1 vccd1 _19049_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_118_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12706__B1 _12543_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16448__A1 _15205_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14459__B1 _14419_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17543__S _17543_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18758__RESET_B repeater195/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09704_ _09788_/A _19405_/Q _09629_/A _19429_/Q vssd1 vssd1 vccd1 vccd1 _09704_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12485__A2 _12457_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19335__CLK _20013_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16667__B _16668_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11693__B1 _10877_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09635_ _09635_/A _09635_/B _09807_/C vssd1 vssd1 vccd1 vccd1 _09787_/C sky130_fd_sc_hd__or3_1
XFILLER_231_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09566_ _09607_/A vssd1 vssd1 vccd1 vccd1 _09585_/A sky130_fd_sc_hd__inv_1
XFILLER_71_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_45_HCLK_A clkbuf_opt_2_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19485__CLK _19510_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09497_ _19303_/Q vssd1 vssd1 vccd1 vccd1 _09497_/Y sky130_fd_sc_hd__inv_2
XPHY_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16683__A _16683_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19546__RESET_B hold346/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10410_ _10410_/A vssd1 vssd1 vccd1 vccd1 _14680_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_99_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11390_ _19559_/Q vssd1 vssd1 vccd1 vccd1 _11572_/A sky130_fd_sc_hd__inv_2
XFILLER_164_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17884__A0 _17880_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17718__S _18546_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10341_ _19865_/Q _10341_/B vssd1 vssd1 vccd1 vccd1 _10341_/X sky130_fd_sc_hd__or2_1
XANTENNA__14147__C1 _14106_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13060_ _13060_/A _13060_/B vssd1 vssd1 vccd1 vccd1 _13061_/B sky130_fd_sc_hd__or2_2
XFILLER_136_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10272_ _10266_/B _14316_/B _19645_/Q _19641_/Q vssd1 vssd1 vccd1 vccd1 _11150_/B
+ sky130_fd_sc_hd__a22o_1
X_12011_ _19357_/Q _12009_/X _09030_/X _12010_/X vssd1 vssd1 vccd1 vccd1 _19357_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12451__A _12458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18499__RESET_B repeater219/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17453__S _17487_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16750_ _16750_/A _16750_/B vssd1 vssd1 vccd1 vccd1 _16750_/Y sky130_fd_sc_hd__nor2_8
X_13962_ _13962_/A vssd1 vssd1 vccd1 vccd1 _13966_/A sky130_fd_sc_hd__inv_2
XFILLER_235_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15701_ _18618_/Q _15697_/A _15700_/Y _15697_/Y vssd1 vssd1 vccd1 vccd1 _15702_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_47_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12913_ _19269_/Q vssd1 vssd1 vccd1 vccd1 _12913_/Y sky130_fd_sc_hd__inv_4
X_16681_ _19050_/Q vssd1 vssd1 vccd1 vccd1 _16681_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13893_ _19195_/Q _13802_/B _19222_/Q _13831_/A _13892_/X vssd1 vssd1 vccd1 vccd1
+ _13897_/C sky130_fd_sc_hd__o221a_1
XFILLER_246_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18420_ _18795_/CLK _18420_/D vssd1 vssd1 vccd1 vccd1 _18420_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16072__C1 _16071_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15632_ _18602_/Q vssd1 vssd1 vccd1 vccd1 _15632_/Y sky130_fd_sc_hd__inv_2
X_12844_ _18940_/Q vssd1 vssd1 vccd1 vccd1 _12964_/A sky130_fd_sc_hd__inv_2
XFILLER_221_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18351_ _18959_/CLK _18351_/D vssd1 vssd1 vccd1 vccd1 _18351_/Q sky130_fd_sc_hd__dfxtp_1
X_15563_ _18584_/Q _15562_/A _15561_/Y _15562_/Y vssd1 vssd1 vccd1 vccd1 _15564_/B
+ sky130_fd_sc_hd__o22a_1
X_12775_ _19255_/Q _13555_/A _12774_/Y _18832_/Q vssd1 vssd1 vccd1 vccd1 _12775_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17798__S0 _17923_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17302_ _17486_/A0 _09924_/Y _17522_/S vssd1 vssd1 vccd1 vccd1 _17302_/X sky130_fd_sc_hd__mux2_1
XPHY_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14514_ _18332_/Q _14504_/A _14513_/X _14505_/A vssd1 vssd1 vccd1 vccd1 _18332_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18282_ _19873_/CLK _18282_/D vssd1 vssd1 vccd1 vccd1 _18282_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11726_ _19509_/Q _11723_/X _16941_/X _11724_/X vssd1 vssd1 vccd1 vccd1 hold223/A
+ sky130_fd_sc_hd__a22o_1
XPHY_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15494_ _15571_/A vssd1 vssd1 vccd1 vccd1 _15535_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__19978__CLK _19992_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17233_ _17232_/X _11393_/Y _17545_/S vssd1 vssd1 vccd1 vccd1 _17233_/X sky130_fd_sc_hd__mux2_1
XFILLER_80_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14445_ _18374_/Q _14436_/X _14415_/X _14439_/X vssd1 vssd1 vccd1 vccd1 _18374_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11657_ _10736_/X _11672_/B _11656_/X _18546_/Q _18520_/Q vssd1 vssd1 vccd1 vccd1
+ _11661_/A sky130_fd_sc_hd__o32a_1
XPHY_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11739__A1 _19500_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11739__B2 _11738_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10608_ _10608_/A vssd1 vssd1 vccd1 vccd1 _10609_/A sky130_fd_sc_hd__inv_2
X_17164_ _15963_/X _12761_/Y _17534_/S vssd1 vssd1 vccd1 vccd1 _17164_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14376_ _18411_/Q _14368_/A _14312_/X _14369_/A vssd1 vssd1 vccd1 vccd1 _18411_/D
+ sky130_fd_sc_hd__a22o_1
X_11588_ _11588_/A vssd1 vssd1 vccd1 vccd1 _11588_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_183_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14138__C1 _14106_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16115_ _16115_/A vssd1 vssd1 vccd1 vccd1 _16433_/B sky130_fd_sc_hd__buf_1
XANTENNA__09000__A _19498_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13327_ _13327_/A vssd1 vssd1 vccd1 vccd1 _13483_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_183_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10539_ _18482_/Q vssd1 vssd1 vccd1 vccd1 _10933_/A sky130_fd_sc_hd__inv_2
XFILLER_170_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10146__A hold322/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17095_ _17094_/X _13838_/Y _17545_/S vssd1 vssd1 vccd1 vccd1 _17095_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16046_ _16436_/B _18739_/Q vssd1 vssd1 vccd1 vccd1 _16046_/X sky130_fd_sc_hd__and2_1
X_13258_ _18749_/Q vssd1 vssd1 vccd1 vccd1 _13259_/B sky130_fd_sc_hd__inv_2
XFILLER_170_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12209_ _19246_/Q _12205_/X _12100_/X _12206_/X vssd1 vssd1 vccd1 vccd1 _19246_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_69_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13189_ _13075_/A _13189_/A2 _13187_/Y _13182_/X vssd1 vssd1 vccd1 vccd1 _18903_/D
+ sky130_fd_sc_hd__a211oi_4
XFILLER_123_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19805_ _19813_/CLK _19805_/D repeater224/X vssd1 vssd1 vccd1 vccd1 _19805_/Q sky130_fd_sc_hd__dfrtp_1
X_17997_ _19849_/CLK _17997_/D vssd1 vssd1 vccd1 vccd1 _17997_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__18851__RESET_B repeater232/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17363__S _17546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19736_ _20055_/CLK _19736_/D repeater208/X vssd1 vssd1 vccd1 vccd1 _19736_/Q sky130_fd_sc_hd__dfrtp_1
X_16948_ _19492_/Q hold130/X _16950_/S vssd1 vssd1 vccd1 vccd1 _16948_/X sky130_fd_sc_hd__mux2_1
XFILLER_238_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16879_ _15963_/X _09560_/Y _17534_/S vssd1 vssd1 vccd1 vccd1 _16879_/X sky130_fd_sc_hd__mux2_1
X_19667_ _19667_/CLK _19667_/D repeater270/X vssd1 vssd1 vccd1 vccd1 _19667_/Q sky130_fd_sc_hd__dfrtp_1
X_09420_ _19391_/Q vssd1 vssd1 vccd1 vccd1 _09420_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18618_ _19577_/CLK _18618_/D repeater269/X vssd1 vssd1 vccd1 vccd1 _18618_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_213_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19598_ _19600_/CLK _19598_/D hold273/X vssd1 vssd1 vccd1 vccd1 _19598_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_241_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09351_ _20026_/Q vssd1 vssd1 vccd1 vccd1 _09486_/A sky130_fd_sc_hd__inv_6
X_18549_ _18633_/CLK _18549_/D repeater229/X vssd1 vssd1 vccd1 vccd1 _18549_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_178_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17789__S0 _19647_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_221_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09282_ _10429_/A vssd1 vssd1 vccd1 vccd1 _14245_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_178_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12536__A hold331/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_108_HCLK clkbuf_4_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19221_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__17538__S _17548_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10705__A2 _10704_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11902__A1 _19415_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08997_ _19519_/Q _18624_/Q vssd1 vssd1 vccd1 vccd1 _13280_/A sky130_fd_sc_hd__nand2_2
XFILLER_102_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13104__B1 _19172_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17273__S _17546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_hold175_A HADDR[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14852__B1 _14812_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09618_ _09618_/A vssd1 vssd1 vccd1 vccd1 _09618_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_hold342_A MSI_S2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_243_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13407__A1 _20108_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10890_ _19694_/Q _10878_/A _10868_/X _10879_/A vssd1 vssd1 vccd1 vccd1 _19694_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19798__RESET_B repeater222/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09549_ _20016_/Q _09547_/Y _20024_/Q _16620_/A vssd1 vssd1 vccd1 vccd1 _09549_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13252__D _13252_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19727__RESET_B repeater205/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12091__B1 _12090_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12560_ _12576_/A vssd1 vssd1 vccd1 vccd1 _12560_/X sky130_fd_sc_hd__buf_1
XPHY_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11511_ _11511_/A vssd1 vssd1 vccd1 vccd1 _11511_/Y sky130_fd_sc_hd__inv_2
XPHY_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12491_ _12529_/A vssd1 vssd1 vccd1 vccd1 _12506_/A sky130_fd_sc_hd__clkbuf_2
XPHY_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19380__RESET_B repeater230/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14230_ _18500_/Q _14230_/B vssd1 vssd1 vccd1 vccd1 _14231_/B sky130_fd_sc_hd__or2_1
XFILLER_11_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11442_ _11548_/A _19129_/Q _11577_/A _19144_/Q vssd1 vssd1 vccd1 vccd1 _11442_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_11_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17448__S _17530_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11373_ _19572_/Q vssd1 vssd1 vccd1 vccd1 _11584_/C sky130_fd_sc_hd__inv_2
X_14161_ _14160_/Y _18682_/Q _19103_/Q _14012_/A vssd1 vssd1 vccd1 vccd1 _14161_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_109_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10324_ _10324_/A _10366_/A vssd1 vssd1 vccd1 vccd1 _10364_/B sky130_fd_sc_hd__nor2_1
X_13112_ _19171_/Q _18900_/Q _13111_/Y _13072_/A vssd1 vssd1 vccd1 vccd1 _13112_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_152_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14092_ _14090_/Y _18673_/Q _19077_/Q _14018_/A _14091_/X vssd1 vssd1 vccd1 vccd1
+ _14093_/D sky130_fd_sc_hd__o221a_1
XFILLER_98_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17920_ _18321_/Q _18441_/Q _18433_/Q _18425_/Q _17923_/S0 _19646_/Q vssd1 vssd1
+ vccd1 vccd1 _17920_/X sky130_fd_sc_hd__mux4_1
X_10255_ _15823_/A _10410_/A vssd1 vssd1 vccd1 vccd1 _15190_/A sky130_fd_sc_hd__or2_4
X_13043_ _18903_/Q vssd1 vssd1 vccd1 vccd1 _13075_/A sky130_fd_sc_hd__inv_2
XANTENNA__10157__B1 _09082_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12181__A _12187_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17851_ _16332_/Y _16333_/Y _16334_/Y _16335_/Y _17913_/S0 _19632_/Q vssd1 vssd1
+ vccd1 vccd1 _17851_/X sky130_fd_sc_hd__mux4_2
XFILLER_78_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10186_ _10186_/A _10186_/B _15749_/C vssd1 vssd1 vccd1 vccd1 _10188_/S sky130_fd_sc_hd__or3_4
XFILLER_120_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16802_ _16801_/X _16707_/Y _17385_/S vssd1 vssd1 vccd1 vccd1 _16802_/X sky130_fd_sc_hd__mux2_1
XANTENNA__17183__S _17490_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17782_ _18325_/Q _18005_/Q _18309_/Q _18301_/Q _17923_/S0 _19646_/Q vssd1 vssd1
+ vccd1 vccd1 _17782_/X sky130_fd_sc_hd__mux4_2
X_14994_ _14994_/A vssd1 vssd1 vccd1 vccd1 _14994_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19521_ _20049_/CLK _19521_/D repeater190/X vssd1 vssd1 vccd1 vccd1 _19521_/Q sky130_fd_sc_hd__dfstp_1
X_16733_ _16784_/X _16513_/A _16786_/X _16002_/X vssd1 vssd1 vccd1 vccd1 _16733_/X
+ sky130_fd_sc_hd__o22a_1
X_13945_ _13945_/A _13962_/A vssd1 vssd1 vccd1 vccd1 _13960_/A sky130_fd_sc_hd__or2_1
XFILLER_207_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19452_ _19841_/CLK _19452_/D repeater272/X vssd1 vssd1 vccd1 vccd1 _19452_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_90_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16664_ _16572_/X _16664_/B _16664_/C vssd1 vssd1 vccd1 vccd1 _16664_/Y sky130_fd_sc_hd__nand3b_2
X_13876_ _19205_/Q _13909_/D _19198_/Q _13946_/A vssd1 vssd1 vccd1 vccd1 _13876_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_201_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15615_ _15618_/B _15613_/X _15614_/X vssd1 vssd1 vccd1 vccd1 _15615_/X sky130_fd_sc_hd__o21a_1
X_18403_ _18954_/CLK _18403_/D vssd1 vssd1 vccd1 vccd1 _18403_/Q sky130_fd_sc_hd__dfxtp_1
X_19383_ _19927_/CLK _19383_/D repeater235/X vssd1 vssd1 vccd1 vccd1 _19383_/Q sky130_fd_sc_hd__dfrtp_2
X_12827_ _19228_/Q vssd1 vssd1 vccd1 vccd1 _12827_/Y sky130_fd_sc_hd__inv_2
XANTENNA__10880__A1 _15364_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16595_ _16595_/A vssd1 vssd1 vccd1 vccd1 _16595_/X sky130_fd_sc_hd__buf_1
XFILLER_61_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19468__RESET_B repeater274/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18334_ _19849_/CLK _18334_/D vssd1 vssd1 vccd1 vccd1 _18334_/Q sky130_fd_sc_hd__dfxtp_1
X_15546_ _15550_/B vssd1 vssd1 vccd1 vccd1 _15552_/B sky130_fd_sc_hd__inv_2
XFILLER_188_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12758_ _12758_/A _12758_/B _12758_/C _12758_/D vssd1 vssd1 vccd1 vccd1 _12834_/A
+ sky130_fd_sc_hd__and4_1
XPHY_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10093__C1 _10107_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11709_ _11737_/A vssd1 vssd1 vccd1 vccd1 _11738_/A sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_91_HCLK_A clkbuf_4_12_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18265_ _20077_/CLK _18265_/D vssd1 vssd1 vccd1 vccd1 _18265_/Q sky130_fd_sc_hd__dfxtp_1
X_15477_ _18564_/Q vssd1 vssd1 vccd1 vccd1 _15477_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12356__A hold251/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12689_ _18973_/Q _12684_/X _12030_/A _12685_/X vssd1 vssd1 vccd1 vccd1 _18973_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17216_ _17486_/A0 _13149_/Y _17543_/S vssd1 vssd1 vccd1 vccd1 _17216_/X sky130_fd_sc_hd__mux2_1
X_14428_ _18384_/Q _14424_/X _14356_/X _14426_/X vssd1 vssd1 vccd1 vccd1 _18384_/D
+ sky130_fd_sc_hd__a22o_1
X_18196_ _18333_/CLK _18196_/D vssd1 vssd1 vccd1 vccd1 _18196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17358__S _17529_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09786__C1 _09813_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17147_ _17486_/A0 _09930_/Y _17543_/S vssd1 vssd1 vccd1 vccd1 _17147_/X sky130_fd_sc_hd__mux2_1
XFILLER_143_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14359_ _14751_/A vssd1 vssd1 vccd1 vccd1 _14359_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17078_ _17077_/X _12925_/Y _17487_/S vssd1 vssd1 vccd1 vccd1 _17078_/X sky130_fd_sc_hd__mux2_1
XFILLER_143_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08920_ _19853_/Q vssd1 vssd1 vccd1 vccd1 _10321_/A sky130_fd_sc_hd__inv_2
X_16029_ _17971_/Q vssd1 vssd1 vccd1 vccd1 _16029_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_226_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10699__A1 _10698_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11896__B1 _09049_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15087__B1 hold236/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17093__S _17546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19719_ _20049_/CLK _19719_/D repeater190/X vssd1 vssd1 vccd1 vccd1 _19719_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_84_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19891__RESET_B repeater207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_240_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09403_ _19914_/Q vssd1 vssd1 vccd1 vccd1 _10086_/A sky130_fd_sc_hd__inv_2
XFILLER_25_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09334_ _19735_/Q _19734_/Q _19736_/Q _19733_/Q _19737_/Q vssd1 vssd1 vccd1 vccd1
+ _10791_/A sky130_fd_sc_hd__a41o_1
XANTENNA__12073__B1 _12069_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19138__RESET_B repeater274/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11820__B1 _10877_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09265_ _09255_/X _20058_/Q _09265_/S vssd1 vssd1 vccd1 vccd1 _20058_/D sky130_fd_sc_hd__mux2_1
XFILLER_178_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18278__CLK _19847_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09196_ _18870_/Q _08919_/A _20123_/Q _17605_/S vssd1 vssd1 vccd1 vccd1 _09197_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__15577__A _15610_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17268__S _17541_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16900__S _17512_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold292_A HWDATA[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10040_ _10040_/A _10040_/B vssd1 vssd1 vccd1 vccd1 _10068_/A sky130_fd_sc_hd__or2_1
XANTENNA__18702__RESET_B hold351/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11887__B1 _09033_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15078__B1 _14793_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16814__A1 _14039_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14825__B1 _14751_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19979__RESET_B repeater192/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11991_ _12313_/A vssd1 vssd1 vccd1 vccd1 _11991_/X sky130_fd_sc_hd__buf_1
XFILLER_152_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17731__S _18508_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19908__RESET_B repeater241/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13730_ _14975_/B vssd1 vssd1 vccd1 vccd1 _14758_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_10942_ _10942_/A _10942_/B _10942_/C vssd1 vssd1 vccd1 vccd1 _15298_/C sky130_fd_sc_hd__or3_1
XFILLER_44_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13661_ _18785_/Q _13656_/X _12030_/A _13658_/X vssd1 vssd1 vccd1 vccd1 _18785_/D
+ sky130_fd_sc_hd__a22o_1
X_10873_ _16053_/A vssd1 vssd1 vccd1 vccd1 _15973_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__19561__RESET_B repeater269/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15400_ _15402_/A _17580_/X vssd1 vssd1 vccd1 vccd1 _18532_/D sky130_fd_sc_hd__and2_1
XFILLER_71_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12612_ _12650_/A vssd1 vssd1 vccd1 vccd1 _12629_/A sky130_fd_sc_hd__clkbuf_2
X_16380_ _19762_/Q vssd1 vssd1 vccd1 vccd1 _16380_/Y sky130_fd_sc_hd__inv_2
XPHY_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13592_ _18817_/Q _13590_/Y _13591_/X _13541_/B vssd1 vssd1 vccd1 vccd1 _18817_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15331_ _18878_/Q vssd1 vssd1 vccd1 vccd1 _15333_/A sky130_fd_sc_hd__inv_2
XFILLER_197_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12543_ _14405_/A vssd1 vssd1 vccd1 vccd1 _12543_/X sky130_fd_sc_hd__buf_6
XANTENNA__11811__B1 _09061_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18050_ _19851_/CLK _18050_/D vssd1 vssd1 vccd1 vccd1 _18050_/Q sky130_fd_sc_hd__dfxtp_1
X_15262_ _15389_/B _15285_/A _18632_/Q _15283_/A _15261_/X vssd1 vssd1 vccd1 vccd1
+ _18632_/D sky130_fd_sc_hd__a32o_1
XFILLER_157_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12474_ _19103_/Q _12471_/X _12356_/X _12472_/X vssd1 vssd1 vccd1 vccd1 _19103_/D
+ sky130_fd_sc_hd__a22o_1
X_17001_ _17000_/X _11341_/Y _17490_/S vssd1 vssd1 vccd1 vccd1 _17001_/X sky130_fd_sc_hd__mux2_1
XANTENNA__16590__B _16622_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13564__B1 _13560_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14213_ _14211_/Y _18702_/Q _14212_/Y _18685_/Q vssd1 vssd1 vccd1 vccd1 _14213_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__17178__S _17542_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11425_ _19156_/Q vssd1 vssd1 vccd1 vccd1 _11425_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15193_ _15193_/A vssd1 vssd1 vccd1 vccd1 _17761_/S sky130_fd_sc_hd__inv_2
XFILLER_137_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14144_ _14007_/A _14144_/A2 _14142_/Y _14106_/X vssd1 vssd1 vccd1 vccd1 _18676_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_125_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11356_ _11463_/A _18964_/Q _11462_/A _18963_/Q vssd1 vssd1 vccd1 vccd1 _11356_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_141_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10307_ _18609_/Q _18608_/Q _18610_/Q vssd1 vssd1 vccd1 vccd1 _15668_/A sky130_fd_sc_hd__or3_1
XFILLER_141_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14075_ _14073_/Y _18697_/Q _14074_/Y _18683_/Q vssd1 vssd1 vccd1 vccd1 _14075_/X
+ sky130_fd_sc_hd__o22a_1
X_18952_ _18954_/CLK _18952_/D repeater257/X vssd1 vssd1 vccd1 vccd1 _18952_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_112_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11287_ _19603_/Q vssd1 vssd1 vccd1 vccd1 _11483_/A sky130_fd_sc_hd__inv_2
XANTENNA__16810__S _17546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17903_ _15931_/Y _15932_/Y _15933_/Y _15934_/Y _17913_/S0 _19632_/Q vssd1 vssd1
+ vccd1 vccd1 _17903_/X sky130_fd_sc_hd__mux4_2
X_13026_ _13021_/A _13021_/B _13021_/C vssd1 vssd1 vccd1 vccd1 _13027_/B sky130_fd_sc_hd__o21a_1
XFILLER_140_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10238_ _10236_/Y _19661_/Q _19834_/Q _10996_/A vssd1 vssd1 vccd1 vccd1 _10238_/X
+ sky130_fd_sc_hd__o22a_1
X_18883_ _19814_/CLK _18883_/D repeater220/X vssd1 vssd1 vccd1 vccd1 _18883_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_239_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15069__B1 _15020_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17834_ _17830_/X _17831_/X _17832_/X _17833_/X _18751_/Q _18752_/Q vssd1 vssd1 vccd1
+ vccd1 _17834_/X sky130_fd_sc_hd__mux4_2
XFILLER_120_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10169_ _19887_/Q _10166_/X _09077_/X _10168_/X vssd1 vssd1 vccd1 vccd1 _19887_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_66_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17765_ _18314_/Q _18434_/Q _18426_/Q _18418_/Q _17923_/S0 _19646_/Q vssd1 vssd1
+ vccd1 vccd1 _17765_/X sky130_fd_sc_hd__mux4_1
X_14977_ hold248/X vssd1 vssd1 vccd1 vccd1 hold247/A sky130_fd_sc_hd__buf_2
XFILLER_207_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrebuffer19 _14024_/B vssd1 vssd1 vccd1 vccd1 _14114_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_81_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19649__RESET_B repeater261/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17641__S _17655_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19504_ _19510_/CLK hold227/X repeater256/X vssd1 vssd1 vccd1 vccd1 _19504_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_35_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16716_ _16716_/A _16718_/B vssd1 vssd1 vccd1 vccd1 _16716_/Y sky130_fd_sc_hd__nor2_1
XFILLER_75_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13928_ _13912_/D _13825_/B _13924_/Y _13927_/X vssd1 vssd1 vccd1 vccd1 _18726_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_235_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17696_ _15446_/Y _19439_/Q _17696_/S vssd1 vssd1 vccd1 vccd1 _18556_/D sky130_fd_sc_hd__mux2_1
XFILLER_222_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17230__A1 _08947_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16647_ _16647_/A _16647_/B vssd1 vssd1 vccd1 vccd1 _16647_/Y sky130_fd_sc_hd__nor2_1
X_19435_ _19435_/CLK _19435_/D repeater259/X vssd1 vssd1 vccd1 vccd1 _19435_/Q sky130_fd_sc_hd__dfrtp_1
X_13859_ _19220_/Q vssd1 vssd1 vccd1 vccd1 _13859_/Y sky130_fd_sc_hd__inv_2
XFILLER_179_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19366_ _19933_/CLK _19366_/D repeater236/X vssd1 vssd1 vccd1 vccd1 _19366_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_34_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16578_ _16688_/A vssd1 vssd1 vccd1 vccd1 _16578_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_188_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18317_ _19637_/CLK _18317_/D vssd1 vssd1 vccd1 vccd1 _18317_/Q sky130_fd_sc_hd__dfxtp_1
X_15529_ _15530_/A vssd1 vssd1 vccd1 vccd1 _15529_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11802__B1 hold314/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19297_ _20013_/CLK _19297_/D repeater241/X vssd1 vssd1 vccd1 vccd1 _19297_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_175_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12086__A hold308/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09050_ _20109_/Q _09041_/X _09049_/X _09043_/X vssd1 vssd1 vccd1 vccd1 _20109_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_175_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrebuffer109 _14020_/B vssd1 vssd1 vccd1 vccd1 _14124_/B1 sky130_fd_sc_hd__dlygate4sd1_1
X_18248_ _19847_/CLK _18248_/D vssd1 vssd1 vccd1 vccd1 _18248_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17088__S _17493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18179_ _18460_/CLK _18179_/D vssd1 vssd1 vccd1 vccd1 _18179_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17916__S0 _17918_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11030__A1 _11023_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09952_ _09990_/A vssd1 vssd1 vccd1 vccd1 _09987_/B sky130_fd_sc_hd__buf_2
XFILLER_103_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20072_ _20124_/CLK _20072_/D repeater207/X vssd1 vssd1 vccd1 vccd1 _20072_/Q sky130_fd_sc_hd__dfrtp_1
X_09883_ _19349_/Q vssd1 vssd1 vccd1 vccd1 _09883_/Y sky130_fd_sc_hd__inv_2
XFILLER_218_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12294__B1 _12223_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12046__B1 _11981_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09317_ _18655_/Q vssd1 vssd1 vccd1 vccd1 _09317_/X sky130_fd_sc_hd__buf_1
XFILLER_167_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09248_ _20063_/Q _20064_/Q _09250_/S vssd1 vssd1 vccd1 vccd1 _20064_/D sky130_fd_sc_hd__mux2_1
XFILLER_182_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18954__RESET_B repeater257/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09179_ _20076_/Q vssd1 vssd1 vccd1 vccd1 _14711_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_193_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17907__S0 _17908_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11210_ _19608_/Q _11205_/Y _11486_/A _19020_/Q _11209_/X vssd1 vssd1 vccd1 vccd1
+ _11223_/B sky130_fd_sc_hd__o221a_1
X_12190_ _12228_/A vssd1 vssd1 vccd1 vccd1 _12229_/A sky130_fd_sc_hd__inv_2
XFILLER_123_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16496__C1 _16495_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11141_ _15232_/A _19225_/Q _12253_/B _11144_/B vssd1 vssd1 vccd1 vccd1 _11141_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_122_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11072_ _11061_/X _11066_/B _11123_/B vssd1 vssd1 vccd1 vccd1 _11072_/Y sky130_fd_sc_hd__o21ai_1
Xoutput88 _16607_/Y vssd1 vssd1 vccd1 vccd1 HRDATA[18] sky130_fd_sc_hd__clkbuf_2
Xoutput99 _16715_/Y vssd1 vssd1 vccd1 vccd1 HRDATA[28] sky130_fd_sc_hd__clkbuf_2
X_10023_ _10023_/A _10101_/B _10023_/C vssd1 vssd1 vccd1 vccd1 _10024_/A sky130_fd_sc_hd__or3_1
XFILLER_88_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14900_ _18112_/Q _14896_/X _14703_/X _14898_/X vssd1 vssd1 vccd1 vccd1 _18112_/D
+ sky130_fd_sc_hd__a22o_1
X_15880_ _19870_/Q vssd1 vssd1 vccd1 vccd1 _15880_/Y sky130_fd_sc_hd__inv_2
XFILLER_248_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14831_ _15058_/A _15034_/B _15034_/C vssd1 vssd1 vccd1 vccd1 _14833_/A sky130_fd_sc_hd__or3_4
XFILLER_56_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17461__S _19498_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19742__RESET_B repeater207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17550_ _15847_/Y _18663_/Q _17550_/S vssd1 vssd1 vccd1 vccd1 _17550_/X sky130_fd_sc_hd__mux2_1
XFILLER_217_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12285__B1 _12107_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14762_ _18193_/Q _14759_/X _14745_/X _14761_/X vssd1 vssd1 vccd1 vccd1 _18193_/D
+ sky130_fd_sc_hd__a22o_1
X_11974_ _19374_/Q _11969_/X _11911_/X _11970_/X vssd1 vssd1 vccd1 vccd1 _19374_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_16_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16501_ _20101_/Q vssd1 vssd1 vccd1 vccd1 _16501_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16585__B _16615_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_217_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13713_ _17761_/X _13710_/B _13712_/X vssd1 vssd1 vccd1 vccd1 _18759_/D sky130_fd_sc_hd__a21oi_1
X_10925_ _17721_/X _10923_/X _19680_/Q _10924_/X vssd1 vssd1 vccd1 vccd1 _19680_/D
+ sky130_fd_sc_hd__a22o_1
X_17481_ _17480_/X _09446_/Y _17529_/S vssd1 vssd1 vccd1 vccd1 _17481_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14693_ hold321/X vssd1 vssd1 vccd1 vccd1 _14693_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_232_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19220_ _19293_/CLK _19220_/D repeater186/X vssd1 vssd1 vccd1 vccd1 _19220_/Q sky130_fd_sc_hd__dfrtp_4
X_16432_ _18113_/Q vssd1 vssd1 vccd1 vccd1 _16432_/Y sky130_fd_sc_hd__inv_2
X_13644_ _13644_/A vssd1 vssd1 vccd1 vccd1 _13644_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__12037__B1 _12035_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10856_ _10856_/A vssd1 vssd1 vccd1 vccd1 _10857_/A sky130_fd_sc_hd__inv_2
XFILLER_220_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19151_ _19576_/CLK _19151_/D repeater255/X vssd1 vssd1 vccd1 vccd1 _19151_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16363_ _17943_/Q _16483_/B vssd1 vssd1 vccd1 vccd1 _16363_/X sky130_fd_sc_hd__and2_1
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13575_ _18827_/Q _13573_/Y _13574_/X _13575_/C1 vssd1 vssd1 vccd1 vccd1 _18827_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA_repeater162_A _17473_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16805__S _17487_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10787_ _19740_/Q _10786_/B _10793_/B _10786_/Y vssd1 vssd1 vccd1 vccd1 _19740_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18102_ _18137_/CLK _18102_/D vssd1 vssd1 vccd1 vccd1 _18102_/Q sky130_fd_sc_hd__dfxtp_1
X_15314_ _15243_/Y _15313_/X _15312_/Y _15306_/X _15266_/X vssd1 vssd1 vccd1 vccd1
+ _18625_/D sky130_fd_sc_hd__o221ai_1
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19082_ _19115_/CLK _19082_/D hold353/X vssd1 vssd1 vccd1 vccd1 _19082_/Q sky130_fd_sc_hd__dfrtp_2
X_12526_ _19069_/Q _12519_/X hold259/X _12520_/X vssd1 vssd1 vccd1 vccd1 _19069_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_158_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16294_ _18803_/Q _16114_/Y _16292_/X _16293_/X _16199_/Y vssd1 vssd1 vccd1 vccd1
+ _16294_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_173_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18033_ _18145_/CLK _18033_/D vssd1 vssd1 vccd1 vccd1 _18033_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__18695__RESET_B hold351/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15245_ _15289_/A _15259_/A _15263_/A vssd1 vssd1 vccd1 vccd1 _15245_/X sky130_fd_sc_hd__or3_4
X_12457_ _12457_/A vssd1 vssd1 vccd1 vccd1 _12457_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_output91_A _16629_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11408_ _19157_/Q vssd1 vssd1 vccd1 vccd1 _11408_/Y sky130_fd_sc_hd__inv_2
X_15176_ _17941_/Q _15170_/X _10698_/X _15172_/X vssd1 vssd1 vccd1 vccd1 _17941_/D
+ sky130_fd_sc_hd__a22o_1
X_12388_ _12400_/A vssd1 vssd1 vccd1 vccd1 _12388_/X sky130_fd_sc_hd__buf_1
XFILLER_141_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14127_ _18687_/Q _14126_/Y _14116_/X _14018_/B vssd1 vssd1 vccd1 vccd1 _18687_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_141_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11339_ _19601_/Q _11338_/Y _11470_/A _18972_/Q vssd1 vssd1 vccd1 vccd1 _11339_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_207_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19984_ _19984_/CLK _19984_/D repeater193/X vssd1 vssd1 vccd1 vccd1 _19984_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__10154__A _10155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18935_ _19315_/CLK _18935_/D repeater214/X vssd1 vssd1 vccd1 vccd1 _18935_/Q sky130_fd_sc_hd__dfrtp_1
X_14058_ _19089_/Q _14030_/A _14057_/Y _18700_/Q vssd1 vssd1 vccd1 vccd1 _14058_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_97_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13009_ _18930_/Q _13008_/Y _12980_/A _12873_/B vssd1 vssd1 vccd1 vccd1 _18930_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_228_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18866_ _18866_/CLK _18866_/D repeater232/X vssd1 vssd1 vccd1 vccd1 _18866_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_95_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17817_ _18357_/Q _17997_/Q _18413_/Q _18397_/Q _17918_/S0 _18750_/Q vssd1 vssd1
+ vccd1 vccd1 _17817_/X sky130_fd_sc_hd__mux4_2
X_18797_ _19435_/CLK _18797_/D repeater258/X vssd1 vssd1 vccd1 vccd1 _18797_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__19483__RESET_B repeater260/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17371__S _17566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17748_ _15318_/Y _11093_/Y _17754_/S vssd1 vssd1 vccd1 vccd1 _17748_/X sky130_fd_sc_hd__mux2_1
XFILLER_63_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19412__RESET_B repeater244/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10826__A1 _10451_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17679_ _15516_/Y _19456_/Q _17683_/S vssd1 vssd1 vccd1 vccd1 _18573_/D sky130_fd_sc_hd__mux2_1
XFILLER_50_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19418_ _19997_/CLK _19418_/D repeater271/X vssd1 vssd1 vccd1 vccd1 _19418_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_22_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19349_ _19352_/CLK _19349_/D hold373/X vssd1 vssd1 vccd1 vccd1 _19349_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__09444__B2 _19380_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09102_ _20093_/Q _09084_/X _09101_/X _09087_/X vssd1 vssd1 vccd1 vccd1 _20093_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_149_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09033_ hold308/X vssd1 vssd1 vccd1 vccd1 _09033_/X sky130_fd_sc_hd__buf_4
XFILLER_248_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12200__B1 _12083_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold310 input47/X vssd1 vssd1 vccd1 vccd1 hold310/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold321 hold321/A vssd1 vssd1 vccd1 vccd1 hold321/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold332 input63/X vssd1 vssd1 vccd1 vccd1 hold332/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold343 hold362/X vssd1 vssd1 vccd1 vccd1 hold343/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17546__S _17546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold354 hold354/A vssd1 vssd1 vccd1 vccd1 hold354/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold365 hold365/A vssd1 vssd1 vccd1 vccd1 hold365/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20124_ _20124_/CLK _20124_/D repeater196/X vssd1 vssd1 vccd1 vccd1 _20124_/Q sky130_fd_sc_hd__dfrtp_1
X_09935_ _19358_/Q vssd1 vssd1 vccd1 vccd1 _09935_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12503__A1 _19084_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20055_ _20055_/CLK _20055_/D repeater204/X vssd1 vssd1 vccd1 vccd1 _20055_/Q sky130_fd_sc_hd__dfrtp_1
X_09866_ _09866_/A _09972_/A vssd1 vssd1 vccd1 vccd1 _09867_/B sky130_fd_sc_hd__or2_1
XFILLER_112_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09797_ _09797_/A vssd1 vssd1 vccd1 vccd1 _09797_/Y sky130_fd_sc_hd__inv_2
Xrepeater160 _17493_/S vssd1 vssd1 vccd1 vccd1 _17490_/S sky130_fd_sc_hd__buf_8
XFILLER_234_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17281__S _17385_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater171 _17482_/S vssd1 vssd1 vccd1 vccd1 _17386_/S sky130_fd_sc_hd__buf_8
XANTENNA__15590__A _15643_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater182 _19631_/Q vssd1 vssd1 vccd1 vccd1 _17913_/S0 sky130_fd_sc_hd__clkbuf_16
XPHY_4314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12267__B1 _12078_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater193 repeater198/X vssd1 vssd1 vccd1 vccd1 repeater193/X sky130_fd_sc_hd__buf_8
XPHY_4336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10710_ _10710_/A vssd1 vssd1 vccd1 vccd1 _19775_/D sky130_fd_sc_hd__inv_2
XANTENNA__12019__B1 hold300/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_242_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11690_ _11691_/A vssd1 vssd1 vccd1 vccd1 _11690_/X sky130_fd_sc_hd__clkbuf_2
XPHY_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10641_ _18509_/Q vssd1 vssd1 vccd1 vccd1 _10660_/A sky130_fd_sc_hd__inv_2
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13360_ _13357_/Y _18868_/Q _20122_/Q _13356_/Y _13359_/X vssd1 vssd1 vccd1 vccd1
+ _13360_/X sky130_fd_sc_hd__a221o_1
X_10572_ _19813_/Q _10572_/B _10572_/C vssd1 vssd1 vccd1 vccd1 _10574_/A sky130_fd_sc_hd__or3_4
XFILLER_220_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15749__B _15749_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12311_ _15776_/A _12316_/B vssd1 vssd1 vccd1 vccd1 _12312_/S sky130_fd_sc_hd__or2_1
XFILLER_158_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13291_ _14392_/A vssd1 vssd1 vccd1 vccd1 _13291_/Y sky130_fd_sc_hd__inv_2
XFILLER_182_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15030_ _18037_/Q _15023_/X _15002_/X _15025_/X vssd1 vssd1 vccd1 vccd1 _18037_/D
+ sky130_fd_sc_hd__a22o_1
X_12242_ _19227_/Q _12205_/A _12241_/X _12206_/A vssd1 vssd1 vccd1 vccd1 _19227_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__15765__A _19764_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17456__S _17544_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12173_ _19268_/Q _12171_/X _11978_/X _12172_/X vssd1 vssd1 vccd1 vccd1 _19268_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18809__CLK _20115_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19994__RESET_B repeater192/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11124_ _11124_/A vssd1 vssd1 vccd1 vccd1 _11127_/A sky130_fd_sc_hd__inv_2
X_16981_ _17809_/X _19899_/Q _16986_/S vssd1 vssd1 vccd1 vccd1 _16981_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19923__RESET_B repeater230/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18720_ _18727_/CLK _18720_/D repeater253/X vssd1 vssd1 vccd1 vccd1 _18720_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__13285__A _13285_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11055_ _14317_/B _11049_/Y _11053_/X vssd1 vssd1 vccd1 vccd1 _19643_/D sky130_fd_sc_hd__o21a_1
X_15932_ _18403_/Q vssd1 vssd1 vccd1 vccd1 _15932_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10702__A hold264/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10006_ _19327_/Q vssd1 vssd1 vccd1 vccd1 _10081_/B sky130_fd_sc_hd__inv_2
XFILLER_37_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17433__A1 _17879_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15863_ _19125_/Q _15863_/B vssd1 vssd1 vccd1 vccd1 _15863_/Y sky130_fd_sc_hd__nor2_1
XFILLER_77_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18651_ _20050_/CLK _18651_/D repeater206/X vssd1 vssd1 vccd1 vccd1 _18651_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_92_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17191__S _17546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17602_ _15322_/X _15321_/Y _17605_/S vssd1 vssd1 vccd1 vccd1 _17602_/X sky130_fd_sc_hd__mux2_1
X_14814_ _14814_/A vssd1 vssd1 vccd1 vccd1 _14814_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_64_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18582_ _19470_/CLK _18582_/D repeater273/X vssd1 vssd1 vccd1 vccd1 _18582_/Q sky130_fd_sc_hd__dfrtp_1
X_15794_ _18338_/Q vssd1 vssd1 vccd1 vccd1 _15794_/Y sky130_fd_sc_hd__inv_2
X_17533_ _17532_/X _15870_/Y _17539_/S vssd1 vssd1 vccd1 vccd1 _17533_/X sky130_fd_sc_hd__mux2_1
XANTENNA__17197__A0 _15768_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14745_ _14745_/A vssd1 vssd1 vccd1 vccd1 _14745_/X sky130_fd_sc_hd__buf_2
X_11957_ _19387_/Q _11955_/X hold314/X _11956_/X vssd1 vssd1 vccd1 vccd1 _19387_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_33_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10908_ _10908_/A vssd1 vssd1 vccd1 vccd1 _10908_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17464_ _17463_/X _16042_/Y _17565_/S vssd1 vssd1 vccd1 vccd1 _17464_/X sky130_fd_sc_hd__mux2_1
X_14676_ _18237_/Q _14669_/X _09180_/X _14671_/X vssd1 vssd1 vccd1 vccd1 _18237_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_220_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11888_ _19425_/Q _11884_/X hold305/X _11885_/X vssd1 vssd1 vccd1 vccd1 _19425_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_199_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16415_ _17316_/X _16415_/B vssd1 vssd1 vccd1 vccd1 _16415_/X sky130_fd_sc_hd__and2_1
X_19203_ _19208_/CLK _19203_/D hold367/X vssd1 vssd1 vccd1 vccd1 _19203_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18876__RESET_B repeater208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13627_ _18801_/Q _13499_/X _13620_/B _13626_/X vssd1 vssd1 vccd1 vccd1 _18801_/D
+ sky130_fd_sc_hd__a31o_1
X_10839_ _10839_/A vssd1 vssd1 vccd1 vccd1 _19718_/D sky130_fd_sc_hd__inv_2
X_17395_ _16203_/Y _16202_/Y _17564_/S vssd1 vssd1 vccd1 vccd1 _17395_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10149__A _12370_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18805__RESET_B repeater231/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16346_ _17345_/X _16435_/B vssd1 vssd1 vccd1 vccd1 _16346_/Y sky130_fd_sc_hd__nand2_1
X_19134_ _19137_/CLK _19134_/D repeater249/X vssd1 vssd1 vccd1 vccd1 _19134_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_192_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13558_ _13558_/A vssd1 vssd1 vccd1 vccd1 _13558_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12430__B1 _12302_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12509_ _19080_/Q _12505_/X _12406_/X _12506_/X vssd1 vssd1 vccd1 vccd1 _19080_/D
+ sky130_fd_sc_hd__a22o_1
X_19065_ _19585_/CLK _19065_/D hold363/X vssd1 vssd1 vccd1 vccd1 _19065_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_172_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16277_ _17950_/Q vssd1 vssd1 vccd1 vccd1 _16277_/Y sky130_fd_sc_hd__inv_2
X_13489_ _13489_/A _13489_/B _13489_/C vssd1 vssd1 vccd1 vccd1 _18838_/D sky130_fd_sc_hd__nor3_1
XFILLER_157_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15228_ _15219_/Y _15226_/Y _15227_/Y _18513_/Q vssd1 vssd1 vccd1 vccd1 _15229_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_172_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14183__B1 _16467_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18016_ _18959_/CLK _18016_/D vssd1 vssd1 vccd1 vccd1 _18016_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_141_HCLK clkbuf_4_3_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19842_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_160_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_146_HCLK_A clkbuf_4_1_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17366__S _17546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17121__A0 _15768_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15159_ _15159_/A vssd1 vssd1 vccd1 vccd1 _15160_/A sky130_fd_sc_hd__inv_2
XANTENNA__10744__B1 _10446_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19734__CLK _20051_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16475__A2 _16505_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19967_ _19970_/CLK _19967_/D repeater274/X vssd1 vssd1 vccd1 vccd1 _19967_/Q sky130_fd_sc_hd__dfrtp_1
X_09720_ _19416_/Q vssd1 vssd1 vccd1 vccd1 _09720_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11708__A _11730_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18918_ _19293_/CLK _18918_/D repeater188/X vssd1 vssd1 vccd1 vccd1 _18918_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12497__B1 _12386_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_234_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19898_ _19900_/CLK _19898_/D repeater195/X vssd1 vssd1 vccd1 vccd1 _19898_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_228_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09651_ _19992_/Q vssd1 vssd1 vccd1 vccd1 _09748_/A sky130_fd_sc_hd__inv_2
XFILLER_228_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18849_ _18866_/CLK _18849_/D repeater232/X vssd1 vssd1 vccd1 vccd1 _18849_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__14238__B2 _17600_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_216_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09582_ _20027_/Q _09580_/Y _09582_/B1 _09581_/X vssd1 vssd1 vccd1 vccd1 _20027_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__17188__A0 _15768_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16656__D _16656_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_224_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12258__B _12487_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_192_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17360__A0 _17486_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09016_ hold284/X vssd1 vssd1 vccd1 vccd1 _09016_/X sky130_fd_sc_hd__buf_4
XFILLER_191_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17276__S _17566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17112__A0 _17473_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold140 HADDR[23] vssd1 vssd1 vccd1 vccd1 input16/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 input35/X vssd1 vssd1 vccd1 vccd1 hold368/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 input3/X vssd1 vssd1 vccd1 vccd1 hold162/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 hold173/A vssd1 vssd1 vccd1 vccd1 hold173/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 HADDR[5] vssd1 vssd1 vccd1 vccd1 input28/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 hold195/A vssd1 vssd1 vccd1 vccd1 hold195/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_68_HCLK_A clkbuf_opt_3_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20107_ _20107_/CLK _20107_/D repeater233/X vssd1 vssd1 vccd1 vccd1 _20107_/Q sky130_fd_sc_hd__dfrtp_4
X_09918_ _19354_/Q vssd1 vssd1 vccd1 vccd1 _09918_/Y sky130_fd_sc_hd__inv_2
XFILLER_144_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19334__RESET_B repeater244/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20038_ _20049_/CLK _20038_/D repeater208/X vssd1 vssd1 vccd1 vccd1 _20038_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_218_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09849_ _09849_/A _10001_/A vssd1 vssd1 vccd1 vccd1 _09850_/B sky130_fd_sc_hd__or2_2
XFILLER_219_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12860_ _18926_/Q vssd1 vssd1 vccd1 vccd1 _13005_/A sky130_fd_sc_hd__inv_2
XPHY_4100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11811_ _19453_/Q _11807_/X _09061_/X _11808_/X vssd1 vssd1 vccd1 vccd1 _19453_/D
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_22_HCLK clkbuf_4_3_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20064_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_4144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17179__A0 _17486_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12791_ _18807_/Q vssd1 vssd1 vccd1 vccd1 _13531_/A sky130_fd_sc_hd__inv_2
XPHY_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14530_ _14532_/A vssd1 vssd1 vccd1 vccd1 _14530_/X sky130_fd_sc_hd__clkbuf_2
XPHY_4188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11742_ _11742_/A vssd1 vssd1 vccd1 vccd1 _15749_/B sky130_fd_sc_hd__clkbuf_2
XPHY_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14461_ _18362_/Q _14452_/A _14405_/X _14453_/A vssd1 vssd1 vccd1 vccd1 _18362_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11673_ _11671_/X _11672_/Y _18626_/Q _19542_/Q _11666_/X vssd1 vssd1 vccd1 vccd1
+ _19542_/D sky130_fd_sc_hd__a32o_1
XFILLER_186_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16200_ _18748_/Q _16114_/Y _16197_/X _16198_/X _16199_/Y vssd1 vssd1 vccd1 vccd1
+ _16200_/X sky130_fd_sc_hd__o221a_1
XPHY_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13412_ _20106_/Q _13430_/A _13409_/Y _18852_/Q _13411_/X vssd1 vssd1 vccd1 vccd1
+ _13417_/C sky130_fd_sc_hd__o221a_1
XFILLER_186_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10624_ _10573_/B _10618_/X _10584_/C _10608_/A vssd1 vssd1 vccd1 vccd1 _19807_/D
+ sky130_fd_sc_hd__o22ai_1
X_17180_ _17179_/X _12942_/Y _17541_/S vssd1 vssd1 vccd1 vccd1 _17180_/X sky130_fd_sc_hd__mux2_1
XPHY_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14392_ _14392_/A _15192_/A vssd1 vssd1 vccd1 vccd1 _14975_/C sky130_fd_sc_hd__or2_2
XPHY_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_164_HCLK clkbuf_4_0_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _18145_/CLK sky130_fd_sc_hd__clkbuf_16
X_16131_ _16123_/Y _16049_/X _16124_/Y _15836_/A _16130_/X vssd1 vssd1 vccd1 vccd1
+ _16131_/X sky130_fd_sc_hd__o221a_2
XFILLER_155_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13343_ _13429_/C _13450_/A vssd1 vssd1 vccd1 vccd1 _13344_/B sky130_fd_sc_hd__or2_1
X_10555_ _19812_/Q _19811_/Q vssd1 vssd1 vccd1 vccd1 _10939_/C sky130_fd_sc_hd__or2_2
XFILLER_182_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17351__A0 _17486_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18631__CLK _19780_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16062_ _19817_/Q vssd1 vssd1 vccd1 vccd1 _16062_/Y sky130_fd_sc_hd__inv_2
XFILLER_154_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13274_ _14270_/A _13274_/B vssd1 vssd1 vccd1 vccd1 _13293_/B sky130_fd_sc_hd__or2_1
X_10486_ _19532_/Q _19531_/Q _19530_/Q _19529_/Q vssd1 vssd1 vccd1 vccd1 _10514_/C
+ sky130_fd_sc_hd__or4_4
XANTENNA__17186__S _17544_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15013_ _18049_/Q _15010_/X _14992_/X _15012_/X vssd1 vssd1 vccd1 vccd1 _18049_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_182_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12225_ hold260/X vssd1 vssd1 vccd1 vccd1 _12225_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_108_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10726__B1 _10418_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19821_ _19822_/CLK _19821_/D repeater218/X vssd1 vssd1 vccd1 vccd1 _19821_/Q sky130_fd_sc_hd__dfrtp_1
X_12156_ _19279_/Q _12150_/X _12104_/X _12151_/X vssd1 vssd1 vccd1 vccd1 _19279_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_78_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11107_ _11105_/Y _17754_/S _19636_/Q _11091_/X vssd1 vssd1 vccd1 vccd1 _11119_/B
+ sky130_fd_sc_hd__o22a_1
X_19752_ _19900_/CLK _19752_/D repeater196/X vssd1 vssd1 vccd1 vccd1 _19752_/Q sky130_fd_sc_hd__dfrtp_1
X_16964_ _16963_/X _20026_/Q _17482_/S vssd1 vssd1 vccd1 vccd1 _16964_/X sky130_fd_sc_hd__mux2_2
X_12087_ _19319_/Q _12082_/X _12086_/X _12084_/X vssd1 vssd1 vccd1 vccd1 _19319_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_238_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18703_ _19119_/CLK _18703_/D hold351/X vssd1 vssd1 vccd1 vccd1 _18703_/Q sky130_fd_sc_hd__dfrtp_1
X_11038_ _17752_/X vssd1 vssd1 vccd1 vccd1 _11039_/A sky130_fd_sc_hd__inv_2
XFILLER_110_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15915_ _15915_/A vssd1 vssd1 vccd1 vccd1 _15915_/X sky130_fd_sc_hd__buf_2
X_19683_ _19795_/CLK _19683_/D repeater219/X vssd1 vssd1 vccd1 vccd1 _19683_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__11151__B1 _19648_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16895_ _17473_/A0 _16710_/Y _17473_/S vssd1 vssd1 vccd1 vccd1 _16895_/X sky130_fd_sc_hd__mux2_1
XANTENNA__19004__RESET_B hold346/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18634_ _19780_/CLK _18634_/D repeater225/X vssd1 vssd1 vccd1 vccd1 _18634_/Q sky130_fd_sc_hd__dfrtp_1
X_15846_ _15846_/A vssd1 vssd1 vccd1 vccd1 _15846_/X sky130_fd_sc_hd__buf_4
XFILLER_218_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18565_ _19841_/CLK _18565_/D repeater194/X vssd1 vssd1 vccd1 vccd1 _18565_/Q sky130_fd_sc_hd__dfrtp_1
X_12989_ _18938_/Q _12988_/Y _12980_/A _12881_/B vssd1 vssd1 vccd1 vccd1 _18938_/D
+ sky130_fd_sc_hd__o211a_1
X_15777_ _19261_/Q _18951_/Q vssd1 vssd1 vccd1 vccd1 _15777_/X sky130_fd_sc_hd__and2_1
XFILLER_18_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_1_0_HCLK clkbuf_4_1_0_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_1_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_221_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17516_ _17515_/X _15877_/Y _17539_/S vssd1 vssd1 vccd1 vccd1 _17516_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16917__A0 _15963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14728_ _18212_/Q _14718_/A _14727_/X _14719_/A vssd1 vssd1 vccd1 vccd1 _18212_/D
+ sky130_fd_sc_hd__a22o_1
X_18496_ _19794_/CLK _18496_/D repeater203/X vssd1 vssd1 vccd1 vccd1 _18496_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_232_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17447_ _17446_/X _09411_/Y _17529_/S vssd1 vssd1 vccd1 vccd1 _17447_/X sky130_fd_sc_hd__mux2_1
X_14659_ _18249_/Q _14656_/X _14600_/X _14658_/X vssd1 vssd1 vccd1 vccd1 _18249_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_21_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12403__B1 _12401_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17378_ _16272_/X _18231_/Q _17564_/S vssd1 vssd1 vccd1 vccd1 _17378_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19117_ _19119_/CLK _19117_/D hold353/X vssd1 vssd1 vccd1 vccd1 _19117_/Q sky130_fd_sc_hd__dfrtp_4
X_16329_ _18024_/Q vssd1 vssd1 vccd1 vccd1 _16329_/Y sky130_fd_sc_hd__inv_2
X_19048_ _19566_/CLK _19048_/D repeater255/X vssd1 vssd1 vccd1 vccd1 _19048_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_106_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19845__RESET_B repeater270/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17096__S _17543_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_247_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09703_ _09693_/X _09703_/B _09703_/C _09703_/D vssd1 vssd1 vccd1 vccd1 _09728_/B
+ sky130_fd_sc_hd__and4b_1
Xclkbuf_leaf_45_HCLK clkbuf_opt_2_HCLK/A vssd1 vssd1 vccd1 vccd1 _19540_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_67_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09634_ _19973_/Q vssd1 vssd1 vccd1 vccd1 _09807_/C sky130_fd_sc_hd__inv_2
XFILLER_228_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18798__RESET_B repeater258/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09565_ _09565_/A _09565_/B _09565_/C _09565_/D vssd1 vssd1 vccd1 vccd1 _09607_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_243_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18727__RESET_B repeater253/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09496_ _20035_/Q vssd1 vssd1 vccd1 vccd1 _09496_/Y sky130_fd_sc_hd__inv_2
XPHY_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12642__B1 _12032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17333__A0 _15768_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16903__S _17386_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10340_ _10340_/A vssd1 vssd1 vccd1 vccd1 _10341_/B sky130_fd_sc_hd__inv_2
XFILLER_164_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10271_ _19641_/Q vssd1 vssd1 vccd1 vccd1 _14316_/B sky130_fd_sc_hd__inv_2
XFILLER_117_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12010_ _12017_/A vssd1 vssd1 vccd1 vccd1 _12010_/X sky130_fd_sc_hd__buf_1
XFILLER_132_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17734__S _18508_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18034__CLK _19851_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10252__A _11936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13961_ _18709_/Q _13960_/Y _13947_/B _13901_/X vssd1 vssd1 vccd1 vccd1 _18709_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_47_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15700_ _18618_/Q vssd1 vssd1 vccd1 vccd1 _15700_/Y sky130_fd_sc_hd__inv_2
X_12912_ _19281_/Q _18938_/Q _12911_/Y _12965_/A vssd1 vssd1 vccd1 vccd1 _12916_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_19_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16680_ _19464_/Q vssd1 vssd1 vccd1 vccd1 _16680_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20073__RESET_B repeater196/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13892_ _19221_/Q _13830_/A _13891_/Y _18709_/Q vssd1 vssd1 vccd1 vccd1 _13892_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_73_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18184__CLK _18198_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15631_ _15629_/Y _15630_/X _15614_/X vssd1 vssd1 vccd1 vccd1 _15631_/X sky130_fd_sc_hd__o21a_1
X_12843_ _18941_/Q vssd1 vssd1 vccd1 vccd1 _12967_/B sky130_fd_sc_hd__inv_2
XFILLER_203_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18350_ _18959_/CLK _18350_/D vssd1 vssd1 vccd1 vccd1 _18350_/Q sky130_fd_sc_hd__dfxtp_1
X_15562_ _15562_/A vssd1 vssd1 vccd1 vccd1 _15562_/Y sky130_fd_sc_hd__inv_2
X_12774_ _19255_/Q vssd1 vssd1 vccd1 vccd1 _12774_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12633__B1 _12406_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17301_ _17300_/X _13538_/A _17386_/S vssd1 vssd1 vccd1 vccd1 _17301_/X sky130_fd_sc_hd__mux2_2
XPHY_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17798__S1 _19646_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14513_ _14727_/A vssd1 vssd1 vccd1 vccd1 _14513_/X sky130_fd_sc_hd__buf_2
XFILLER_214_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11725_ _19510_/Q _11723_/X _16942_/X _11724_/X vssd1 vssd1 vccd1 vccd1 hold217/A
+ sky130_fd_sc_hd__a22o_1
X_18281_ _19847_/CLK _18281_/D vssd1 vssd1 vccd1 vccd1 _18281_/Q sky130_fd_sc_hd__dfxtp_1
X_15493_ _18568_/Q vssd1 vssd1 vccd1 vccd1 _15493_/Y sky130_fd_sc_hd__inv_2
XPHY_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14394__A _14395_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14444_ _18375_/Q _14436_/X _14443_/X _14439_/X vssd1 vssd1 vccd1 vccd1 _18375_/D
+ sky130_fd_sc_hd__a22o_1
X_17232_ _17231_/X _11308_/Y _17459_/S vssd1 vssd1 vccd1 vccd1 _17232_/X sky130_fd_sc_hd__mux2_1
XPHY_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11656_ _11656_/A _15271_/A _15389_/C _11655_/X vssd1 vssd1 vccd1 vccd1 _11656_/X
+ sky130_fd_sc_hd__or4b_4
XPHY_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09450__A2_N _19383_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11739__A2 _11737_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10607_ _15224_/A _10617_/A vssd1 vssd1 vccd1 vccd1 _10608_/A sky130_fd_sc_hd__or2_2
X_17163_ _17162_/X _20018_/Q _17386_/S vssd1 vssd1 vccd1 vccd1 _17163_/X sky130_fd_sc_hd__mux2_2
XPHY_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17324__A0 _15963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14375_ _18412_/Q _14368_/A _14329_/X _14369_/A vssd1 vssd1 vccd1 vccd1 _18412_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16813__S _17546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11587_ _11592_/A vssd1 vssd1 vccd1 vccd1 _11588_/A sky130_fd_sc_hd__clkbuf_2
XPHY_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16114_ _17964_/Q vssd1 vssd1 vccd1 vccd1 _16114_/Y sky130_fd_sc_hd__inv_2
X_13326_ _18837_/Q vssd1 vssd1 vccd1 vccd1 _13327_/A sky130_fd_sc_hd__inv_2
X_10538_ _19814_/Q _10537_/B _15443_/A _10537_/Y vssd1 vssd1 vccd1 vccd1 _19814_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_171_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17094_ _17093_/X _14061_/Y _17490_/S vssd1 vssd1 vccd1 vccd1 _17094_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16045_ _20061_/Q _16204_/A vssd1 vssd1 vccd1 vccd1 _16045_/X sky130_fd_sc_hd__and2_1
X_13257_ _18750_/Q vssd1 vssd1 vccd1 vccd1 _13259_/A sky130_fd_sc_hd__inv_2
X_10469_ _19823_/Q _18549_/Q _10468_/Y _10460_/C vssd1 vssd1 vccd1 vccd1 _10470_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_89_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12208_ _19247_/Q _12205_/X _12098_/X _12206_/X vssd1 vssd1 vccd1 vccd1 _19247_/D
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_68_HCLK clkbuf_opt_3_HCLK/A vssd1 vssd1 vccd1 vccd1 _19920_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_170_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13188_ _18904_/Q _13187_/Y _13188_/B1 _13176_/X vssd1 vssd1 vccd1 vccd1 _18904_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_111_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19804_ _19808_/CLK _19804_/D repeater222/X vssd1 vssd1 vccd1 vccd1 _19804_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__11258__A _19023_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17644__S _17655_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12139_ _19292_/Q _12134_/X _12074_/X _12137_/X vssd1 vssd1 vccd1 vccd1 _19292_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_123_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17996_ _18412_/CLK _17996_/D vssd1 vssd1 vccd1 vccd1 _17996_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_51_HCLK_A clkbuf_opt_1_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14310__B1 _13676_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19735_ _20051_/CLK _19735_/D repeater208/X vssd1 vssd1 vccd1 vccd1 _19735_/Q sky130_fd_sc_hd__dfrtp_1
X_16947_ _19491_/Q hold142/X _16950_/S vssd1 vssd1 vccd1 vccd1 _16947_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19666_ _19855_/CLK _19666_/D repeater264/X vssd1 vssd1 vccd1 vccd1 _19666_/Q sky130_fd_sc_hd__dfrtp_4
X_16878_ _16877_/X _09482_/A _17482_/S vssd1 vssd1 vccd1 vccd1 _16878_/X sky130_fd_sc_hd__mux2_1
X_18617_ _19577_/CLK _18617_/D repeater269/X vssd1 vssd1 vccd1 vccd1 _18617_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_64_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15829_ _15858_/C _15829_/B _16492_/A vssd1 vssd1 vccd1 vccd1 _15830_/A sky130_fd_sc_hd__or3_4
X_19597_ _19597_/CLK _19597_/D hold273/X vssd1 vssd1 vccd1 vccd1 _19597_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_213_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18820__RESET_B repeater231/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09350_ _20027_/Q vssd1 vssd1 vccd1 vccd1 _09487_/A sky130_fd_sc_hd__inv_2
X_18548_ _19780_/CLK _18548_/D repeater229/X vssd1 vssd1 vccd1 vccd1 _18548_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__11427__B2 _19130_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12624__B1 _12389_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17789__S1 _19648_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09281_ _19498_/Q vssd1 vssd1 vccd1 vccd1 _10429_/A sky130_fd_sc_hd__inv_2
X_18479_ _19780_/CLK _18479_/D repeater227/X vssd1 vssd1 vccd1 vccd1 _18479_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_221_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14377__B1 _14314_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18057__CLK _18169_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15863__A _19125_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08996_ _12130_/A _12130_/B _13279_/C vssd1 vssd1 vccd1 vccd1 _15890_/A sky130_fd_sc_hd__or3_4
XFILLER_125_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16678__B _16678_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_217_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18908__RESET_B repeater188/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09617_ _09467_/A _09467_/B _09615_/Y _09607_/X vssd1 vssd1 vccd1 vccd1 _20006_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_18_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_243_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09548_ _19314_/Q vssd1 vssd1 vccd1 vccd1 _16620_/A sky130_fd_sc_hd__inv_2
XFILLER_243_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12091__A1 _19317_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09479_ _09479_/A _09595_/A vssd1 vssd1 vccd1 vccd1 _09480_/B sky130_fd_sc_hd__or2_2
XPHY_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11510_ _11478_/A _11478_/B _11506_/X _11508_/Y vssd1 vssd1 vccd1 vccd1 _19598_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12490_ _12528_/A vssd1 vssd1 vccd1 vccd1 _12529_/A sky130_fd_sc_hd__inv_2
XFILLER_211_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17729__S _18508_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11441_ _19564_/Q vssd1 vssd1 vccd1 vccd1 _11577_/A sky130_fd_sc_hd__inv_2
XFILLER_7_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14160_ _19103_/Q vssd1 vssd1 vccd1 vccd1 _14160_/Y sky130_fd_sc_hd__inv_2
X_11372_ _19552_/Q vssd1 vssd1 vccd1 vccd1 _11622_/A sky130_fd_sc_hd__inv_2
XFILLER_152_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13111_ _19171_/Q vssd1 vssd1 vccd1 vccd1 _13111_/Y sky130_fd_sc_hd__inv_2
X_10323_ _10323_/A _10371_/A vssd1 vssd1 vccd1 vccd1 _10366_/A sky130_fd_sc_hd__or2_1
XFILLER_3_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14091_ _19092_/Q _14034_/Y _19085_/Q _14026_/A vssd1 vssd1 vccd1 vccd1 _14091_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_124_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14540__B1 hold330/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13042_ _18904_/Q vssd1 vssd1 vccd1 vccd1 _13076_/A sky130_fd_sc_hd__inv_2
X_10254_ _19496_/Q _19495_/Q vssd1 vssd1 vccd1 vccd1 _10410_/A sky130_fd_sc_hd__or2_4
XFILLER_106_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12181__B _12309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17464__S _17565_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17850_ _16328_/Y _16329_/Y _16330_/Y _16331_/Y _17913_/S0 _19632_/Q vssd1 vssd1
+ vccd1 vccd1 _17850_/X sky130_fd_sc_hd__mux4_2
X_10185_ _17631_/X _10181_/A _19876_/Q _15715_/B vssd1 vssd1 vccd1 vccd1 _19876_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_239_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16588__B _16615_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16801_ _15963_/X _09522_/Y _17534_/S vssd1 vssd1 vccd1 vccd1 _16801_/X sky130_fd_sc_hd__mux2_1
X_17781_ _18389_/Q _18381_/Q _18373_/Q _18365_/Q _17923_/S0 _19646_/Q vssd1 vssd1
+ vccd1 vccd1 _17781_/X sky130_fd_sc_hd__mux4_2
X_14993_ _14993_/A vssd1 vssd1 vccd1 vccd1 _14994_/A sky130_fd_sc_hd__inv_2
X_19520_ _19814_/CLK _19520_/D repeater223/X vssd1 vssd1 vccd1 vccd1 _19520_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_115_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16732_ _16891_/X _16683_/X _16894_/X _16684_/X _16731_/X vssd1 vssd1 vccd1 vccd1
+ _16735_/B sky130_fd_sc_hd__o221a_2
X_13944_ _13964_/A _13964_/B _13944_/C vssd1 vssd1 vccd1 vccd1 _13962_/A sky130_fd_sc_hd__or3_1
XFILLER_235_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19945__CLK _19976_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19451_ _19841_/CLK _19451_/D repeater271/X vssd1 vssd1 vccd1 vccd1 _19451_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_235_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16663_ _16989_/X _16577_/X _17045_/X _16578_/X _16662_/X vssd1 vssd1 vccd1 vccd1
+ _16664_/C sky130_fd_sc_hd__o221a_1
X_13875_ _19200_/Q vssd1 vssd1 vccd1 vccd1 _13875_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16808__S _17535_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_repeater192_A repeater193/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18402_ _18954_/CLK _18402_/D vssd1 vssd1 vccd1 vccd1 _18402_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12826_ _12821_/Y _18810_/Q _12822_/Y _18820_/Q _12825_/X vssd1 vssd1 vccd1 vccd1
+ _12833_/C sky130_fd_sc_hd__o221a_1
X_15614_ _15643_/A vssd1 vssd1 vccd1 vccd1 _15614_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_62_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19382_ _19920_/CLK _19382_/D repeater230/X vssd1 vssd1 vccd1 vccd1 _19382_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12606__B1 _12538_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16594_ _16594_/A vssd1 vssd1 vccd1 vccd1 _16594_/X sky130_fd_sc_hd__buf_1
XFILLER_222_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18333_ _18333_/CLK _18333_/D vssd1 vssd1 vccd1 vccd1 _18333_/Q sky130_fd_sc_hd__dfxtp_1
X_12757_ _12752_/Y _18811_/Q _19232_/Q _13533_/A _12756_/X vssd1 vssd1 vccd1 vccd1
+ _12758_/D sky130_fd_sc_hd__o221a_1
X_15545_ _18580_/Q _15547_/B vssd1 vssd1 vccd1 vccd1 _15550_/B sky130_fd_sc_hd__or2_1
XPHY_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12637__A _12651_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11708_ _11730_/A vssd1 vssd1 vccd1 vccd1 _11708_/X sky130_fd_sc_hd__clkbuf_2
X_15476_ _15474_/Y _15475_/Y _15459_/X vssd1 vssd1 vccd1 vccd1 _15476_/X sky130_fd_sc_hd__o21a_1
X_18264_ _20079_/CLK _18264_/D vssd1 vssd1 vccd1 vccd1 _18264_/Q sky130_fd_sc_hd__dfxtp_1
X_12688_ _18974_/Q _12684_/X _12028_/A _12685_/X vssd1 vssd1 vccd1 vccd1 _18974_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14427_ _18385_/Q _14424_/X _14351_/X _14426_/X vssd1 vssd1 vccd1 vccd1 _18385_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17639__S _17655_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17215_ _16484_/X _08934_/Y _17566_/S vssd1 vssd1 vccd1 vccd1 _17215_/X sky130_fd_sc_hd__mux2_1
X_11639_ _11639_/A _11639_/B _11639_/C vssd1 vssd1 vccd1 vccd1 _11642_/A sky130_fd_sc_hd__or3_4
XFILLER_30_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18195_ _18333_/CLK _18195_/D vssd1 vssd1 vccd1 vccd1 _18195_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__19437__RESET_B repeater269/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17146_ _17145_/X _09479_/A _17536_/S vssd1 vssd1 vccd1 vccd1 _17146_/X sky130_fd_sc_hd__mux2_2
X_14358_ hold245/X vssd1 vssd1 vccd1 vccd1 _14751_/A sky130_fd_sc_hd__clkbuf_2
X_13309_ _18856_/Q vssd1 vssd1 vccd1 vccd1 _13429_/C sky130_fd_sc_hd__inv_6
X_17077_ _17486_/A0 _13115_/Y _17543_/S vssd1 vssd1 vccd1 vccd1 _17077_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12372__A _12372_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14289_ _14289_/A vssd1 vssd1 vccd1 vccd1 _14290_/A sky130_fd_sc_hd__inv_2
XFILLER_115_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16028_ _17947_/Q vssd1 vssd1 vccd1 vccd1 _16028_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17374__S _17564_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09681__A _19422_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17979_ _20123_/CLK _17979_/D vssd1 vssd1 vccd1 vccd1 _17979_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19718_ _19720_/CLK _19718_/D repeater190/X vssd1 vssd1 vccd1 vccd1 _19718_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__11716__A _11730_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_242_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19649_ _19867_/CLK _19649_/D repeater261/X vssd1 vssd1 vccd1 vccd1 _19649_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_38_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09402_ _19925_/Q vssd1 vssd1 vccd1 vccd1 _10041_/A sky130_fd_sc_hd__inv_2
XFILLER_19_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09333_ _09333_/A _09333_/B _18661_/D _09332_/X vssd1 vssd1 vccd1 vccd1 _13766_/D
+ sky130_fd_sc_hd__or4b_4
XFILLER_179_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12073__A1 _19325_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09264_ _10186_/A _09340_/B _15961_/A vssd1 vssd1 vccd1 vccd1 _09265_/S sky130_fd_sc_hd__or3_1
XFILLER_193_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15858__A _15858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09195_ _09192_/A _08983_/X _09192_/Y vssd1 vssd1 vccd1 vccd1 _20071_/D sky130_fd_sc_hd__a21oi_1
XANTENNA__19178__RESET_B repeater212/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16511__B2 _16235_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14522__B1 _14441_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17284__S _17318_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold285_A HWDATA[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08979_ _17605_/S _10133_/C vssd1 vssd1 vccd1 vccd1 _08982_/B sky130_fd_sc_hd__or2_1
XFILLER_217_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11990_ _11841_/X _19365_/Q _11990_/S vssd1 vssd1 vccd1 vccd1 _19365_/D sky130_fd_sc_hd__mux2_1
X_10941_ _10583_/A _10940_/X _10584_/C vssd1 vssd1 vccd1 vccd1 _10942_/B sky130_fd_sc_hd__o21ai_1
XFILLER_217_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13660_ _18786_/Q _13656_/X _12028_/A _13658_/X vssd1 vssd1 vccd1 vccd1 _18786_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_16_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_244_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10872_ _15349_/A vssd1 vssd1 vccd1 vccd1 _15364_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__17870__S0 _17913_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12611_ _15769_/A _12659_/B vssd1 vssd1 vccd1 vccd1 _12650_/A sky130_fd_sc_hd__or2_4
XANTENNA__19948__RESET_B hold371/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13591_ _13591_/A vssd1 vssd1 vccd1 vccd1 _13591_/X sky130_fd_sc_hd__clkbuf_2
XPHY_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12457__A _12457_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10075__B1 _10026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15330_ _15330_/A _15832_/A vssd1 vssd1 vccd1 vccd1 _18476_/D sky130_fd_sc_hd__nor2_2
XPHY_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12542_ _19062_/Q _12505_/A _12541_/X _12506_/A vssd1 vssd1 vccd1 vccd1 _19062_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_212_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15261_ _15437_/B _18632_/Q _15263_/A _15250_/Y _15260_/X vssd1 vssd1 vccd1 vccd1
+ _15261_/X sky130_fd_sc_hd__a32o_1
XANTENNA__17459__S _17459_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15768__A _15863_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12473_ _19104_/Q _12471_/X _12353_/X _12472_/X vssd1 vssd1 vccd1 vccd1 _19104_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_184_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19530__RESET_B repeater221/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17000_ _15768_/Y _11283_/Y _17546_/S vssd1 vssd1 vccd1 vccd1 _17000_/X sky130_fd_sc_hd__mux2_1
X_14212_ _19106_/Q vssd1 vssd1 vccd1 vccd1 _14212_/Y sky130_fd_sc_hd__inv_2
X_11424_ _19576_/Q vssd1 vssd1 vccd1 vccd1 _11561_/A sky130_fd_sc_hd__inv_2
XFILLER_6_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15192_ _15192_/A _15192_/B vssd1 vssd1 vccd1 vccd1 _15192_/Y sky130_fd_sc_hd__nor2_1
Xclkbuf_3_5_0_HCLK clkbuf_3_5_0_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_14143_ _18677_/Q _14142_/Y _14143_/B1 _14112_/X vssd1 vssd1 vccd1 vccd1 _18677_/D
+ sky130_fd_sc_hd__o211a_1
X_11355_ _18980_/Q vssd1 vssd1 vccd1 vccd1 _11355_/Y sky130_fd_sc_hd__inv_2
XFILLER_180_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10306_ _18604_/Q _18607_/Q _18611_/Q vssd1 vssd1 vccd1 vccd1 _10308_/C sky130_fd_sc_hd__or3_2
XFILLER_152_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14074_ _19072_/Q vssd1 vssd1 vccd1 vccd1 _14074_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18951_ _20035_/CLK _18951_/D repeater216/X vssd1 vssd1 vccd1 vccd1 _18951_/Q sky130_fd_sc_hd__dfrtp_1
X_11286_ _19017_/Q vssd1 vssd1 vccd1 vccd1 _11286_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17194__S _17546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17902_ _15927_/Y _15928_/Y _15929_/Y _15930_/Y _17913_/S0 _19632_/Q vssd1 vssd1
+ vccd1 vccd1 _17902_/X sky130_fd_sc_hd__mux4_1
X_13025_ _12859_/B _13024_/A _18921_/Q _13027_/A _12962_/X vssd1 vssd1 vccd1 vccd1
+ _18921_/D sky130_fd_sc_hd__o221a_1
X_10237_ _19661_/Q vssd1 vssd1 vccd1 vccd1 _10996_/A sky130_fd_sc_hd__inv_2
X_18882_ _19814_/CLK _18882_/D repeater220/X vssd1 vssd1 vccd1 vccd1 _18882_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_79_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater205_A repeater207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17833_ _17934_/Q _18456_/Q _18464_/Q _18064_/Q _17918_/S0 _18750_/Q vssd1 vssd1
+ vccd1 vccd1 _17833_/X sky130_fd_sc_hd__mux4_2
XFILLER_86_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10168_ _10175_/A vssd1 vssd1 vccd1 vccd1 _10168_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_66_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17764_ _15192_/Y _13254_/Y _17764_/S vssd1 vssd1 vccd1 vccd1 _17764_/X sky130_fd_sc_hd__mux2_2
X_10099_ _10099_/A vssd1 vssd1 vccd1 vccd1 _10103_/A sky130_fd_sc_hd__inv_2
X_14976_ _14978_/A vssd1 vssd1 vccd1 vccd1 _14976_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_212_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19503_ _19510_/CLK hold232/X repeater256/X vssd1 vssd1 vccd1 vccd1 _19503_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_63_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16715_ _16682_/X _16715_/B _16715_/C vssd1 vssd1 vccd1 vccd1 _16715_/Y sky130_fd_sc_hd__nand3b_4
XFILLER_75_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13927_ _13927_/A vssd1 vssd1 vccd1 vccd1 _13927_/X sky130_fd_sc_hd__clkbuf_4
X_17695_ _15451_/Y _19440_/Q _17696_/S vssd1 vssd1 vccd1 vccd1 _18557_/D sky130_fd_sc_hd__mux2_1
XFILLER_207_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19434_ _19513_/CLK _19434_/D repeater259/X vssd1 vssd1 vccd1 vccd1 _19434_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_222_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16646_ _16646_/A _16647_/B vssd1 vssd1 vccd1 vccd1 _16646_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__17861__S0 _17913_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13858_ _19195_/Q vssd1 vssd1 vccd1 vccd1 _13858_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14044__A2 _18701_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12809_ _18808_/Q vssd1 vssd1 vccd1 vccd1 _13532_/A sky130_fd_sc_hd__inv_2
X_19365_ _19905_/CLK _19365_/D repeater210/X vssd1 vssd1 vccd1 vccd1 _19365_/Q sky130_fd_sc_hd__dfrtp_1
X_16577_ _16687_/A vssd1 vssd1 vccd1 vccd1 _16577_/X sky130_fd_sc_hd__clkbuf_2
X_13789_ _18723_/Q vssd1 vssd1 vccd1 vccd1 _13910_/C sky130_fd_sc_hd__inv_2
XFILLER_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19618__RESET_B repeater230/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11271__A _19009_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18316_ _18435_/CLK _18316_/D vssd1 vssd1 vccd1 vccd1 _18316_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15528_ _18576_/Q vssd1 vssd1 vccd1 vccd1 _15530_/A sky130_fd_sc_hd__clkbuf_2
X_19296_ _20013_/CLK _19296_/D repeater241/X vssd1 vssd1 vccd1 vccd1 _19296_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_187_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17369__S _19498_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18247_ _18465_/CLK _18247_/D vssd1 vssd1 vccd1 vccd1 _18247_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15459_ _15512_/A vssd1 vssd1 vccd1 vccd1 _15459_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_129_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16741__B2 _16002_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14752__B1 _14751_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18178_ _18460_/CLK _18178_/D vssd1 vssd1 vccd1 vccd1 _18178_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17916__S1 _18750_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17129_ _17128_/X _09862_/A _17414_/S vssd1 vssd1 vccd1 vccd1 _17129_/X sky130_fd_sc_hd__mux2_1
X_09951_ _19970_/Q _09878_/Y _09879_/Y _09878_/A _09950_/X vssd1 vssd1 vccd1 vccd1
+ _19970_/D sky130_fd_sc_hd__o221a_1
XANTENNA__20105__RESET_B repeater230/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09882_ _09879_/Y _19362_/Q _19948_/Q _09880_/Y _09881_/X vssd1 vssd1 vccd1 vccd1
+ _09895_/A sky130_fd_sc_hd__o221a_1
X_20071_ _20124_/CLK _20071_/D repeater207/X vssd1 vssd1 vccd1 vccd1 _20071_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_98_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18245__CLK _19847_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17852__S0 _17913_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09316_ _18654_/Q vssd1 vssd1 vccd1 vccd1 _15721_/A sky130_fd_sc_hd__buf_1
XFILLER_139_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16691__B _16691_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17279__S _17318_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09247_ _20064_/Q _20065_/Q _09250_/S vssd1 vssd1 vccd1 vccd1 _20065_/D sky130_fd_sc_hd__mux2_1
XFILLER_167_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold200_A HADDR[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09178_ _14709_/A _09163_/X _09177_/X _09165_/X vssd1 vssd1 vccd1 vccd1 _20077_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_147_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17907__S1 _18759_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16911__S _17523_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16496__B1 _17221_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11140_ _19226_/Q vssd1 vssd1 vccd1 vccd1 _15232_/A sky130_fd_sc_hd__buf_1
XFILLER_123_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11071_ _14378_/B _11064_/B _14489_/B _19631_/Q _11070_/Y vssd1 vssd1 vccd1 vccd1
+ _11076_/B sky130_fd_sc_hd__a221o_1
XFILLER_248_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput89 _16614_/Y vssd1 vssd1 vccd1 vccd1 HRDATA[19] sky130_fd_sc_hd__clkbuf_2
XANTENNA__16248__B1 _17399_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10022_ _10047_/C _10048_/A _10022_/C _10051_/A vssd1 vssd1 vccd1 vccd1 _10023_/C
+ sky130_fd_sc_hd__or4_4
XFILLER_88_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17742__S _18508_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14830_ _18154_/Q _14821_/A _14782_/X _14822_/A vssd1 vssd1 vccd1 vccd1 _18154_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10260__A _19873_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11973_ _19375_/Q _11969_/X _11909_/X _11970_/X vssd1 vssd1 vccd1 vccd1 _19375_/D
+ sky130_fd_sc_hd__a22o_1
X_14761_ _14761_/A vssd1 vssd1 vccd1 vccd1 _14761_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_91_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16500_ _19272_/Q vssd1 vssd1 vccd1 vccd1 _16500_/Y sky130_fd_sc_hd__inv_2
X_10924_ _10924_/A vssd1 vssd1 vccd1 vccd1 _10924_/X sky130_fd_sc_hd__clkbuf_2
X_13712_ _13706_/A _13704_/B _13704_/A vssd1 vssd1 vccd1 vccd1 _13712_/X sky130_fd_sc_hd__o21a_1
XFILLER_232_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10835__A2 _10831_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17480_ _15963_/X _09551_/Y _17534_/S vssd1 vssd1 vccd1 vccd1 _17480_/X sky130_fd_sc_hd__mux2_1
X_14692_ _18227_/Q _14683_/A _14691_/X _14684_/A vssd1 vssd1 vccd1 vccd1 _18227_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17843__S0 _17913_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19782__RESET_B repeater204/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16431_ _18105_/Q vssd1 vssd1 vccd1 vccd1 _16431_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13234__B1 _18545_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10855_ _10856_/A vssd1 vssd1 vccd1 vccd1 _10855_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_31_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13643_ _13646_/A vssd1 vssd1 vccd1 vccd1 _13644_/A sky130_fd_sc_hd__inv_2
XANTENNA__18738__CLK _20051_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12187__A _12187_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19150_ _19597_/CLK _19150_/D repeater281/X vssd1 vssd1 vccd1 vccd1 _19150_/Q sky130_fd_sc_hd__dfrtp_4
X_13574_ _13591_/A vssd1 vssd1 vccd1 vccd1 _13574_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_31_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14982__B1 hold236/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16362_ _18112_/Q vssd1 vssd1 vccd1 vccd1 _16362_/Y sky130_fd_sc_hd__inv_2
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10786_ _19740_/Q _10786_/B vssd1 vssd1 vccd1 vccd1 _10786_/Y sky130_fd_sc_hd__nand2_1
XFILLER_169_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11796__B1 _09033_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18101_ _18137_/CLK _18101_/D vssd1 vssd1 vccd1 vccd1 _18101_/Q sky130_fd_sc_hd__dfxtp_1
X_15313_ _11648_/A _15437_/B _15312_/Y _15245_/X vssd1 vssd1 vccd1 vccd1 _15313_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_9_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17189__S _17544_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12525_ hold260/X vssd1 vssd1 vccd1 vccd1 hold259/A sky130_fd_sc_hd__clkbuf_4
XFILLER_9_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19081_ _19115_/CLK _19081_/D hold353/X vssd1 vssd1 vccd1 vccd1 _19081_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16293_ _18802_/Q _16043_/Y _18803_/Q _16114_/Y vssd1 vssd1 vccd1 vccd1 _16293_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA_repeater155_A _17517_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18032_ _18142_/CLK _18032_/D vssd1 vssd1 vccd1 vccd1 _18032_/Q sky130_fd_sc_hd__dfxtp_1
X_15244_ _19824_/Q _19823_/Q _19825_/Q vssd1 vssd1 vccd1 vccd1 _15263_/A sky130_fd_sc_hd__or3_4
XFILLER_173_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12456_ _19115_/Q _12450_/X _12398_/X _12451_/X vssd1 vssd1 vccd1 vccd1 _19115_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_172_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11407_ _19561_/Q vssd1 vssd1 vccd1 vccd1 _11574_/A sky130_fd_sc_hd__inv_2
X_15175_ _17942_/Q _15170_/X hold244/X _15172_/X vssd1 vssd1 vccd1 vccd1 _17942_/D
+ sky130_fd_sc_hd__a22o_1
X_12387_ _19153_/Q _12374_/X _12386_/X _12378_/X vssd1 vssd1 vccd1 vccd1 _19153_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16821__S _17542_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output84_A _16559_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14126_ _14126_/A vssd1 vssd1 vccd1 vccd1 _14126_/Y sky130_fd_sc_hd__clkinv_1
X_11338_ _18983_/Q vssd1 vssd1 vccd1 vccd1 _11338_/Y sky130_fd_sc_hd__inv_2
XFILLER_180_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19983_ _19992_/CLK _19983_/D repeater192/X vssd1 vssd1 vccd1 vccd1 _19983_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_125_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18934_ _19315_/CLK _18934_/D repeater213/X vssd1 vssd1 vccd1 vccd1 _18934_/Q sky130_fd_sc_hd__dfrtp_4
X_14057_ _19089_/Q vssd1 vssd1 vccd1 vccd1 _14057_/Y sky130_fd_sc_hd__inv_2
X_11269_ _19006_/Q vssd1 vssd1 vccd1 vccd1 _16542_/A sky130_fd_sc_hd__inv_2
XANTENNA__12650__A _12650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13008_ _13008_/A _13008_/B vssd1 vssd1 vccd1 vccd1 _13008_/Y sky130_fd_sc_hd__nor2_1
XFILLER_79_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18865_ _20107_/CLK _18865_/D repeater233/X vssd1 vssd1 vccd1 vccd1 _18865_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_121_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18666__SET_B repeater222/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17652__S _17655_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17816_ _18189_/Q _18181_/Q _18173_/Q _18157_/Q _17918_/S0 _18750_/Q vssd1 vssd1
+ vccd1 vccd1 _17816_/X sky130_fd_sc_hd__mux4_1
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18796_ _19435_/CLK _18796_/D repeater258/X vssd1 vssd1 vccd1 vccd1 _18796_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_67_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17747_ _15318_/Y _11059_/Y _17755_/S vssd1 vssd1 vccd1 vccd1 _17747_/X sky130_fd_sc_hd__mux2_2
X_14959_ _18077_/Q _14952_/X _14931_/X _14954_/X vssd1 vssd1 vccd1 vccd1 _18077_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_223_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17834__S0 _18751_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_106_HCLK_A clkbuf_4_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17678_ _15521_/X _19457_/Q _17696_/S vssd1 vssd1 vccd1 vccd1 _18574_/D sky130_fd_sc_hd__mux2_1
XFILLER_51_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19417_ _19905_/CLK _19417_/D repeater210/X vssd1 vssd1 vccd1 vccd1 _19417_/Q sky130_fd_sc_hd__dfrtp_4
X_16629_ _16629_/A _16629_/B _16629_/C _16629_/D vssd1 vssd1 vccd1 vccd1 _16629_/X
+ sky130_fd_sc_hd__or4_4
XFILLER_22_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_3_2_0_HCLK_A clkbuf_3_3_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19452__RESET_B repeater272/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19348_ _19352_/CLK _19348_/D repeater245/X vssd1 vssd1 vccd1 vccd1 _19348_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_188_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09101_ _10423_/A vssd1 vssd1 vccd1 vccd1 _09101_/X sky130_fd_sc_hd__buf_4
XANTENNA__17099__S _17534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19279_ _19283_/CLK _19279_/D repeater212/X vssd1 vssd1 vccd1 vccd1 _19279_/Q sky130_fd_sc_hd__dfrtp_4
X_09032_ _20117_/Q _09029_/X _09030_/X _09031_/X vssd1 vssd1 vccd1 vccd1 _20117_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_176_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold300 hold300/A vssd1 vssd1 vccd1 vccd1 hold300/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold311 HWDATA[18] vssd1 vssd1 vccd1 vccd1 input47/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold322 input38/X vssd1 vssd1 vccd1 vccd1 hold322/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold333 HWDATA[3] vssd1 vssd1 vccd1 vccd1 input63/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16478__B1 _16903_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold344 input74/X vssd1 vssd1 vccd1 vccd1 hold344/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold355 hold355/A vssd1 vssd1 vccd1 vccd1 hold355/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold366 hold366/A vssd1 vssd1 vccd1 vccd1 hold366/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20123_ _20123_/CLK _20123_/D repeater196/X vssd1 vssd1 vccd1 vccd1 _20123_/Q sky130_fd_sc_hd__dfrtp_2
X_09934_ _19332_/Q vssd1 vssd1 vccd1 vccd1 _09934_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20054_ _20055_/CLK _20054_/D repeater205/X vssd1 vssd1 vccd1 vccd1 _20054_/Q sky130_fd_sc_hd__dfrtp_1
X_09865_ _09865_/A _09865_/B vssd1 vssd1 vccd1 vccd1 _09972_/A sky130_fd_sc_hd__or2_1
XANTENNA__20020__CLK _20091_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11176__A _11191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17562__S _17567_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09796_ _09794_/A _09794_/B _09734_/A _09794_/Y vssd1 vssd1 vccd1 vccd1 _19982_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_133_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater150 _17487_/S vssd1 vssd1 vccd1 vccd1 _17541_/S sky130_fd_sc_hd__buf_8
XFILLER_246_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater161 _17547_/S vssd1 vssd1 vccd1 vccd1 _17493_/S sky130_fd_sc_hd__buf_8
Xrepeater172 _17488_/S vssd1 vssd1 vccd1 vccd1 _17542_/S sky130_fd_sc_hd__buf_8
XPHY_4304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater183 _18758_/Q vssd1 vssd1 vccd1 vccd1 _17908_/S0 sky130_fd_sc_hd__clkbuf_16
XPHY_4315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater194 repeater198/X vssd1 vssd1 vccd1 vccd1 repeater194/X sky130_fd_sc_hd__buf_6
XPHY_4326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17825__S0 _17918_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16906__S _17490_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_242_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10640_ _10640_/A vssd1 vssd1 vccd1 vccd1 _19797_/D sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_28_HCLK_A clkbuf_4_9_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10571_ _19807_/Q vssd1 vssd1 vccd1 vccd1 _10573_/B sky130_fd_sc_hd__inv_2
XFILLER_210_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16207__A _16721_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12310_ _12180_/X _19192_/Q _12310_/S vssd1 vssd1 vccd1 vccd1 _19192_/D sky130_fd_sc_hd__mux2_1
XFILLER_158_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13290_ _14270_/B _17918_/S0 _14286_/B _13259_/B _17758_/X vssd1 vssd1 vccd1 vccd1
+ _13299_/B sky130_fd_sc_hd__o221ai_1
XFILLER_213_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20027__RESET_B repeater239/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17737__S _18508_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12241_ _14405_/A vssd1 vssd1 vccd1 vccd1 _12241_/X sky130_fd_sc_hd__buf_4
XANTENNA__14192__B2 _18681_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10255__A _15823_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12172_ _12172_/A vssd1 vssd1 vccd1 vccd1 _12172_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_122_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11950__B1 _09030_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11123_ _11123_/A _11123_/B vssd1 vssd1 vccd1 vccd1 _11124_/A sky130_fd_sc_hd__or2_1
XFILLER_174_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15141__B1 _10715_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16980_ _17804_/X _19898_/Q _16986_/S vssd1 vssd1 vccd1 vccd1 _16980_/X sky130_fd_sc_hd__mux2_1
XFILLER_107_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11054_ _14517_/A _14317_/B _11049_/Y _14335_/A _11053_/X vssd1 vssd1 vccd1 vccd1
+ _19644_/D sky130_fd_sc_hd__a32o_1
XFILLER_77_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15931_ _18339_/Q vssd1 vssd1 vccd1 vccd1 _15931_/Y sky130_fd_sc_hd__inv_2
XFILLER_190_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17472__S _17568_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10005_ _19938_/Q _09990_/X _10004_/Y vssd1 vssd1 vccd1 vccd1 _19938_/D sky130_fd_sc_hd__o21a_1
XFILLER_67_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18650_ _20050_/CLK _18650_/D repeater206/X vssd1 vssd1 vccd1 vccd1 _18650_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_209_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15862_ _19024_/Q _15863_/B vssd1 vssd1 vccd1 vccd1 _15862_/Y sky130_fd_sc_hd__nor2_1
XFILLER_77_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19963__RESET_B hold370/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17601_ _10133_/X _16986_/S _17605_/S vssd1 vssd1 vccd1 vccd1 _17601_/X sky130_fd_sc_hd__mux2_1
X_14813_ _18165_/Q _14801_/X _14812_/X _14804_/X vssd1 vssd1 vccd1 vccd1 _18165_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18581_ _19561_/CLK _18581_/D repeater274/X vssd1 vssd1 vccd1 vccd1 _18581_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_236_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15793_ _18346_/Q vssd1 vssd1 vccd1 vccd1 _15793_/Y sky130_fd_sc_hd__inv_2
XANTENNA_output122_A _15750_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18560__CLK _19992_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10269__B1 _19648_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17532_ _17531_/X _12733_/Y _17548_/S vssd1 vssd1 vccd1 vccd1 _17532_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11814__A _11821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_217_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14744_ _14746_/A vssd1 vssd1 vccd1 vccd1 _14744_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__17816__S0 _17918_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11956_ _11956_/A vssd1 vssd1 vccd1 vccd1 _11956_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_33_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10907_ _15215_/B _10907_/B vssd1 vssd1 vccd1 vccd1 _10908_/A sky130_fd_sc_hd__or2_2
X_17463_ _16044_/Y _16043_/Y _17564_/S vssd1 vssd1 vccd1 vccd1 _17463_/X sky130_fd_sc_hd__mux2_1
X_11887_ _19426_/Q _11884_/X _09033_/X _11885_/X vssd1 vssd1 vccd1 vccd1 _19426_/D
+ sky130_fd_sc_hd__a22o_1
X_14675_ _18238_/Q _14669_/X _09177_/X _14671_/X vssd1 vssd1 vccd1 vccd1 _18238_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16816__S _17534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19202_ _19585_/CLK _19202_/D hold365/X vssd1 vssd1 vccd1 vccd1 _19202_/Q sky130_fd_sc_hd__dfrtp_1
X_16414_ _18249_/Q _16433_/B vssd1 vssd1 vccd1 vccd1 _16414_/X sky130_fd_sc_hd__or2_1
X_10838_ _15349_/A _10831_/B _15735_/A _10712_/Y _10840_/S vssd1 vssd1 vccd1 vccd1
+ _10839_/A sky130_fd_sc_hd__o32a_1
X_13626_ _18800_/Q _13616_/B _13617_/A _13620_/Y vssd1 vssd1 vccd1 vccd1 _13626_/X
+ sky130_fd_sc_hd__o211a_1
X_17394_ _16205_/Y _09229_/Y _19498_/Q vssd1 vssd1 vccd1 vccd1 _17394_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10149__B _12130_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19133_ _19137_/CLK _19133_/D repeater249/X vssd1 vssd1 vccd1 vccd1 _19133_/Q sky130_fd_sc_hd__dfrtp_1
X_16345_ _17346_/X _16415_/B vssd1 vssd1 vccd1 vccd1 _16345_/X sky130_fd_sc_hd__and2_1
X_13557_ _13557_/A _13557_/B vssd1 vssd1 vccd1 vccd1 _13558_/A sky130_fd_sc_hd__or2_1
XFILLER_9_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10769_ _19751_/Q _10767_/B _10758_/B _10767_/Y vssd1 vssd1 vccd1 vccd1 _19751_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_12_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12508_ _19081_/Q _12505_/X _12404_/X _12506_/X vssd1 vssd1 vccd1 vccd1 _19081_/D
+ sky130_fd_sc_hd__a22o_1
X_19064_ _19585_/CLK _19064_/D hold361/X vssd1 vssd1 vccd1 vccd1 _19064_/Q sky130_fd_sc_hd__dfrtp_1
X_13488_ _13483_/A _13483_/B _13483_/C vssd1 vssd1 vccd1 vccd1 _13489_/B sky130_fd_sc_hd__o21a_1
X_16276_ _18095_/Q vssd1 vssd1 vccd1 vccd1 _16276_/Y sky130_fd_sc_hd__inv_2
XFILLER_172_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18015_ _18169_/CLK _18015_/D vssd1 vssd1 vccd1 vccd1 _18015_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__18845__RESET_B repeater233/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15227_ _19723_/Q vssd1 vssd1 vccd1 vccd1 _15227_/Y sky130_fd_sc_hd__inv_2
XFILLER_145_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17647__S _17655_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12439_ _15769_/A _12487_/B vssd1 vssd1 vccd1 vccd1 _12478_/A sky130_fd_sc_hd__or2_4
XFILLER_172_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12194__B1 _12074_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15158_ _15159_/A vssd1 vssd1 vccd1 vccd1 _15158_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_5_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20043__CLK _20051_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14109_ _18697_/Q _14108_/Y _14096_/X _14109_/C1 vssd1 vssd1 vccd1 vccd1 _18697_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_141_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12380__A hold291/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15089_ _17998_/Q _15083_/X _14791_/X _15085_/X vssd1 vssd1 vccd1 vccd1 _17998_/D
+ sky130_fd_sc_hd__a22o_1
X_19966_ _19976_/CLK _19966_/D repeater185/X vssd1 vssd1 vccd1 vccd1 _19966_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_101_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18917_ _19293_/CLK _18917_/D repeater187/X vssd1 vssd1 vccd1 vccd1 _18917_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__13694__A0 _12313_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19897_ _19900_/CLK _19897_/D repeater195/X vssd1 vssd1 vccd1 vccd1 _19897_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_79_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17382__S _17414_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09650_ _19993_/Q vssd1 vssd1 vccd1 vccd1 _09749_/A sky130_fd_sc_hd__inv_2
X_18848_ _18866_/CLK _18848_/D repeater232/X vssd1 vssd1 vccd1 vccd1 _18848_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_228_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09581_ _09585_/A vssd1 vssd1 vccd1 vccd1 _09581_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_67_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18779_ _19667_/CLK _18779_/D repeater264/X vssd1 vssd1 vccd1 vccd1 _18779_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_243_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19633__RESET_B repeater258/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11724__A _11731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17807__S0 _17918_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16396__C1 _16393_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_224_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19409__CLK _19984_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_opt_3_HCLK clkbuf_opt_3_HCLK/A vssd1 vssd1 vccd1 vccd1 _18506_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_192_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09015_ _09041_/A vssd1 vssd1 vccd1 vccd1 _09015_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_164_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18586__RESET_B repeater272/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold130 input14/X vssd1 vssd1 vccd1 vccd1 hold130/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09050__B1 _09049_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold141 hold141/A vssd1 vssd1 vccd1 vccd1 hold141/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold152 HSEL vssd1 vssd1 vccd1 vccd1 input35/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 HADDR[11] vssd1 vssd1 vccd1 vccd1 input3/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold174 input4/X vssd1 vssd1 vccd1 vccd1 hold174/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 hold185/A vssd1 vssd1 vccd1 vccd1 hold185/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold196 input27/X vssd1 vssd1 vccd1 vccd1 hold196/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_160_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20106_ _20107_/CLK _20106_/D repeater230/X vssd1 vssd1 vccd1 vccd1 _20106_/Q sky130_fd_sc_hd__dfrtp_4
X_09917_ _19334_/Q vssd1 vssd1 vccd1 vccd1 _09917_/Y sky130_fd_sc_hd__inv_2
XFILLER_132_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17292__S _17513_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20037_ _20064_/CLK _20037_/D repeater198/X vssd1 vssd1 vccd1 vccd1 _20037_/Q sky130_fd_sc_hd__dfrtp_2
X_09848_ _09848_/A _09848_/B vssd1 vssd1 vccd1 vccd1 _10001_/A sky130_fd_sc_hd__or2_2
XFILLER_85_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09779_ _19989_/Q _09778_/Y _09763_/X _09746_/B vssd1 vssd1 vccd1 vccd1 _19989_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_4112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19374__RESET_B repeater241/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11810_ _19454_/Q _11807_/X _09058_/X _11808_/X vssd1 vssd1 vccd1 vccd1 _19454_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12790_ _19232_/Q vssd1 vssd1 vccd1 vccd1 _12790_/Y sky130_fd_sc_hd__inv_2
XFILLER_160_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11741_ _15749_/A _11737_/X _16930_/X _11738_/X vssd1 vssd1 vccd1 vccd1 _19498_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09104__A _14780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_152_HCLK_A clkbuf_4_1_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11672_ _15311_/A _11672_/B _11672_/C vssd1 vssd1 vccd1 vccd1 _11672_/Y sky130_fd_sc_hd__nor3_4
XFILLER_159_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14460_ _18363_/Q _14452_/A _14403_/X _14453_/A vssd1 vssd1 vccd1 vccd1 _18363_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10623_ _19808_/Q _10609_/A _10575_/A _10606_/X vssd1 vssd1 vccd1 vccd1 _19808_/D
+ sky130_fd_sc_hd__o22a_1
X_13411_ _20108_/Q _13429_/B _13410_/Y _18858_/Q vssd1 vssd1 vccd1 vccd1 _13411_/X
+ sky130_fd_sc_hd__o2bb2a_1
XPHY_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14391_ _18755_/Q vssd1 vssd1 vccd1 vccd1 _14731_/B sky130_fd_sc_hd__buf_1
XPHY_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13342_ _13429_/A _13342_/B vssd1 vssd1 vccd1 vccd1 _13450_/A sky130_fd_sc_hd__or2_1
X_16130_ _16125_/Y _15866_/A _16126_/Y _15840_/A _16129_/X vssd1 vssd1 vccd1 vccd1
+ _16130_/X sky130_fd_sc_hd__o221a_1
X_10554_ _19805_/Q vssd1 vssd1 vccd1 vccd1 _10558_/B sky130_fd_sc_hd__inv_2
XFILLER_210_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17467__S _17568_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16061_ _18874_/Q vssd1 vssd1 vccd1 vccd1 _16061_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14165__B2 _14003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13273_ _18754_/Q vssd1 vssd1 vccd1 vccd1 _14270_/A sky130_fd_sc_hd__inv_2
XANTENNA__15776__A _15776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10485_ _19544_/Q _19543_/Q vssd1 vssd1 vccd1 vccd1 _10501_/C sky130_fd_sc_hd__or2_1
XFILLER_154_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12176__B1 _11920_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12224_ _19236_/Q _12219_/X _12223_/X _12220_/X vssd1 vssd1 vccd1 vccd1 _19236_/D
+ sky130_fd_sc_hd__a22o_1
X_15012_ _15012_/A vssd1 vssd1 vccd1 vccd1 _15012_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__11923__B1 _11922_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19820_ _19822_/CLK _19820_/D repeater218/X vssd1 vssd1 vccd1 vccd1 _19820_/Q sky130_fd_sc_hd__dfrtp_1
X_12155_ _19280_/Q _12150_/X _12102_/X _12151_/X vssd1 vssd1 vccd1 vccd1 _19280_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16862__A0 _17473_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11106_ _11106_/A vssd1 vssd1 vccd1 vccd1 _17754_/S sky130_fd_sc_hd__inv_2
XFILLER_96_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19751_ _20070_/CLK _19751_/D repeater197/X vssd1 vssd1 vccd1 vccd1 _19751_/Q sky130_fd_sc_hd__dfrtp_1
X_16963_ _16647_/Y _16963_/A1 _17529_/S vssd1 vssd1 vccd1 vccd1 _16963_/X sky130_fd_sc_hd__mux2_1
X_12086_ hold308/X vssd1 vssd1 vccd1 vccd1 _12086_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__10432__B _15199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18702_ _19119_/CLK _18702_/D hold351/X vssd1 vssd1 vccd1 vccd1 _18702_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_204_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11037_ _19649_/Q _11029_/Y _19649_/Q _11029_/Y vssd1 vssd1 vccd1 vccd1 _19649_/D
+ sky130_fd_sc_hd__o2bb2a_1
X_15914_ _15914_/A vssd1 vssd1 vccd1 vccd1 _15915_/A sky130_fd_sc_hd__buf_1
X_19682_ _19795_/CLK _19682_/D repeater219/X vssd1 vssd1 vccd1 vccd1 _19682_/Q sky130_fd_sc_hd__dfrtp_1
X_16894_ _16893_/X _13089_/A _17488_/S vssd1 vssd1 vccd1 vccd1 _16894_/X sky130_fd_sc_hd__mux2_1
XFILLER_237_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18633_ _18633_/CLK _18633_/D repeater225/X vssd1 vssd1 vccd1 vccd1 _18633_/Q sky130_fd_sc_hd__dfrtp_4
X_15845_ _15858_/A _15858_/B _15858_/C _15845_/D vssd1 vssd1 vccd1 vccd1 _15846_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_225_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18564_ _19841_/CLK _18564_/D repeater194/X vssd1 vssd1 vccd1 vccd1 _18564_/Q sky130_fd_sc_hd__dfrtp_1
X_15776_ _15776_/A vssd1 vssd1 vccd1 vccd1 _17537_/S sky130_fd_sc_hd__clkinv_4
XFILLER_220_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12988_ _12988_/A vssd1 vssd1 vccd1 vccd1 _12988_/Y sky130_fd_sc_hd__inv_2
XFILLER_206_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09014__A _09084_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17515_ _17514_/X _10109_/Y _17548_/S vssd1 vssd1 vccd1 vccd1 _17515_/X sky130_fd_sc_hd__mux2_1
X_14727_ _14727_/A vssd1 vssd1 vccd1 vccd1 _14727_/X sky130_fd_sc_hd__clkbuf_2
X_11939_ _11955_/A vssd1 vssd1 vccd1 vccd1 _11939_/X sky130_fd_sc_hd__buf_1
X_18495_ _20089_/CLK _18495_/D repeater203/X vssd1 vssd1 vccd1 vccd1 _18495_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_221_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17446_ _15963_/X _09513_/Y _17534_/S vssd1 vssd1 vccd1 vccd1 _17446_/X sky130_fd_sc_hd__mux2_1
XFILLER_221_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14658_ _14658_/A vssd1 vssd1 vccd1 vccd1 _14658_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_60_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13609_ _13530_/A _13530_/B _13588_/A _13607_/Y vssd1 vssd1 vccd1 vccd1 _18806_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_20_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12403__A1 _19147_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_11_HCLK_A clkbuf_4_2_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17377_ _17376_/X _17864_/X _17568_/S vssd1 vssd1 vccd1 vccd1 _17377_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09668__B _09807_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14589_ _14589_/A vssd1 vssd1 vccd1 vccd1 _14589_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__12375__A hold284/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_74_HCLK_A clkbuf_opt_4_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19116_ _19119_/CLK _19116_/D hold353/X vssd1 vssd1 vccd1 vccd1 _19116_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_174_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16328_ _18144_/Q vssd1 vssd1 vccd1 vccd1 _16328_/Y sky130_fd_sc_hd__inv_2
XFILLER_158_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17342__A1 _18778_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17377__S _17568_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19047_ _19566_/CLK _19047_/D repeater255/X vssd1 vssd1 vccd1 vccd1 _19047_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_173_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16259_ _18055_/Q vssd1 vssd1 vccd1 vccd1 _16259_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12167__B1 _12038_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09032__B1 _09030_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19851__CLK _19851_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13667__B1 hold267/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19949_ _19964_/CLK _19949_/D hold371/X vssd1 vssd1 vccd1 vccd1 _19949_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_228_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09702_ _09791_/A _19408_/Q _19979_/Q _09700_/Y _09701_/X vssd1 vssd1 vccd1 vccd1
+ _09703_/D sky130_fd_sc_hd__o221a_1
XFILLER_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09633_ _19974_/Q vssd1 vssd1 vccd1 vccd1 _09635_/B sky130_fd_sc_hd__inv_2
XFILLER_215_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09564_ _09564_/A _09564_/B _09564_/C _09564_/D vssd1 vssd1 vccd1 vccd1 _09565_/D
+ sky130_fd_sc_hd__and4_1
XANTENNA__09099__B1 _09098_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09495_ _09495_/A vssd1 vssd1 vccd1 vccd1 _09495_/Y sky130_fd_sc_hd__inv_2
XPHY_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18767__RESET_B repeater271/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17287__S _17545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16541__C1 _16540_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10270_ _14517_/A _10269_/X _14517_/A _10269_/X vssd1 vssd1 vccd1 vccd1 _10281_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_105_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19555__RESET_B hold348/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13960_ _13960_/A vssd1 vssd1 vccd1 vccd1 _13960_/Y sky130_fd_sc_hd__inv_2
XFILLER_47_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12330__B1 _12086_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12911_ _19281_/Q vssd1 vssd1 vccd1 vccd1 _12911_/Y sky130_fd_sc_hd__inv_4
XFILLER_235_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13891_ _19198_/Q vssd1 vssd1 vccd1 vccd1 _13891_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16072__A1 _17448_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_234_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15630_ _18600_/Q _15621_/A _18601_/Q vssd1 vssd1 vccd1 vccd1 _15630_/X sky130_fd_sc_hd__o21a_1
XFILLER_234_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12842_ _18942_/Q vssd1 vssd1 vccd1 vccd1 _12967_/C sky130_fd_sc_hd__inv_2
XFILLER_62_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_131_HCLK clkbuf_4_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19137_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_199_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15561_ _18584_/Q vssd1 vssd1 vccd1 vccd1 _15561_/Y sky130_fd_sc_hd__inv_2
XFILLER_199_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12773_ _18832_/Q vssd1 vssd1 vccd1 vccd1 _13555_/A sky130_fd_sc_hd__inv_2
XPHY_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17300_ _17299_/X _13358_/Y _17535_/S vssd1 vssd1 vccd1 vccd1 _17300_/X sky130_fd_sc_hd__mux2_1
XPHY_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18479__CLK _19780_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14512_ _18333_/Q _14503_/X hold330/X _14505_/X vssd1 vssd1 vccd1 vccd1 _18333_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_203_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11724_ _11731_/A vssd1 vssd1 vccd1 vccd1 _11724_/X sky130_fd_sc_hd__buf_1
X_18280_ _19847_/CLK _18280_/D vssd1 vssd1 vccd1 vccd1 _18280_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_202_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15492_ _15490_/Y _15491_/Y _15483_/X vssd1 vssd1 vccd1 vccd1 _15492_/X sky130_fd_sc_hd__o21a_1
XANTENNA__17572__A1 _19771_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17231_ _15768_/Y _11294_/Y _17546_/S vssd1 vssd1 vccd1 vccd1 _17231_/X sky130_fd_sc_hd__mux2_1
XFILLER_80_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11655_ _11655_/A _11655_/B vssd1 vssd1 vccd1 vccd1 _11655_/X sky130_fd_sc_hd__or2_1
X_14443_ _14751_/A vssd1 vssd1 vccd1 vccd1 _14443_/X sky130_fd_sc_hd__clkbuf_2
XPHY_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10708__A hold336/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12397__B1 _12396_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10606_ _10606_/A vssd1 vssd1 vccd1 vccd1 _10606_/X sky130_fd_sc_hd__clkbuf_2
X_17162_ _16547_/Y _19380_/Q _17385_/S vssd1 vssd1 vccd1 vccd1 _17162_/X sky130_fd_sc_hd__mux2_1
XFILLER_168_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11586_ _11586_/A vssd1 vssd1 vccd1 vccd1 _11586_/Y sky130_fd_sc_hd__inv_2
X_14374_ _18413_/Q _14367_/X _14326_/X _14369_/X vssd1 vssd1 vccd1 vccd1 _18413_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17197__S _17546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16113_ _18770_/Q vssd1 vssd1 vccd1 vccd1 _16113_/Y sky130_fd_sc_hd__inv_2
X_10537_ _10537_/A _10537_/B vssd1 vssd1 vccd1 vccd1 _10537_/Y sky130_fd_sc_hd__nor2_1
X_13325_ _18842_/Q vssd1 vssd1 vccd1 vccd1 _13465_/A sky130_fd_sc_hd__inv_2
XFILLER_128_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17093_ _15768_/Y _14199_/Y _17546_/S vssd1 vssd1 vccd1 vccd1 _17093_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12149__B1 _12092_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16044_ _17939_/Q _16096_/B vssd1 vssd1 vccd1 vccd1 _16044_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__15886__B2 _15858_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10468_ _19823_/Q vssd1 vssd1 vccd1 vccd1 _10468_/Y sky130_fd_sc_hd__inv_2
X_13256_ _18751_/Q vssd1 vssd1 vccd1 vccd1 _13256_/X sky130_fd_sc_hd__buf_1
XFILLER_108_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12207_ _19248_/Q _12205_/X _12095_/X _12206_/X vssd1 vssd1 vccd1 vccd1 _19248_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_89_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13187_ _13187_/A vssd1 vssd1 vccd1 vccd1 _13187_/Y sky130_fd_sc_hd__inv_2
X_10399_ _11096_/A _14476_/A vssd1 vssd1 vccd1 vccd1 _10400_/B sky130_fd_sc_hd__or2_1
XFILLER_97_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16835__A0 _17486_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19803_ _19812_/CLK _19803_/D repeater222/X vssd1 vssd1 vccd1 vccd1 _19803_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_111_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12138_ _19293_/Q _12134_/X _12069_/X _12137_/X vssd1 vssd1 vccd1 vccd1 _19293_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_229_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17995_ _18465_/CLK _17995_/D vssd1 vssd1 vccd1 vccd1 _17995_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19296__RESET_B repeater241/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19734_ _20051_/CLK _19734_/D repeater207/X vssd1 vssd1 vccd1 vccd1 _19734_/Q sky130_fd_sc_hd__dfrtp_1
X_16946_ _19490_/Q hold171/X _16946_/S vssd1 vssd1 vccd1 vccd1 _16946_/X sky130_fd_sc_hd__mux2_1
X_12069_ hold284/X vssd1 vssd1 vccd1 vccd1 _12069_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_237_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19225__RESET_B repeater257/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19665_ _19855_/CLK _19665_/D repeater264/X vssd1 vssd1 vccd1 vccd1 _19665_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_49_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16877_ _16876_/X _09414_/Y _17529_/S vssd1 vssd1 vccd1 vccd1 _16877_/X sky130_fd_sc_hd__mux2_1
X_18616_ _19577_/CLK _18616_/D repeater268/X vssd1 vssd1 vccd1 vccd1 _18616_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_37_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15828_ _15828_/A vssd1 vssd1 vccd1 vccd1 _15828_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__10883__B1 _10882_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_231_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19596_ _19597_/CLK _19596_/D hold273/X vssd1 vssd1 vccd1 vccd1 _19596_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_80_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18547_ _19814_/CLK _18547_/D repeater220/X vssd1 vssd1 vccd1 vccd1 _18547_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_64_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15759_ _18886_/Q _18884_/Q _18885_/Q _15758_/X vssd1 vssd1 vccd1 vccd1 _18525_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12624__A1 _19018_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17012__A0 _17473_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09280_ _19499_/Q vssd1 vssd1 vccd1 vccd1 _15749_/C sky130_fd_sc_hd__clkbuf_2
X_18478_ _19780_/CLK _19684_/Q repeater227/X vssd1 vssd1 vccd1 vccd1 _18478_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17563__A1 _17909_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18860__RESET_B repeater232/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17429_ _16116_/Y _16114_/Y _17564_/S vssd1 vssd1 vccd1 vccd1 _17429_/X sky130_fd_sc_hd__mux2_1
XFILLER_221_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09253__A0 _18652_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_12_HCLK clkbuf_4_2_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _18765_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_114_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15863__B _15863_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08995_ _19516_/Q _09259_/B _10250_/C vssd1 vssd1 vccd1 vccd1 _13279_/C sky130_fd_sc_hd__or3_4
XFILLER_88_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_154_HCLK clkbuf_4_1_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _18435_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_84_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11184__A _11191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09616_ _20007_/Q _09615_/Y _09585_/A _09616_/C1 vssd1 vssd1 vccd1 vccd1 _20007_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_141_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19747__CLK _20070_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_243_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09547_ _19306_/Q vssd1 vssd1 vccd1 vccd1 _09547_/Y sky130_fd_sc_hd__inv_2
XFILLER_71_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17003__A0 _17473_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09478_ _09478_/A _09478_/B vssd1 vssd1 vccd1 vccd1 _09595_/A sky130_fd_sc_hd__or2_1
XPHY_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16914__S _17386_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19897__CLK _19900_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12379__B1 _12375_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11440_ _19549_/Q vssd1 vssd1 vccd1 vccd1 _11548_/A sky130_fd_sc_hd__inv_2
XFILLER_196_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11371_ _19549_/Q _11366_/Y _11547_/A _19154_/Q _11370_/Y vssd1 vssd1 vccd1 vccd1
+ _11389_/A sky130_fd_sc_hd__o221a_1
XFILLER_137_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10322_ _10322_/A _10375_/A vssd1 vssd1 vccd1 vccd1 _10371_/A sky130_fd_sc_hd__or2_1
X_13110_ _19160_/Q vssd1 vssd1 vccd1 vccd1 _13110_/Y sky130_fd_sc_hd__inv_2
X_14090_ _19062_/Q vssd1 vssd1 vccd1 vccd1 _14090_/Y sky130_fd_sc_hd__inv_2
XFILLER_166_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19736__RESET_B repeater208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13041_ _18905_/Q vssd1 vssd1 vccd1 vccd1 _13077_/A sky130_fd_sc_hd__inv_2
X_10253_ _19498_/Q _19497_/Q _10430_/A vssd1 vssd1 vccd1 vccd1 _15823_/A sky130_fd_sc_hd__or3_4
XFILLER_124_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10263__A _19647_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10184_ _19877_/Q _10181_/A _10290_/B vssd1 vssd1 vccd1 vccd1 _19877_/D sky130_fd_sc_hd__a21o_1
XFILLER_182_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16800_ _16799_/X _18916_/Q _17542_/S vssd1 vssd1 vccd1 vccd1 _16800_/X sky130_fd_sc_hd__mux2_1
XFILLER_182_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17780_ _18317_/Q _18437_/Q _18429_/Q _18421_/Q _17923_/S0 _19646_/Q vssd1 vssd1
+ vccd1 vccd1 _17780_/X sky130_fd_sc_hd__mux4_1
XFILLER_47_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14992_ _18959_/Q vssd1 vssd1 vccd1 vccd1 _14992_/X sky130_fd_sc_hd__buf_2
XANTENNA__12303__B1 _12302_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16731_ _16774_/X _16493_/A _16777_/X _16512_/A vssd1 vssd1 vccd1 vccd1 _16731_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_59_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13943_ _13909_/D _13815_/B _13941_/Y _13919_/X vssd1 vssd1 vccd1 vccd1 _18716_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_47_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17480__S _17534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19450_ _19841_/CLK _19450_/D repeater271/X vssd1 vssd1 vccd1 vccd1 _19450_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_19_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16662_ _17014_/X _16637_/X _17043_/X _16638_/X vssd1 vssd1 vccd1 vccd1 _16662_/X
+ sky130_fd_sc_hd__o22a_1
X_13874_ _13846_/Y _18705_/Q _13871_/Y _18727_/Q _13873_/X vssd1 vssd1 vccd1 vccd1
+ _13882_/B sky130_fd_sc_hd__o221a_1
XFILLER_235_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18401_ _19637_/CLK _18401_/D vssd1 vssd1 vccd1 vccd1 _18401_/Q sky130_fd_sc_hd__dfxtp_1
X_15613_ _18596_/Q _15605_/A _18597_/Q vssd1 vssd1 vccd1 vccd1 _15613_/X sky130_fd_sc_hd__o21a_1
X_19381_ _19927_/CLK _19381_/D repeater230/X vssd1 vssd1 vccd1 vccd1 _19381_/Q sky130_fd_sc_hd__dfrtp_1
X_12825_ _19235_/Q _13536_/A _19252_/Q _13552_/A vssd1 vssd1 vccd1 vccd1 _12825_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__18689__RESET_B hold359/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16593_ _17252_/X _16555_/X _17247_/X _16556_/X vssd1 vssd1 vccd1 vccd1 _16600_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_201_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_repeater185_A hold371/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18332_ _18333_/CLK _18332_/D vssd1 vssd1 vccd1 vccd1 _18332_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__18618__RESET_B repeater269/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15544_ _18580_/Q vssd1 vssd1 vccd1 vccd1 _15544_/Y sky130_fd_sc_hd__inv_2
XFILLER_91_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12756_ _16719_/A _18833_/Q _19234_/Q _13535_/A vssd1 vssd1 vccd1 vccd1 _12756_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11707_ _11737_/A vssd1 vssd1 vccd1 vccd1 _11730_/A sky130_fd_sc_hd__buf_2
X_18263_ _20077_/CLK _18263_/D vssd1 vssd1 vccd1 vccd1 _18263_/Q sky130_fd_sc_hd__dfxtp_1
X_15475_ _15475_/A _15475_/B vssd1 vssd1 vccd1 vccd1 _15475_/Y sky130_fd_sc_hd__nor2_1
XFILLER_129_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16824__S _17482_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12687_ _18975_/Q _12684_/X hold233/X _12685_/X vssd1 vssd1 vccd1 vccd1 _18975_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17214_ _17213_/X _09857_/B _17524_/S vssd1 vssd1 vccd1 vccd1 _17214_/X sky130_fd_sc_hd__mux2_1
XFILLER_147_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14426_ _14426_/A vssd1 vssd1 vccd1 vccd1 _14426_/X sky130_fd_sc_hd__clkbuf_2
XPHY_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11638_ _19550_/Q _11641_/A _11635_/A _11563_/X vssd1 vssd1 vccd1 vccd1 _19550_/D
+ sky130_fd_sc_hd__o211a_1
X_18194_ _18333_/CLK _18194_/D vssd1 vssd1 vccd1 vccd1 _18194_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_35_HCLK _18641_/CLK vssd1 vssd1 vccd1 vccd1 _20077_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17145_ _17144_/X _09453_/Y _17529_/S vssd1 vssd1 vccd1 vccd1 _17145_/X sky130_fd_sc_hd__mux2_1
X_14357_ _18424_/Q _14349_/X _14356_/X _14353_/X vssd1 vssd1 vccd1 vccd1 _18424_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_128_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11569_ _11569_/A _11569_/B _11569_/C vssd1 vssd1 vccd1 vccd1 _19576_/D sky130_fd_sc_hd__nor3_1
X_13308_ _18857_/Q vssd1 vssd1 vccd1 vccd1 _13428_/B sky130_fd_sc_hd__inv_2
X_17076_ _17075_/X _19148_/Q _17548_/S vssd1 vssd1 vccd1 vccd1 _17076_/X sky130_fd_sc_hd__mux2_2
X_14288_ _14289_/A vssd1 vssd1 vccd1 vccd1 _14288_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__16520__A2 _15904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17655__S _17655_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16027_ _18092_/Q vssd1 vssd1 vccd1 vccd1 _16027_/Y sky130_fd_sc_hd__inv_2
X_13239_ _15404_/A vssd1 vssd1 vccd1 vccd1 _15419_/A sky130_fd_sc_hd__buf_2
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12542__B1 _12541_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19406__RESET_B repeater210/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17978_ _20123_/CLK _17978_/D vssd1 vssd1 vccd1 vccd1 _17978_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14295__B1 _13676_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19717_ _19720_/CLK _19717_/D repeater202/X vssd1 vssd1 vccd1 vccd1 _19717_/Q sky130_fd_sc_hd__dfrtp_2
X_16929_ _19473_/Q hold199/X _16950_/S vssd1 vssd1 vccd1 vccd1 _16929_/X sky130_fd_sc_hd__mux2_4
XFILLER_66_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17390__S _17545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19648_ _19859_/CLK _19648_/D repeater262/X vssd1 vssd1 vccd1 vccd1 _19648_/Q sky130_fd_sc_hd__dfrtp_2
X_09401_ _19385_/Q vssd1 vssd1 vccd1 vccd1 _09401_/Y sky130_fd_sc_hd__inv_2
XFILLER_225_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19579_ _19600_/CLK _19579_/D hold355/X vssd1 vssd1 vccd1 vccd1 _19579_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_41_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09332_ _09313_/Y _09315_/Y _20047_/Q _15725_/A _09331_/X vssd1 vssd1 vccd1 vccd1
+ _09332_/X sky130_fd_sc_hd__o221a_1
XFILLER_40_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09263_ _14245_/C vssd1 vssd1 vccd1 vccd1 _15961_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_193_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09194_ _20072_/Q _09192_/Y _09192_/B _09193_/Y vssd1 vssd1 vccd1 vccd1 _20072_/D
+ sky130_fd_sc_hd__o22a_1
XANTENNA__15858__B _15858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18174__CLK _18198_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17565__S _17565_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08978_ _08978_/A _09199_/A vssd1 vssd1 vccd1 vccd1 _10133_/C sky130_fd_sc_hd__or2_1
XFILLER_29_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold278_A HWDATA[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_229_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16909__S _17542_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10847__B1 _10448_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10940_ _10940_/A vssd1 vssd1 vccd1 vccd1 _10940_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_217_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10871_ _19701_/Q _10856_/A _10870_/X _10857_/A vssd1 vssd1 vccd1 vccd1 _19701_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17870__S1 _19632_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12610_ _12313_/X _19024_/Q _12610_/S vssd1 vssd1 vccd1 vccd1 _19024_/D sky130_fd_sc_hd__mux2_1
XPHY_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18711__RESET_B repeater253/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13590_ _13590_/A vssd1 vssd1 vccd1 vccd1 _13590_/Y sky130_fd_sc_hd__inv_2
XPHY_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_58_HCLK clkbuf_4_12_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19905_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12541_ hold335/X vssd1 vssd1 vccd1 vccd1 _12541_/X sky130_fd_sc_hd__buf_6
XFILLER_40_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10258__A _15296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_opt_2_HCLK_A clkbuf_opt_2_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15260_ _15268_/A _19777_/Q _15257_/Y _15259_/Y vssd1 vssd1 vccd1 vccd1 _15260_/X
+ sky130_fd_sc_hd__a31o_1
XPHY_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19988__RESET_B repeater192/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12472_ _12479_/A vssd1 vssd1 vccd1 vccd1 _12472_/X sky130_fd_sc_hd__buf_1
XFILLER_184_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14211_ _19123_/Q vssd1 vssd1 vccd1 vccd1 _14211_/Y sky130_fd_sc_hd__inv_2
XFILLER_184_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11423_ _19152_/Q vssd1 vssd1 vccd1 vccd1 _11423_/Y sky130_fd_sc_hd__inv_2
X_15191_ _15191_/A vssd1 vssd1 vccd1 vccd1 _17764_/S sky130_fd_sc_hd__inv_2
XFILLER_153_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11354_ _18972_/Q vssd1 vssd1 vccd1 vccd1 _11354_/Y sky130_fd_sc_hd__inv_2
X_14142_ _14142_/A vssd1 vssd1 vccd1 vccd1 _14142_/Y sky130_fd_sc_hd__clkinv_1
X_10305_ _18603_/Q _18602_/Q _15629_/A vssd1 vssd1 vccd1 vccd1 _15640_/B sky130_fd_sc_hd__or3_4
XANTENNA__17475__S _17517_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11285_ _19583_/Q _11280_/Y _19598_/Q _16615_/A _11284_/X vssd1 vssd1 vccd1 vccd1
+ _11298_/B sky130_fd_sc_hd__o221a_1
X_14073_ _19086_/Q vssd1 vssd1 vccd1 vccd1 _14073_/Y sky130_fd_sc_hd__inv_2
X_18950_ _19290_/CLK _18950_/D repeater211/X vssd1 vssd1 vccd1 vccd1 _18950_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_153_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13298__A1_N _18752_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12524__B1 hold267/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17901_ _15923_/Y _15924_/Y _15925_/Y _15926_/Y _17913_/S0 _19632_/Q vssd1 vssd1
+ vccd1 vccd1 _17901_/X sky130_fd_sc_hd__mux4_2
X_10236_ _19834_/Q vssd1 vssd1 vccd1 vccd1 _10236_/Y sky130_fd_sc_hd__inv_2
X_13024_ _13024_/A vssd1 vssd1 vccd1 vccd1 _13027_/A sky130_fd_sc_hd__inv_2
X_18881_ _19814_/CLK _18881_/D repeater220/X vssd1 vssd1 vccd1 vccd1 _18881_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_121_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17832_ _18360_/Q _18000_/Q _18416_/Q _18400_/Q _17918_/S0 _18750_/Q vssd1 vssd1
+ vccd1 vccd1 _17832_/X sky130_fd_sc_hd__mux4_2
XFILLER_126_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10167_ _10174_/A vssd1 vssd1 vccd1 vccd1 _10175_/A sky130_fd_sc_hd__inv_2
XFILLER_208_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17763_ _15192_/Y _13289_/Y _17763_/S vssd1 vssd1 vccd1 vccd1 _17763_/X sky130_fd_sc_hd__mux2_1
X_10098_ _19911_/Q _10097_/Y _10084_/B _10026_/X vssd1 vssd1 vccd1 vccd1 _19911_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_66_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14975_ _15082_/A _14975_/B _14975_/C vssd1 vssd1 vccd1 vccd1 _14978_/A sky130_fd_sc_hd__or3_4
XANTENNA__16819__S _17543_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19502_ _19510_/CLK hold229/X repeater256/X vssd1 vssd1 vccd1 vccd1 _19502_/Q sky130_fd_sc_hd__dfrtp_1
X_16714_ _16844_/X _16687_/X _16896_/X _16688_/X _16713_/X vssd1 vssd1 vccd1 vccd1
+ _16715_/C sky130_fd_sc_hd__o221a_1
XFILLER_212_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13926_ _18727_/Q _13924_/Y _13827_/B _13925_/X vssd1 vssd1 vccd1 vccd1 _18727_/D
+ sky130_fd_sc_hd__o211a_1
X_17694_ _15455_/Y _19441_/Q _17696_/S vssd1 vssd1 vccd1 vccd1 _18558_/D sky130_fd_sc_hd__mux2_1
X_19433_ _19513_/CLK _19433_/D repeater259/X vssd1 vssd1 vccd1 vccd1 _19433_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_207_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16645_ _16645_/A _16647_/B vssd1 vssd1 vccd1 vccd1 _16645_/Y sky130_fd_sc_hd__nor2_1
XFILLER_62_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13857_ _19201_/Q _13949_/A _13855_/Y _18712_/Q _13856_/X vssd1 vssd1 vccd1 vccd1
+ _13867_/B sky130_fd_sc_hd__o221a_1
XANTENNA__17861__S1 _19632_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12808_ _12808_/A _12808_/B _12808_/C _12808_/D vssd1 vssd1 vccd1 vccd1 _12834_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_90_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19364_ _19984_/CLK _19364_/D repeater243/X vssd1 vssd1 vccd1 vccd1 _19364_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__09456__B1 _10039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16576_ _17123_/X _16573_/X _17111_/X _16574_/X _16575_/X vssd1 vssd1 vccd1 vccd1
+ _16581_/B sky130_fd_sc_hd__o221a_4
XFILLER_222_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13788_ _18724_/Q vssd1 vssd1 vccd1 vccd1 _13909_/B sky130_fd_sc_hd__inv_2
XFILLER_188_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18315_ _18435_/CLK _18315_/D vssd1 vssd1 vccd1 vccd1 _18315_/Q sky130_fd_sc_hd__dfxtp_1
X_15527_ _15525_/Y _15526_/Y _15512_/X vssd1 vssd1 vccd1 vccd1 _15527_/X sky130_fd_sc_hd__o21a_1
X_12739_ _12734_/Y _18835_/Q _19236_/Q _13537_/B _12738_/X vssd1 vssd1 vccd1 vccd1
+ _12758_/A sky130_fd_sc_hd__o221a_1
X_19295_ _20115_/CLK _19295_/D repeater239/X vssd1 vssd1 vccd1 vccd1 _19295_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_187_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18246_ _19847_/CLK _18246_/D vssd1 vssd1 vccd1 vccd1 _18246_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__19712__SET_B repeater219/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15458_ _18558_/Q _15453_/A _18559_/Q vssd1 vssd1 vccd1 vccd1 _15458_/X sky130_fd_sc_hd__o21a_1
XANTENNA__16741__A2 _16513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14409_ _14410_/A vssd1 vssd1 vccd1 vccd1 _14409_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__19658__RESET_B repeater270/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18177_ _18216_/CLK _18177_/D vssd1 vssd1 vccd1 vccd1 _18177_/Q sky130_fd_sc_hd__dfxtp_1
X_15389_ _15389_/A _15389_/B _15389_/C vssd1 vssd1 vccd1 vccd1 _18519_/D sky130_fd_sc_hd__and3_1
XFILLER_117_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17128_ _17127_/X _09720_/Y _17517_/S vssd1 vssd1 vccd1 vccd1 _17128_/X sky130_fd_sc_hd__mux2_1
XANTENNA__17385__S _17385_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17059_ _16668_/Y _20115_/Q _17385_/S vssd1 vssd1 vccd1 vccd1 _17059_/X sky130_fd_sc_hd__mux2_1
X_09950_ _09968_/A vssd1 vssd1 vccd1 vccd1 _09950_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_leaf_129_HCLK_A clkbuf_4_4_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19240__RESET_B repeater239/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12515__B1 _12344_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20070_ _20070_/CLK _20070_/D repeater207/X vssd1 vssd1 vccd1 vccd1 _20070_/Q sky130_fd_sc_hd__dfrtp_1
X_09881_ _09856_/A _19339_/Q _09864_/A _19348_/Q vssd1 vssd1 vccd1 vccd1 _09881_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_140_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17206__A0 _15963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_214_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17852__S1 _19632_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12558__A _12659_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17509__A1 _15610_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14440__B1 _14437_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09315_ _15725_/A vssd1 vssd1 vccd1 vccd1 _09315_/Y sky130_fd_sc_hd__inv_2
XFILLER_210_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09246_ _20065_/Q _20066_/Q _09250_/S vssd1 vssd1 vccd1 vccd1 _20066_/D sky130_fd_sc_hd__mux2_1
XFILLER_194_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19399__RESET_B repeater271/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09177_ _14707_/A vssd1 vssd1 vccd1 vccd1 _09177_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_175_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19328__RESET_B repeater241/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17295__S _17541_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11309__B2 _18977_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11070_ _17754_/X vssd1 vssd1 vccd1 vccd1 _11070_/Y sky130_fd_sc_hd__inv_2
XFILLER_150_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput79 _15918_/Y vssd1 vssd1 vccd1 vccd1 HRDATA[0] sky130_fd_sc_hd__clkbuf_2
XANTENNA__16212__B _16212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10021_ _10033_/B _10021_/B _10021_/C vssd1 vssd1 vccd1 vccd1 _10051_/A sky130_fd_sc_hd__or3_1
XFILLER_49_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16248__B2 _15999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09107__A hold322/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10280__A1_N _19646_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14760_ _14760_/A vssd1 vssd1 vccd1 vccd1 _14761_/A sky130_fd_sc_hd__inv_2
X_11972_ _19376_/Q _11969_/X _09075_/X _11970_/X vssd1 vssd1 vccd1 vccd1 _19376_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17748__A1 _11093_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13711_ _13500_/Y _13710_/Y _13707_/Y vssd1 vssd1 vccd1 vccd1 _18760_/D sky130_fd_sc_hd__a21oi_1
XFILLER_244_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10923_ _10923_/A vssd1 vssd1 vccd1 vccd1 _10923_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_16_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14691_ _14780_/A vssd1 vssd1 vccd1 vccd1 _14691_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__17843__S1 _19632_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_232_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16430_ _18089_/Q vssd1 vssd1 vccd1 vccd1 _16430_/Y sky130_fd_sc_hd__inv_2
X_13642_ _17614_/X _13642_/B _15233_/B _13642_/D vssd1 vssd1 vccd1 vccd1 _13646_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_232_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10854_ _15823_/A _14245_/D vssd1 vssd1 vccd1 vccd1 _10856_/A sky130_fd_sc_hd__or2_2
XANTENNA__13234__B2 _17584_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14431__B1 _14417_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12187__B _12187_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16361_ _18104_/Q vssd1 vssd1 vccd1 vccd1 _16361_/Y sky130_fd_sc_hd__inv_2
X_13573_ _13573_/A vssd1 vssd1 vccd1 vccd1 _13573_/Y sky130_fd_sc_hd__inv_2
XFILLER_169_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10785_ _18653_/Q vssd1 vssd1 vccd1 vccd1 _10793_/B sky130_fd_sc_hd__buf_1
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18100_ _18260_/CLK _18100_/D vssd1 vssd1 vccd1 vccd1 _18100_/Q sky130_fd_sc_hd__dfxtp_1
X_15312_ _18625_/Q vssd1 vssd1 vccd1 vccd1 _15312_/Y sky130_fd_sc_hd__inv_2
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19080_ _19115_/CLK _19080_/D hold353/X vssd1 vssd1 vccd1 vccd1 _19080_/Q sky130_fd_sc_hd__dfrtp_1
X_12524_ _19070_/Q _12519_/X hold267/X _12520_/X vssd1 vssd1 vccd1 vccd1 _19070_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16292_ _18802_/Q _16043_/Y _18801_/Q _15957_/Y _16291_/X vssd1 vssd1 vccd1 vccd1
+ _16292_/X sky130_fd_sc_hd__o221a_1
XFILLER_9_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18031_ _18145_/CLK _18031_/D vssd1 vssd1 vccd1 vccd1 _18031_/Q sky130_fd_sc_hd__dfxtp_1
X_15243_ _18632_/Q vssd1 vssd1 vccd1 vccd1 _15243_/Y sky130_fd_sc_hd__inv_2
XFILLER_200_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12455_ _19116_/Q _12450_/X _12396_/X _12451_/X vssd1 vssd1 vccd1 vccd1 _19116_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_repeater148_A _17486_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11406_ _19546_/Q vssd1 vssd1 vccd1 vccd1 _11549_/A sky130_fd_sc_hd__inv_2
XFILLER_153_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15174_ _17943_/Q _15170_/X hold236/X _15172_/X vssd1 vssd1 vccd1 vccd1 _17943_/D
+ sky130_fd_sc_hd__a22o_1
X_12386_ hold286/X vssd1 vssd1 vccd1 vccd1 _12386_/X sky130_fd_sc_hd__buf_2
XFILLER_126_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14125_ _14018_/A _14018_/B _14123_/Y _14118_/X vssd1 vssd1 vccd1 vccd1 _18688_/D
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__16487__B2 _16506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11337_ _18963_/Q vssd1 vssd1 vccd1 vccd1 _11337_/Y sky130_fd_sc_hd__inv_2
X_19982_ _19992_/CLK _19982_/D repeater192/X vssd1 vssd1 vccd1 vccd1 _19982_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_98_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18933_ _19315_/CLK _18933_/D repeater215/X vssd1 vssd1 vccd1 vccd1 _18933_/Q sky130_fd_sc_hd__dfrtp_1
X_14056_ _19063_/Q _14005_/A _14053_/Y _18674_/Q _14055_/X vssd1 vssd1 vccd1 vccd1
+ _14064_/B sky130_fd_sc_hd__a221o_1
XFILLER_140_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11268_ _19589_/Q vssd1 vssd1 vccd1 vccd1 _11469_/A sky130_fd_sc_hd__inv_2
XFILLER_122_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13007_ _13007_/A _13011_/A vssd1 vssd1 vccd1 vccd1 _13008_/B sky130_fd_sc_hd__or2_2
X_10219_ _19838_/Q vssd1 vssd1 vccd1 vccd1 _10219_/Y sky130_fd_sc_hd__inv_2
X_18864_ _18866_/CLK _18864_/D repeater231/X vssd1 vssd1 vccd1 vccd1 _18864_/Q sky130_fd_sc_hd__dfrtp_4
X_11199_ _19592_/Q vssd1 vssd1 vccd1 vccd1 _11472_/A sky130_fd_sc_hd__inv_2
XFILLER_79_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10451__A _10451_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09017__A _09084_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17815_ _18333_/Q _18213_/Q _18205_/Q _18197_/Q _17918_/S0 _18750_/Q vssd1 vssd1
+ vccd1 vccd1 _17815_/X sky130_fd_sc_hd__mux4_1
X_18795_ _18795_/CLK _18795_/D repeater261/X vssd1 vssd1 vccd1 vccd1 _18795_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_95_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17746_ _17756_/S _11153_/Y _17753_/S vssd1 vssd1 vccd1 vccd1 _17746_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14958_ _18078_/Q _14952_/X _14929_/X _14954_/X vssd1 vssd1 vccd1 vccd1 _18078_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_223_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13909_ _13909_/A _13909_/B _13909_/C _13909_/D vssd1 vssd1 vccd1 vccd1 _13911_/C
+ sky130_fd_sc_hd__or4_4
X_17677_ _15527_/X _19458_/Q _17683_/S vssd1 vssd1 vccd1 vccd1 _18575_/D sky130_fd_sc_hd__mux2_1
XFILLER_35_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14889_ _18118_/Q _14883_/X _14810_/X _14885_/X vssd1 vssd1 vccd1 vccd1 _18118_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12378__A _12402_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17834__S1 _18752_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11282__A _19003_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16628_ _16959_/X _16597_/X _17074_/X _16598_/X vssd1 vssd1 vccd1 vccd1 _16629_/D
+ sky130_fd_sc_hd__a22o_2
X_19416_ _19905_/CLK _19416_/D repeater210/X vssd1 vssd1 vccd1 vccd1 _19416_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_51_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14422__B1 _14405_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19839__RESET_B repeater270/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16559_ _16504_/X _16552_/X _16554_/X _16558_/Y vssd1 vssd1 vccd1 vccd1 _16559_/Y
+ sky130_fd_sc_hd__o211ai_4
X_19347_ _19952_/CLK _19347_/D repeater245/X vssd1 vssd1 vccd1 vccd1 _19347_/Q sky130_fd_sc_hd__dfrtp_4
X_09100_ hold264/X vssd1 vssd1 vccd1 vccd1 _10423_/A sky130_fd_sc_hd__clkbuf_2
X_19278_ _19315_/CLK _19278_/D repeater215/X vssd1 vssd1 vccd1 vccd1 _19278_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_31_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_176_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09031_ _09043_/A vssd1 vssd1 vccd1 vccd1 _09031_/X sky130_fd_sc_hd__buf_1
XFILLER_176_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18229_ _18412_/CLK _18229_/D vssd1 vssd1 vccd1 vccd1 _18229_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold301 input50/X vssd1 vssd1 vccd1 vccd1 hold301/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold312 input72/X vssd1 vssd1 vccd1 vccd1 hold312/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 HWDATA[0] vssd1 vssd1 vccd1 vccd1 input38/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold334 hold334/A vssd1 vssd1 vccd1 vccd1 hold334/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold345 hold345/A vssd1 vssd1 vccd1 vccd1 hold361/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold356 hold356/A vssd1 vssd1 vccd1 vccd1 hold356/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17770__S0 _17923_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold367 hold367/A vssd1 vssd1 vccd1 vccd1 hold367/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20122_ _20122_/CLK _20122_/D repeater234/X vssd1 vssd1 vccd1 vccd1 _20122_/Q sky130_fd_sc_hd__dfrtp_1
X_09933_ _19943_/Q _16215_/A _09851_/A _19334_/Q _09932_/X vssd1 vssd1 vccd1 vccd1
+ _09947_/A sky130_fd_sc_hd__o221a_1
XANTENNA__15150__B2 _15148_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20053_ _20055_/CLK _20053_/D repeater205/X vssd1 vssd1 vccd1 vccd1 _20053_/Q sky130_fd_sc_hd__dfrtp_1
X_09864_ _09864_/A _09975_/A vssd1 vssd1 vccd1 vccd1 _09865_/B sky130_fd_sc_hd__or2_2
XFILLER_86_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15871__B _15878_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09795_ _19983_/Q _09794_/Y _09731_/A _09740_/B vssd1 vssd1 vccd1 vccd1 _19983_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_246_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater151 _17459_/S vssd1 vssd1 vccd1 vccd1 _17487_/S sky130_fd_sc_hd__buf_8
Xrepeater162 _17473_/S vssd1 vssd1 vccd1 vccd1 _17547_/S sky130_fd_sc_hd__buf_8
XANTENNA__14110__C1 _14135_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater173 _17524_/S vssd1 vssd1 vccd1 vccd1 _17488_/S sky130_fd_sc_hd__buf_8
XPHY_4305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14661__B1 _14606_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater184 _18749_/Q vssd1 vssd1 vccd1 vccd1 _17918_/S0 sky130_fd_sc_hd__clkbuf_16
Xrepeater195 repeater199/X vssd1 vssd1 vccd1 vccd1 repeater195/X sky130_fd_sc_hd__buf_8
XPHY_4327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17825__S1 _18750_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_214_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11192__A _11192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_214_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold143_A HADDR[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10570_ _10613_/A _10615_/A vssd1 vssd1 vccd1 vccd1 _10938_/B sky130_fd_sc_hd__nor2_1
XFILLER_210_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09229_ _19882_/Q vssd1 vssd1 vccd1 vccd1 _09229_/Y sky130_fd_sc_hd__inv_2
XFILLER_158_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16922__S _17534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19162__RESET_B hold370/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12240_ hold322/X vssd1 vssd1 vccd1 vccd1 _14405_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_108_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10255__B _10410_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12171_ _12171_/A vssd1 vssd1 vccd1 vccd1 _12171_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_150_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20067__RESET_B repeater207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11122_ _17747_/X vssd1 vssd1 vccd1 vccd1 _11123_/A sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_112_HCLK_A clkbuf_opt_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17418__A0 _17486_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11053_ _11056_/A _11053_/B vssd1 vssd1 vccd1 vccd1 _11053_/X sky130_fd_sc_hd__or2_1
X_15930_ _18347_/Q vssd1 vssd1 vccd1 vccd1 _15930_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10004_ _19363_/Q vssd1 vssd1 vccd1 vccd1 _10004_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15861_ _19126_/Q vssd1 vssd1 vccd1 vccd1 _15861_/Y sky130_fd_sc_hd__inv_2
XFILLER_190_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17600_ _18490_/Q _15335_/Y _17600_/S vssd1 vssd1 vccd1 vccd1 _17600_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14812_ _14812_/A vssd1 vssd1 vccd1 vccd1 _14812_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_190_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18580_ _19561_/CLK _18580_/D hold348/A vssd1 vssd1 vccd1 vccd1 _18580_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_17_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15792_ _18146_/Q vssd1 vssd1 vccd1 vccd1 _15792_/Y sky130_fd_sc_hd__inv_2
XFILLER_123_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17531_ _15871_/Y _13483_/A _17537_/S vssd1 vssd1 vccd1 vccd1 _17531_/X sky130_fd_sc_hd__mux2_1
X_14743_ _14743_/A _18755_/Q _14975_/C vssd1 vssd1 vccd1 vccd1 _14746_/A sky130_fd_sc_hd__or3_4
X_11955_ _11955_/A vssd1 vssd1 vccd1 vccd1 _11955_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__17816__S1 _18750_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10906_ _18637_/Q vssd1 vssd1 vccd1 vccd1 _10907_/B sky130_fd_sc_hd__inv_2
XFILLER_33_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17462_ _16045_/X _19880_/Q _19498_/Q vssd1 vssd1 vccd1 vccd1 _17462_/X sky130_fd_sc_hd__mux2_1
XFILLER_178_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14674_ _18239_/Q _14669_/X _09174_/X _14671_/X vssd1 vssd1 vccd1 vccd1 _18239_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_232_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14404__B1 _14403_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11886_ _19427_/Q _11884_/X _09030_/X _11885_/X vssd1 vssd1 vccd1 vccd1 _19427_/D
+ sky130_fd_sc_hd__a22o_1
X_19201_ _19585_/CLK _19201_/D hold365/X vssd1 vssd1 vccd1 vccd1 _19201_/Q sky130_fd_sc_hd__dfrtp_4
X_16413_ _18049_/Q vssd1 vssd1 vccd1 vccd1 _16413_/Y sky130_fd_sc_hd__inv_2
X_13625_ _13622_/X _13621_/X _13622_/X _13621_/X vssd1 vssd1 vccd1 vccd1 _18802_/D
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_220_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10837_ _19718_/Q vssd1 vssd1 vccd1 vccd1 _15735_/A sky130_fd_sc_hd__inv_2
XFILLER_158_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17393_ _16206_/Y _09320_/Y _19498_/Q vssd1 vssd1 vccd1 vccd1 _17393_/X sky130_fd_sc_hd__mux2_1
XANTENNA_repeater265_A repeater267/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19132_ _19970_/CLK _19132_/D repeater249/X vssd1 vssd1 vccd1 vccd1 _19132_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_186_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16344_ _18248_/Q _16344_/B vssd1 vssd1 vccd1 vccd1 _16344_/X sky130_fd_sc_hd__and2_1
X_13556_ _13556_/A _13563_/A vssd1 vssd1 vccd1 vccd1 _13557_/B sky130_fd_sc_hd__or2_2
X_10768_ _10764_/Y _10767_/Y _10286_/A _10762_/X vssd1 vssd1 vccd1 vccd1 _19752_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_118_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12507_ _19082_/Q _12505_/X _12401_/X _12506_/X vssd1 vssd1 vccd1 vccd1 _19082_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_8_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19063_ _19585_/CLK _19063_/D hold361/X vssd1 vssd1 vccd1 vccd1 _19063_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_118_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16275_ _18127_/Q vssd1 vssd1 vccd1 vccd1 _16275_/Y sky130_fd_sc_hd__inv_2
X_13487_ _13322_/B _13486_/A _18839_/Q _13489_/A _13421_/X vssd1 vssd1 vccd1 vccd1
+ _18839_/D sky130_fd_sc_hd__o221a_1
XANTENNA__16832__S _17534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10446__A _10446_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10699_ _10698_/X _17749_/X _17749_/S _10694_/Y _19777_/Q vssd1 vssd1 vccd1 vccd1
+ _19777_/D sky130_fd_sc_hd__a32o_1
XFILLER_185_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_218_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18014_ _18169_/CLK _18014_/D vssd1 vssd1 vccd1 vccd1 _18014_/Q sky130_fd_sc_hd__dfxtp_1
X_15226_ _19721_/Q vssd1 vssd1 vccd1 vccd1 _15226_/Y sky130_fd_sc_hd__inv_2
XFILLER_172_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12438_ _12313_/X _19125_/Q _12438_/S vssd1 vssd1 vccd1 vccd1 _19125_/D sky130_fd_sc_hd__mux2_1
XFILLER_160_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15157_ _18765_/Q _18764_/Q _15157_/C vssd1 vssd1 vccd1 vccd1 _15159_/A sky130_fd_sc_hd__or3_4
X_12369_ _19158_/Q _12334_/A _12241_/X _12335_/A vssd1 vssd1 vccd1 vccd1 _19158_/D
+ sky130_fd_sc_hd__a22o_1
X_14108_ _14108_/A vssd1 vssd1 vccd1 vccd1 _14108_/Y sky130_fd_sc_hd__clkinv_1
XFILLER_114_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15088_ _17999_/Q _15083_/X hold244/X _15085_/X vssd1 vssd1 vccd1 vccd1 _17999_/D
+ sky130_fd_sc_hd__a22o_1
X_19965_ _19965_/CLK _19965_/D repeater185/X vssd1 vssd1 vccd1 vccd1 _19965_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_102_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17409__A0 _17486_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16880__A1 _09426_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18814__RESET_B repeater239/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14039_ _19080_/Q vssd1 vssd1 vccd1 vccd1 _14039_/Y sky130_fd_sc_hd__inv_2
X_18916_ _19222_/CLK _18916_/D repeater186/X vssd1 vssd1 vccd1 vccd1 _18916_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_67_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19896_ _20064_/CLK _19896_/D repeater198/X vssd1 vssd1 vccd1 vccd1 _19896_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_110_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18847_ _18866_/CLK _18847_/D repeater232/X vssd1 vssd1 vccd1 vccd1 _18847_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_34_HCLK_A _18641_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13492__A _15858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_97_HCLK_A clkbuf_4_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_243_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09580_ _09580_/A vssd1 vssd1 vccd1 vccd1 _09580_/Y sky130_fd_sc_hd__inv_2
X_18778_ _19855_/CLK _18778_/D repeater264/X vssd1 vssd1 vccd1 vccd1 _18778_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_208_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_236_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17729_ _15380_/X _19716_/Q _18508_/D vssd1 vssd1 vccd1 vccd1 _17729_/X sky130_fd_sc_hd__mux2_1
XFILLER_208_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17807__S1 _18750_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_224_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19780__CLK _19780_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09014_ _09084_/A vssd1 vssd1 vccd1 vccd1 _09041_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_117_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold131 HADDR[21] vssd1 vssd1 vccd1 vccd1 input14/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold142 input13/X vssd1 vssd1 vccd1 vccd1 hold142/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold153 input9/X vssd1 vssd1 vccd1 vccd1 hold153/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11932__A1 _15512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold164 hold164/A vssd1 vssd1 vccd1 vccd1 hold164/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 HADDR[12] vssd1 vssd1 vccd1 vccd1 input4/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold186 input30/X vssd1 vssd1 vccd1 vccd1 hold186/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold197 HADDR[4] vssd1 vssd1 vccd1 vccd1 input27/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17573__S _17584_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20105_ _20107_/CLK _20105_/D repeater230/X vssd1 vssd1 vccd1 vccd1 _20105_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_160_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09916_ _19960_/Q _09912_/Y _19956_/Q _16588_/A _09915_/X vssd1 vssd1 vccd1 vccd1
+ _09928_/A sky130_fd_sc_hd__o221a_1
XFILLER_247_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20036_ _20036_/CLK _20036_/D repeater198/X vssd1 vssd1 vccd1 vccd1 _20036_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__11696__B1 _10861_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09847_ _19939_/Q vssd1 vssd1 vccd1 vccd1 _09848_/A sky130_fd_sc_hd__inv_2
XFILLER_219_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09778_ _09778_/A vssd1 vssd1 vccd1 vccd1 _09778_/Y sky130_fd_sc_hd__inv_2
XFILLER_246_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_233_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_233_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16917__S _17534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11740_ _15749_/C _11737_/X _16931_/X _11738_/X vssd1 vssd1 vccd1 vccd1 _19499_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16387__B1 _15333_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11671_ _11674_/A vssd1 vssd1 vccd1 vccd1 _11671_/X sky130_fd_sc_hd__clkbuf_2
XPHY_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13410_ _20112_/Q vssd1 vssd1 vccd1 vccd1 _13410_/Y sky130_fd_sc_hd__inv_2
XFILLER_168_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19343__RESET_B repeater244/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10622_ _10939_/B _10618_/X _10574_/X _10608_/A vssd1 vssd1 vccd1 vccd1 _19809_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_186_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14390_ _18402_/Q _14381_/A _14268_/X _14382_/A vssd1 vssd1 vccd1 vccd1 _18402_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13341_ _13429_/B _13453_/A vssd1 vssd1 vccd1 vccd1 _13342_/B sky130_fd_sc_hd__or2_2
XFILLER_128_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10553_ _10553_/A vssd1 vssd1 vccd1 vccd1 _10616_/C sky130_fd_sc_hd__inv_2
XFILLER_139_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_194_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16060_ _19758_/Q vssd1 vssd1 vccd1 vccd1 _16060_/Y sky130_fd_sc_hd__inv_2
XFILLER_154_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19503__CLK _19510_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13272_ _14366_/B _13271_/Y _14366_/B _13271_/Y vssd1 vssd1 vccd1 vccd1 _13278_/C
+ sky130_fd_sc_hd__a2bb2o_1
X_10484_ _19540_/Q vssd1 vssd1 vccd1 vccd1 _10491_/B sky130_fd_sc_hd__inv_2
XFILLER_182_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15011_ _15011_/A vssd1 vssd1 vccd1 vccd1 _15012_/A sky130_fd_sc_hd__inv_2
X_12223_ hold268/X vssd1 vssd1 vccd1 vccd1 _12223_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__10187__A0 _09339_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12154_ _19281_/Q _12150_/X _12100_/X _12151_/X vssd1 vssd1 vccd1 vccd1 _19281_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17483__S _17534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11105_ _19636_/Q vssd1 vssd1 vccd1 vccd1 _11105_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19750_ _19900_/CLK _19750_/D repeater197/X vssd1 vssd1 vccd1 vccd1 _19750_/Q sky130_fd_sc_hd__dfrtp_1
X_16962_ _16961_/X _13552_/A _17536_/S vssd1 vssd1 vccd1 vccd1 _16962_/X sky130_fd_sc_hd__mux2_1
X_12085_ _19320_/Q _12082_/X _12083_/X _12084_/X vssd1 vssd1 vccd1 vccd1 _19320_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_111_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18701_ _18701_/CLK _18701_/D hold351/X vssd1 vssd1 vccd1 vccd1 _18701_/Q sky130_fd_sc_hd__dfrtp_2
X_11036_ _19650_/Q _11022_/X _11029_/B _11035_/X vssd1 vssd1 vccd1 vccd1 _19650_/D
+ sky130_fd_sc_hd__a31o_1
X_15913_ _17554_/X vssd1 vssd1 vccd1 vccd1 _15913_/Y sky130_fd_sc_hd__inv_2
X_19681_ _19795_/CLK _19681_/D repeater219/X vssd1 vssd1 vccd1 vccd1 _19681_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_76_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16893_ _16892_/X _12938_/Y _17487_/S vssd1 vssd1 vccd1 vccd1 _16893_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18632_ _18633_/CLK _18632_/D repeater225/X vssd1 vssd1 vccd1 vccd1 _18632_/Q sky130_fd_sc_hd__dfrtp_1
X_15844_ _15834_/Y _15836_/X _15837_/Y _15838_/X _15843_/X vssd1 vssd1 vccd1 vccd1
+ _15844_/X sky130_fd_sc_hd__o221a_1
XFILLER_225_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18563_ _20058_/CLK _18563_/D repeater194/X vssd1 vssd1 vccd1 vccd1 _18563_/Q sky130_fd_sc_hd__dfrtp_1
X_15775_ _19192_/Q _18736_/Q vssd1 vssd1 vccd1 vccd1 _15775_/X sky130_fd_sc_hd__and2_1
X_12987_ _12964_/B _12881_/B _12983_/Y _12986_/X vssd1 vssd1 vccd1 vccd1 _18939_/D
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__16827__S _17524_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_233_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14726_ _18213_/Q _14717_/X _14725_/X _14719_/X vssd1 vssd1 vccd1 vccd1 _18213_/D
+ sky130_fd_sc_hd__a22o_1
X_17514_ _15878_/Y _15479_/A _17537_/S vssd1 vssd1 vccd1 vccd1 _17514_/X sky130_fd_sc_hd__mux2_1
XFILLER_206_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11938_ _11977_/A vssd1 vssd1 vccd1 vccd1 _11955_/A sky130_fd_sc_hd__clkbuf_2
X_18494_ _20089_/CLK _18494_/D repeater203/X vssd1 vssd1 vccd1 vccd1 _18494_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_33_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_220_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17445_ _17444_/X _09850_/A _17518_/S vssd1 vssd1 vccd1 vccd1 _17445_/X sky130_fd_sc_hd__mux2_1
X_14657_ _14657_/A vssd1 vssd1 vccd1 vccd1 _14658_/A sky130_fd_sc_hd__inv_2
XFILLER_220_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11869_ _11869_/A _11869_/B vssd1 vssd1 vccd1 vccd1 _11869_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__15050__B1 _14992_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19084__RESET_B hold351/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13608_ _18807_/Q _13607_/Y _13591_/X _13608_/C1 vssd1 vssd1 vccd1 vccd1 _18807_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_32_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17376_ _17375_/X _16271_/Y _17567_/S vssd1 vssd1 vccd1 vccd1 _17376_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14588_ _14588_/A vssd1 vssd1 vccd1 vccd1 _14589_/A sky130_fd_sc_hd__inv_2
XANTENNA__20010__CLK _20091_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09030__A hold303/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19115_ _19115_/CLK _19115_/D hold353/X vssd1 vssd1 vccd1 vccd1 _19115_/Q sky130_fd_sc_hd__dfrtp_1
X_16327_ _15846_/A _16310_/X _15859_/A _16319_/X _16326_/X vssd1 vssd1 vccd1 vccd1
+ _16327_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_201_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13539_ _13539_/A _13539_/B vssd1 vssd1 vccd1 vccd1 _13590_/A sky130_fd_sc_hd__or2_1
XANTENNA__11611__B1 _11617_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19046_ _19566_/CLK _19046_/D repeater255/X vssd1 vssd1 vccd1 vccd1 _19046_/Q sky130_fd_sc_hd__dfrtp_1
X_16258_ _18039_/Q vssd1 vssd1 vccd1 vccd1 _16258_/Y sky130_fd_sc_hd__inv_2
X_15209_ _15205_/Y _18635_/Q _15206_/Y _15208_/Y vssd1 vssd1 vccd1 vccd1 _15209_/X
+ sky130_fd_sc_hd__a31o_1
X_16189_ _15218_/Y _15388_/A _15216_/C _15213_/X vssd1 vssd1 vccd1 vccd1 _16189_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_161_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10178__B1 _09101_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13116__B1 _19169_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17393__S _19498_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19948_ _19976_/CLK _19948_/D hold371/X vssd1 vssd1 vccd1 vccd1 _19948_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_229_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09701_ _19996_/Q _19425_/Q _19996_/Q _19425_/Q vssd1 vssd1 vccd1 vccd1 _09701_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_19879_ _20059_/CLK _19879_/D repeater199/X vssd1 vssd1 vccd1 vccd1 _19879_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_110_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16605__B2 _15887_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09632_ _19975_/Q vssd1 vssd1 vccd1 vccd1 _09635_/A sky130_fd_sc_hd__inv_2
XFILLER_55_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09563_ _09466_/A _19295_/Q _20020_/Q _09559_/Y _09562_/X vssd1 vssd1 vccd1 vccd1
+ _09564_/D sky130_fd_sc_hd__o221a_1
XFILLER_82_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09494_ _09494_/A _09494_/B vssd1 vssd1 vccd1 vccd1 _09495_/A sky130_fd_sc_hd__or2_1
XPHY_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15041__B1 _15000_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_91_HCLK clkbuf_4_12_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19984_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_183_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17568__S _17568_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18736__RESET_B repeater244/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10169__B1 _09077_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16501__A _20101_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20019_ _20120_/CLK _20019_/D repeater238/X vssd1 vssd1 vccd1 vccd1 _20019_/Q sky130_fd_sc_hd__dfrtp_1
X_12910_ _19286_/Q _18943_/Q _12909_/Y _12885_/A vssd1 vssd1 vccd1 vccd1 _12916_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_207_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13890_ _13886_/Y _18729_/Q _19211_/Q _13910_/A _13889_/X vssd1 vssd1 vccd1 vccd1
+ _13897_/B sky130_fd_sc_hd__o221a_1
XFILLER_234_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14607__B1 _14606_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_80_HCLK_A clkbuf_4_13_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12841_ _18943_/Q vssd1 vssd1 vccd1 vccd1 _12885_/A sky130_fd_sc_hd__inv_4
XFILLER_73_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15560_ _15559_/Y _15556_/A _18583_/Q _15556_/Y _15512_/A vssd1 vssd1 vccd1 vccd1
+ _15560_/X sky130_fd_sc_hd__o221a_1
X_12772_ _19246_/Q vssd1 vssd1 vccd1 vccd1 _12772_/Y sky130_fd_sc_hd__inv_2
XPHY_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_242_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14511_ hold331/X vssd1 vssd1 vccd1 vccd1 hold330/A sky130_fd_sc_hd__clkbuf_2
XFILLER_70_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ _11730_/A vssd1 vssd1 vccd1 vccd1 _11723_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_202_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15491_ _15491_/A _15491_/B vssd1 vssd1 vccd1 vccd1 _15491_/Y sky130_fd_sc_hd__nor2_1
XFILLER_9_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15032__B1 _15006_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17230_ _16484_/X _08947_/Y _17566_/S vssd1 vssd1 vccd1 vccd1 _17230_/X sky130_fd_sc_hd__mux2_1
XPHY_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14442_ _18376_/Q _14436_/X _14441_/X _14439_/X vssd1 vssd1 vccd1 vccd1 _18376_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_42_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11654_ _11654_/A _11654_/B vssd1 vssd1 vccd1 vccd1 _11655_/B sky130_fd_sc_hd__or2_1
XFILLER_187_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10605_ _10617_/A vssd1 vssd1 vccd1 vccd1 _10606_/A sky130_fd_sc_hd__buf_1
XFILLER_196_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17161_ _17160_/X _09476_/A _17482_/S vssd1 vssd1 vccd1 vccd1 _17161_/X sky130_fd_sc_hd__mux2_2
XANTENNA__17478__S _17523_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14373_ _18414_/Q _14367_/X hold324/X _14369_/X vssd1 vssd1 vccd1 vccd1 _18414_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20082__RESET_B repeater204/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11585_ _11585_/A _11594_/A vssd1 vssd1 vccd1 vccd1 _11586_/A sky130_fd_sc_hd__or2_2
XANTENNA__14691__A _14780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16112_ _18109_/Q vssd1 vssd1 vccd1 vccd1 _16112_/Y sky130_fd_sc_hd__inv_2
X_13324_ _18843_/Q vssd1 vssd1 vccd1 vccd1 _13466_/A sky130_fd_sc_hd__inv_2
X_10536_ _11648_/A vssd1 vssd1 vccd1 vccd1 _15443_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_183_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17092_ _17091_/X _13067_/A _17488_/S vssd1 vssd1 vccd1 vccd1 _17092_/X sky130_fd_sc_hd__mux2_1
XFILLER_116_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16043_ _17963_/Q vssd1 vssd1 vccd1 vccd1 _16043_/Y sky130_fd_sc_hd__inv_2
X_13255_ _18752_/Q vssd1 vssd1 vccd1 vccd1 _13255_/Y sky130_fd_sc_hd__inv_2
X_10467_ _19824_/Q _10466_/X _18548_/Q _10462_/Y vssd1 vssd1 vccd1 vccd1 _19824_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_89_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12206_ _12206_/A vssd1 vssd1 vccd1 vccd1 _12206_/X sky130_fd_sc_hd__clkbuf_2
X_13186_ _13077_/A _13186_/A2 _13184_/Y _13182_/X vssd1 vssd1 vccd1 vccd1 _18905_/D
+ sky130_fd_sc_hd__a211oi_4
X_10398_ _19850_/Q vssd1 vssd1 vccd1 vccd1 _11096_/A sky130_fd_sc_hd__inv_2
XFILLER_69_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19802_ _19808_/CLK _19802_/D repeater224/X vssd1 vssd1 vccd1 vccd1 _19802_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_97_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12137_ _12151_/A vssd1 vssd1 vccd1 vccd1 _12137_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_124_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17994_ _18412_/CLK _17994_/D vssd1 vssd1 vccd1 vccd1 _17994_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19733_ _20051_/CLK _19733_/D repeater208/X vssd1 vssd1 vccd1 vccd1 _19733_/Q sky130_fd_sc_hd__dfrtp_1
X_12068_ _12094_/A vssd1 vssd1 vccd1 vccd1 _12068_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_1_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16945_ _19489_/Q hold133/X _16946_/S vssd1 vssd1 vccd1 vccd1 _16945_/X sky130_fd_sc_hd__mux2_1
XFILLER_237_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11019_ _19654_/Q _19653_/Q _10224_/X _10211_/X vssd1 vssd1 vccd1 vccd1 _11019_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_65_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19664_ _19667_/CLK _19664_/D repeater264/X vssd1 vssd1 vccd1 vccd1 _19664_/Q sky130_fd_sc_hd__dfrtp_1
X_16876_ _15963_/X _09500_/Y _17534_/S vssd1 vssd1 vccd1 vccd1 _16876_/X sky130_fd_sc_hd__mux2_1
XFILLER_64_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16599__B1 _17245_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_231_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17260__A1 _19143_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_237_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18615_ _19157_/CLK _18615_/D repeater267/X vssd1 vssd1 vccd1 vccd1 _18615_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__09025__A hold279/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15827_ _15866_/A vssd1 vssd1 vccd1 vccd1 _15828_/A sky130_fd_sc_hd__clkbuf_2
X_19595_ _19595_/CLK _19595_/D repeater282/X vssd1 vssd1 vccd1 vccd1 _19595_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__19265__RESET_B repeater245/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15758_ _18886_/Q _18884_/Q vssd1 vssd1 vccd1 vccd1 _15758_/X sky130_fd_sc_hd__or2_1
X_18546_ _19920_/CLK _18546_/D repeater220/X vssd1 vssd1 vccd1 vccd1 _18546_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__12085__B1 _12083_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17012__A1 _09918_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10096__C1 _10107_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14709_ _14709_/A vssd1 vssd1 vccd1 vccd1 _14709_/X sky130_fd_sc_hd__clkbuf_2
X_18477_ _19780_/CLK _18477_/D repeater227/X vssd1 vssd1 vccd1 vccd1 _18477_/Q sky130_fd_sc_hd__dfrtp_1
X_15689_ _15687_/Y _15688_/Y _15673_/X vssd1 vssd1 vccd1 vccd1 _15689_/X sky130_fd_sc_hd__o21a_1
XANTENNA__12386__A hold286/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14377__A2 _14368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17428_ _16117_/X _19881_/Q _19498_/Q vssd1 vssd1 vccd1 vccd1 _17428_/X sky130_fd_sc_hd__mux2_1
XFILLER_178_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17388__S _17488_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19699__CLK _20051_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17359_ _17358_/X _13533_/A _17386_/S vssd1 vssd1 vccd1 vccd1 _17359_/X sky130_fd_sc_hd__mux2_4
XFILLER_118_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19029_ _19667_/CLK _19029_/D repeater264/X vssd1 vssd1 vccd1 vccd1 _19029_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_134_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08994_ _18620_/Q vssd1 vssd1 vccd1 vccd1 _10250_/C sky130_fd_sc_hd__inv_2
XFILLER_248_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14837__B1 _14808_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_229_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16678__D _16678_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_229_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17251__A1 _19383_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09615_ _09615_/A vssd1 vssd1 vccd1 vccd1 _09615_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09546_ _19298_/Q vssd1 vssd1 vccd1 vccd1 _16212_/A sky130_fd_sc_hd__inv_2
XFILLER_24_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_221_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11823__B1 _10882_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09477_ _09477_/A _09598_/A vssd1 vssd1 vccd1 vccd1 _09478_/B sky130_fd_sc_hd__or2_1
XPHY_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12296__A _14273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15014__B1 _14996_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17298__S _17524_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11370_ _11620_/A _19130_/Q _11576_/A _19143_/Q vssd1 vssd1 vccd1 vccd1 _11370_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_50_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16514__B1 _17282_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16215__B _16469_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10321_ _10321_/A _10321_/B _10321_/C _10321_/D vssd1 vssd1 vccd1 vccd1 _10375_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_166_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16930__S _16950_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13040_ _18906_/Q vssd1 vssd1 vccd1 vccd1 _13078_/A sky130_fd_sc_hd__inv_2
X_10252_ _11936_/A _15899_/A vssd1 vssd1 vccd1 vccd1 _10409_/A sky130_fd_sc_hd__or2_2
XFILLER_105_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10183_ _15715_/B _10759_/C vssd1 vssd1 vccd1 vccd1 _10290_/B sky130_fd_sc_hd__and2_1
XFILLER_132_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14828__B1 hold263/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14991_ _14993_/A vssd1 vssd1 vccd1 vccd1 _14991_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_219_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16730_ _19055_/Q vssd1 vssd1 vccd1 vccd1 _16730_/Y sky130_fd_sc_hd__inv_2
X_13942_ _18717_/Q _13941_/Y _13925_/A _13817_/B vssd1 vssd1 vccd1 vccd1 _18717_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_87_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_247_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16661_ _16995_/X _16573_/X _17024_/X _16574_/X _16660_/X vssd1 vssd1 vccd1 vccd1
+ _16664_/B sky130_fd_sc_hd__o221a_4
X_13873_ _13872_/Y _18710_/Q _13838_/Y _13873_/B2 vssd1 vssd1 vccd1 vccd1 _13873_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_35_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15612_ _15612_/A vssd1 vssd1 vccd1 vccd1 _15618_/B sky130_fd_sc_hd__inv_2
X_18400_ _18416_/CLK _18400_/D vssd1 vssd1 vccd1 vccd1 _18400_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12824_ _18829_/Q vssd1 vssd1 vccd1 vccd1 _13552_/A sky130_fd_sc_hd__inv_2
X_19380_ _19927_/CLK _19380_/D repeater230/X vssd1 vssd1 vccd1 vccd1 _19380_/Q sky130_fd_sc_hd__dfrtp_2
X_16592_ _17248_/X _16563_/X _17237_/X _16591_/X vssd1 vssd1 vccd1 vccd1 _16600_/A
+ sky130_fd_sc_hd__o22ai_2
XFILLER_131_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_243_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15543_ _18579_/Q _15538_/Y _15541_/Y _15538_/A _15542_/X vssd1 vssd1 vccd1 vccd1
+ _15543_/X sky130_fd_sc_hd__o221a_1
X_18331_ _18412_/CLK _18331_/D vssd1 vssd1 vccd1 vccd1 _18331_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12755_ _18811_/Q vssd1 vssd1 vccd1 vccd1 _13535_/A sky130_fd_sc_hd__inv_2
XFILLER_187_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15005__B1 _15004_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_repeater178_A _17414_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11706_ _18622_/D hold213/X vssd1 vssd1 vccd1 vccd1 _11737_/A sky130_fd_sc_hd__or2b_1
X_18262_ _20077_/CLK _18262_/D vssd1 vssd1 vccd1 vccd1 _18262_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15474_ _15474_/A vssd1 vssd1 vccd1 vccd1 _15474_/Y sky130_fd_sc_hd__inv_2
XFILLER_203_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12686_ _18976_/Q _12684_/X hold277/X _12685_/X vssd1 vssd1 vccd1 vccd1 _18976_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13567__B1 _13560_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14425_ _14425_/A vssd1 vssd1 vccd1 vccd1 _14426_/A sky130_fd_sc_hd__inv_2
X_17213_ _17212_/X _09694_/Y _17523_/S vssd1 vssd1 vccd1 vccd1 _17213_/X sky130_fd_sc_hd__mux2_1
XPHY_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11637_ _11637_/A vssd1 vssd1 vccd1 vccd1 _11641_/A sky130_fd_sc_hd__inv_2
X_18193_ _18216_/CLK _18193_/D vssd1 vssd1 vccd1 vccd1 _18193_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18658__RESET_B repeater210/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17001__S _17490_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17144_ _15963_/X _09531_/Y _17534_/S vssd1 vssd1 vccd1 vccd1 _17144_/X sky130_fd_sc_hd__mux2_1
XPHY_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14356_ _14749_/A vssd1 vssd1 vccd1 vccd1 _14356_/X sky130_fd_sc_hd__clkbuf_2
XPHY_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11568_ _11561_/C _11590_/B _11561_/A vssd1 vssd1 vccd1 vccd1 _11569_/C sky130_fd_sc_hd__o21a_1
XANTENNA__19991__CLK _19992_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13307_ _18858_/Q vssd1 vssd1 vccd1 vccd1 _13428_/A sky130_fd_sc_hd__inv_2
X_10519_ _10530_/C _10530_/A _19543_/Q _10519_/D vssd1 vssd1 vccd1 vccd1 _11651_/B
+ sky130_fd_sc_hd__and4b_1
X_17075_ _16643_/Y _18982_/Q _17493_/S vssd1 vssd1 vccd1 vccd1 _17075_/X sky130_fd_sc_hd__mux2_1
X_14287_ _14366_/A _14758_/B _15082_/C vssd1 vssd1 vccd1 vccd1 _14289_/A sky130_fd_sc_hd__or3_4
XFILLER_128_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11499_ _11484_/A _11484_/B _11528_/A _11497_/Y vssd1 vssd1 vccd1 vccd1 _19604_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_226_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16026_ _18124_/Q vssd1 vssd1 vccd1 vccd1 _16026_/Y sky130_fd_sc_hd__inv_2
X_13238_ _18627_/Q _11647_/Y _18880_/Q _15389_/A vssd1 vssd1 vccd1 vccd1 _18880_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_170_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10002__C1 _09964_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13169_ _13169_/A vssd1 vssd1 vccd1 vccd1 _13169_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17977_ _18260_/CLK _17977_/D vssd1 vssd1 vccd1 vccd1 _17977_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17671__S _17683_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19716_ _19794_/CLK _19716_/D repeater201/X vssd1 vssd1 vccd1 vccd1 _19716_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_38_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16928_ _19472_/Q hold202/X _16946_/S vssd1 vssd1 vccd1 vccd1 _16928_/X sky130_fd_sc_hd__mux2_2
XFILLER_38_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19647_ _19647_/CLK _19647_/D repeater261/X vssd1 vssd1 vccd1 vccd1 _19647_/Q sky130_fd_sc_hd__dfrtp_2
X_16859_ _16858_/X _09483_/A _17482_/S vssd1 vssd1 vccd1 vccd1 _16859_/X sky130_fd_sc_hd__mux2_1
XFILLER_81_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09400_ _19930_/Q _19390_/Q _10046_/A _09399_/Y vssd1 vssd1 vccd1 vccd1 _09400_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_92_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19578_ _19600_/CLK _19578_/D hold355/X vssd1 vssd1 vccd1 vccd1 _19578_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_92_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13404__A1_N _20105_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09331_ _20045_/Q _15723_/A _09323_/X _09327_/X _09330_/X vssd1 vssd1 vccd1 vccd1
+ _09331_/X sky130_fd_sc_hd__o2111a_1
XFILLER_240_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18529_ _19937_/CLK _18529_/D repeater189/X vssd1 vssd1 vccd1 vccd1 _18529_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__11805__B1 _09049_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09262_ _19499_/Q vssd1 vssd1 vccd1 vccd1 _14245_/C sky130_fd_sc_hd__inv_2
XFILLER_194_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09193_ _20072_/Q _20071_/Q _08917_/A vssd1 vssd1 vccd1 vccd1 _09193_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__17919__S0 _18751_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12230__B1 _11978_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_121_HCLK clkbuf_opt_0_HCLK/A vssd1 vssd1 vccd1 vccd1 _19600_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_103_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17472__A1 _17894_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08977_ _09203_/A _09205_/A _08977_/C vssd1 vssd1 vccd1 vccd1 _09199_/A sky130_fd_sc_hd__or3_4
XANTENNA__17581__S _17584_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15890__A _15890_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12297__B1 _12296_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_229_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12836__A2 _13597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_232_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12049__B1 _11922_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10870_ _11926_/A vssd1 vssd1 vccd1 vccd1 _10870_/X sky130_fd_sc_hd__buf_2
XFILLER_232_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09529_ _19315_/Q vssd1 vssd1 vccd1 vccd1 _09529_/Y sky130_fd_sc_hd__inv_2
XPHY_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16925__S _16950_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_212_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12540_ hold336/X vssd1 vssd1 vccd1 vccd1 hold335/A sky130_fd_sc_hd__clkbuf_2
XFILLER_240_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_236_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12471_ _12478_/A vssd1 vssd1 vccd1 vccd1 _12471_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__18751__RESET_B repeater195/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14210_ _19097_/Q vssd1 vssd1 vccd1 vccd1 _16209_/A sky130_fd_sc_hd__inv_2
X_11422_ _19562_/Q _11418_/Y _19556_/Q _11419_/Y _11421_/X vssd1 vssd1 vccd1 vccd1
+ _11433_/B sky130_fd_sc_hd__o221a_1
XANTENNA__11024__A1 _11023_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12221__B1 _12035_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15190_ _15190_/A vssd1 vssd1 vccd1 vccd1 _17568_/S sky130_fd_sc_hd__clkinv_8
XANTENNA__16499__C1 _16496_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14141_ _14009_/A _14141_/A2 _14139_/Y _14106_/X vssd1 vssd1 vccd1 vccd1 _18678_/D
+ sky130_fd_sc_hd__a211oi_2
X_11353_ _11479_/A _18981_/Q _11468_/B _18969_/Q _11352_/X vssd1 vssd1 vccd1 vccd1
+ _11361_/B sky130_fd_sc_hd__o221a_1
X_10304_ _18601_/Q _18600_/Q _15621_/A vssd1 vssd1 vccd1 vccd1 _15629_/A sky130_fd_sc_hd__or3_4
XFILLER_4_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14072_ _19061_/Q vssd1 vssd1 vccd1 vccd1 _14072_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19957__RESET_B hold371/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11284_ _19589_/Q _11282_/Y _19604_/Q _11283_/Y vssd1 vssd1 vccd1 vccd1 _11284_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_106_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17900_ _15919_/Y _15920_/Y _15921_/Y _15922_/Y _17913_/S0 _19632_/Q vssd1 vssd1
+ vccd1 vccd1 _17900_/X sky130_fd_sc_hd__mux4_2
X_13023_ _13023_/A _13023_/B _13027_/C vssd1 vssd1 vccd1 vccd1 _18922_/D sky130_fd_sc_hd__nor3_1
X_10235_ _19663_/Q vssd1 vssd1 vccd1 vccd1 _10963_/A sky130_fd_sc_hd__inv_2
XFILLER_79_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18880_ _19814_/CLK _18880_/D repeater223/X vssd1 vssd1 vccd1 vccd1 _18880_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_86_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17831_ _18192_/Q _18184_/Q _18176_/Q _18160_/Q _17918_/S0 _18750_/Q vssd1 vssd1
+ vccd1 vccd1 _17831_/X sky130_fd_sc_hd__mux4_2
XFILLER_39_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10166_ _10174_/A vssd1 vssd1 vccd1 vccd1 _10166_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_output145_A _19764_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17491__S _17545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12288__B1 _12030_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17762_ _17761_/S _13491_/Y _17762_/S vssd1 vssd1 vccd1 vccd1 _17762_/X sky130_fd_sc_hd__mux2_1
X_10097_ _10097_/A vssd1 vssd1 vccd1 vccd1 _10097_/Y sky130_fd_sc_hd__inv_2
X_14974_ _18066_/Q _14965_/A _14842_/X _14966_/A vssd1 vssd1 vccd1 vccd1 _18066_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_235_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19501_ _19510_/CLK hold231/X repeater256/X vssd1 vssd1 vccd1 vccd1 _19501_/Q sky130_fd_sc_hd__dfrtp_1
X_16713_ _16899_/X _16513_/A _16901_/X _16002_/X vssd1 vssd1 vccd1 vccd1 _16713_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_47_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13925_ _13925_/A vssd1 vssd1 vccd1 vccd1 _13925_/X sky130_fd_sc_hd__clkbuf_2
X_17693_ _15460_/X _19442_/Q _17696_/S vssd1 vssd1 vccd1 vccd1 _18559_/D sky130_fd_sc_hd__mux2_1
XFILLER_19_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19432_ _20003_/CLK _19432_/D repeater185/X vssd1 vssd1 vccd1 vccd1 _19432_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__11833__A _12558_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16644_ _16644_/A _16647_/B vssd1 vssd1 vccd1 vccd1 _16644_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__17986__CLK _19851_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13856_ _19217_/Q _18728_/Q _19217_/Q _18728_/Q vssd1 vssd1 vccd1 vccd1 _13856_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_74_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12807_ _19237_/Q _13537_/A _16211_/A _18808_/Q _12806_/X vssd1 vssd1 vccd1 vccd1
+ _12808_/D sky130_fd_sc_hd__o221a_1
XFILLER_50_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19363_ _19984_/CLK _19363_/D repeater243/X vssd1 vssd1 vccd1 vccd1 _19363_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18839__RESET_B repeater233/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16575_ _17202_/X _16394_/X _17205_/X _15898_/X vssd1 vssd1 vccd1 vccd1 _16575_/X
+ sky130_fd_sc_hd__o22a_2
X_13787_ _18725_/Q vssd1 vssd1 vccd1 vccd1 _13909_/A sky130_fd_sc_hd__inv_2
XANTENNA__16835__S _17543_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09456__B2 _19383_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10999_ _19660_/Q _10999_/B vssd1 vssd1 vccd1 vccd1 _10999_/X sky130_fd_sc_hd__or2_1
XFILLER_15_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18314_ _18435_/CLK _18314_/D vssd1 vssd1 vccd1 vccd1 _18314_/Q sky130_fd_sc_hd__dfxtp_1
X_12738_ _16469_/A _18812_/Q _16586_/A _18821_/Q vssd1 vssd1 vccd1 vccd1 _12738_/X
+ sky130_fd_sc_hd__o22a_1
X_15526_ _15526_/A _15526_/B vssd1 vssd1 vccd1 vccd1 _15526_/Y sky130_fd_sc_hd__nor2_1
X_19294_ _20032_/CLK _19294_/D repeater240/X vssd1 vssd1 vccd1 vccd1 _19294_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12460__B1 _12404_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18245_ _19847_/CLK _18245_/D vssd1 vssd1 vccd1 vccd1 _18245_/Q sky130_fd_sc_hd__dfxtp_1
X_15457_ _15457_/A vssd1 vssd1 vccd1 vccd1 _15463_/B sky130_fd_sc_hd__inv_2
XPHY_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12669_ _18987_/Q _12661_/X hold286/X _12664_/X vssd1 vssd1 vccd1 vccd1 _18987_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_187_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14408_ _14450_/A _14450_/B _14571_/C vssd1 vssd1 vccd1 vccd1 _14410_/A sky130_fd_sc_hd__or3_4
XFILLER_129_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15388_ _15388_/A _15388_/B vssd1 vssd1 vccd1 vccd1 _18513_/D sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_144_HCLK clkbuf_4_1_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19847_/CLK sky130_fd_sc_hd__clkbuf_16
X_18176_ _18198_/CLK _18176_/D vssd1 vssd1 vccd1 vccd1 _18176_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_190_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17666__S _17683_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14339_ _18433_/Q _14336_/X _14273_/X _14338_/X vssd1 vssd1 vccd1 vccd1 _18433_/D
+ sky130_fd_sc_hd__a22o_1
X_17127_ _17486_/A0 _09914_/Y _17543_/S vssd1 vssd1 vccd1 vccd1 _17127_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17058_ _17057_/X _15683_/A _17318_/S vssd1 vssd1 vccd1 vccd1 _17058_/X sky130_fd_sc_hd__mux2_1
XANTENNA__19737__CLK _20051_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11318__A2 _18973_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16009_ _18028_/Q vssd1 vssd1 vccd1 vccd1 _16009_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19627__RESET_B repeater261/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09880_ _19340_/Q vssd1 vssd1 vccd1 vccd1 _09880_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_4_7_0_HCLK clkbuf_4_7_0_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_7_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_100_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19887__CLK _20051_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12279__B1 _12098_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20114__RESET_B repeater217/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12558__B _12558_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09314_ _18658_/Q _09329_/A _09302_/A vssd1 vssd1 vccd1 vccd1 _15725_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__18509__RESET_B repeater222/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15869__B _15878_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18141__CLK _19510_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09245_ _09253_/S vssd1 vssd1 vccd1 vccd1 _09250_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_194_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12203__B1 _12090_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09176_ _20077_/Q vssd1 vssd1 vccd1 vccd1 _14709_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_181_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17576__S _17584_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16496__A2 _15896_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11309__A2 _18968_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19368__RESET_B repeater241/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11918__A _12232_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10822__A _10831_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold290_A HWDATA[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10020_ _10045_/A _10044_/A _10047_/A _10046_/A vssd1 vssd1 vccd1 vccd1 _10021_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_48_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_25_HCLK clkbuf_4_9_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20050_/CLK sky130_fd_sc_hd__clkbuf_16
X_11971_ _19377_/Q _11969_/X _09071_/X _11970_/X vssd1 vssd1 vccd1 vccd1 _19377_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_29_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13710_ _17761_/X _13710_/B vssd1 vssd1 vccd1 vccd1 _13710_/Y sky130_fd_sc_hd__nand2_1
X_10922_ _18510_/Q _10922_/B vssd1 vssd1 vccd1 vccd1 _19681_/D sky130_fd_sc_hd__or2_1
X_14690_ _18228_/Q _14683_/A _14582_/X _14684_/A vssd1 vssd1 vccd1 vccd1 _18228_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12690__B1 _12032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_244_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13641_ _13641_/A _13641_/B vssd1 vssd1 vccd1 vccd1 _15233_/B sky130_fd_sc_hd__or2_2
XFILLER_71_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10853_ _19709_/Q _10844_/A _10427_/X _10845_/A vssd1 vssd1 vccd1 vccd1 _19709_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_32_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_232_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16360_ _18088_/Q vssd1 vssd1 vccd1 vccd1 _16360_/Y sky130_fd_sc_hd__inv_2
X_13572_ _13551_/A _13572_/A2 _13571_/X _13569_/Y vssd1 vssd1 vccd1 vccd1 _18828_/D
+ sky130_fd_sc_hd__a211oi_4
XFILLER_13_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10784_ _10805_/A _19741_/Q _19740_/Q vssd1 vssd1 vccd1 vccd1 _19741_/D sky130_fd_sc_hd__a21o_1
XFILLER_188_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_135_HCLK_A clkbuf_4_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_212_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15311_ _15311_/A _18551_/Q vssd1 vssd1 vccd1 vccd1 _15753_/B sky130_fd_sc_hd__or2_2
XFILLER_169_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12523_ hold268/X vssd1 vssd1 vccd1 vccd1 hold267/A sky130_fd_sc_hd__clkbuf_4
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16291_ _18801_/Q _15957_/Y _18800_/Q _15819_/Y vssd1 vssd1 vccd1 vccd1 _16291_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_200_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15242_ _18633_/Q vssd1 vssd1 vccd1 vccd1 _15242_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18634__CLK _19780_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18030_ _18142_/CLK _18030_/D vssd1 vssd1 vccd1 vccd1 _18030_/Q sky130_fd_sc_hd__dfxtp_1
X_12454_ _19117_/Q _12450_/X _12394_/X _12451_/X vssd1 vssd1 vccd1 vccd1 _19117_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_126_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11405_ _11548_/B _19128_/Q _11547_/B _19153_/Q _11404_/X vssd1 vssd1 vccd1 vccd1
+ _11412_/C sky130_fd_sc_hd__o221a_1
XANTENNA__17486__S _17543_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15173_ _17944_/Q _15170_/X hold247/X _15172_/X vssd1 vssd1 vccd1 vccd1 _17944_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17133__A0 _17486_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12385_ _19154_/Q _12374_/X _12384_/X _12378_/X vssd1 vssd1 vccd1 vccd1 _19154_/D
+ sky130_fd_sc_hd__a22o_1
X_14124_ _18689_/Q _14123_/Y _14124_/B1 _14112_/X vssd1 vssd1 vccd1 vccd1 _18689_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__19791__RESET_B repeater203/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11336_ _19599_/Q _11332_/Y _19595_/Q _11333_/Y _11335_/X vssd1 vssd1 vccd1 vccd1
+ _11347_/A sky130_fd_sc_hd__o221a_1
XFILLER_4_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16487__A2 _16505_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19981_ _19992_/CLK _19981_/D repeater192/X vssd1 vssd1 vccd1 vccd1 _19981_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_207_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14055_ _19074_/Q _18685_/Q _14054_/Y _14015_/A vssd1 vssd1 vccd1 vccd1 _14055_/X
+ sky130_fd_sc_hd__o22a_1
X_18932_ _19325_/CLK _18932_/D repeater215/X vssd1 vssd1 vccd1 vccd1 _18932_/Q sky130_fd_sc_hd__dfrtp_1
X_11267_ _11478_/A _19012_/Q _11485_/A _19019_/Q _11266_/X vssd1 vssd1 vccd1 vccd1
+ _11299_/B sky130_fd_sc_hd__o221a_1
XFILLER_97_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13006_ _13006_/A _13006_/B vssd1 vssd1 vccd1 vccd1 _13011_/A sky130_fd_sc_hd__or2_1
X_10218_ _19827_/Q vssd1 vssd1 vccd1 vccd1 _10218_/Y sky130_fd_sc_hd__inv_2
X_18863_ _18866_/CLK _18863_/D repeater231/X vssd1 vssd1 vccd1 vccd1 _18863_/Q sky130_fd_sc_hd__dfrtp_1
X_11198_ _17720_/X _11191_/A _19611_/Q _11192_/A vssd1 vssd1 vccd1 vccd1 _19611_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_223_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18014__CLK _18169_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17814_ _17810_/X _17811_/X _17812_/X _17813_/X _18751_/Q _18752_/Q vssd1 vssd1 vccd1
+ vccd1 _17814_/X sky130_fd_sc_hd__mux4_2
X_10149_ _12370_/A _12130_/B _12370_/C vssd1 vssd1 vccd1 vccd1 _15883_/A sky130_fd_sc_hd__or3_4
X_18794_ _19647_/CLK _18794_/D repeater261/X vssd1 vssd1 vccd1 vccd1 _18794_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_67_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17745_ _17764_/S _13289_/Y _17763_/S vssd1 vssd1 vccd1 vccd1 _17745_/X sky130_fd_sc_hd__mux2_1
XFILLER_236_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14957_ _18079_/Q _14952_/X _14927_/X _14954_/X vssd1 vssd1 vccd1 vccd1 _18079_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12659__A _12659_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13908_ _18733_/Q _13916_/A _13907_/X _13832_/B vssd1 vssd1 vccd1 vccd1 _18733_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12681__B1 hold318/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17676_ _15532_/Y _19459_/Q _17683_/S vssd1 vssd1 vccd1 vccd1 _18576_/D sky130_fd_sc_hd__mux2_1
X_14888_ _18119_/Q _14883_/X _14808_/X _14885_/X vssd1 vssd1 vccd1 vccd1 _18119_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_63_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_15_0_HCLK clkbuf_3_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_4_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09033__A hold308/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19415_ _19984_/CLK _19415_/D repeater193/X vssd1 vssd1 vccd1 vccd1 _19415_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16627_ _16978_/X _16594_/X _16976_/X _16595_/X vssd1 vssd1 vccd1 vccd1 _16629_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18673__RESET_B repeater252/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13839_ _13838_/Y _18730_/Q _19197_/Q _13945_/A vssd1 vssd1 vccd1 vccd1 _13839_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_51_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19346_ _19952_/CLK _19346_/D repeater245/X vssd1 vssd1 vccd1 vccd1 _19346_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_15_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12433__B1 _12236_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16558_ _17163_/X _16555_/X _17154_/X _16556_/X _16557_/X vssd1 vssd1 vccd1 vccd1
+ _16558_/Y sky130_fd_sc_hd__a221oi_2
X_15509_ _18572_/Q _15509_/B vssd1 vssd1 vccd1 vccd1 _15518_/C sky130_fd_sc_hd__or2_2
X_19277_ _19315_/CLK _19277_/D repeater215/X vssd1 vssd1 vccd1 vccd1 _19277_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12394__A hold306/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16489_ _19887_/Q vssd1 vssd1 vccd1 vccd1 _16489_/Y sky130_fd_sc_hd__inv_2
X_09030_ hold303/X vssd1 vssd1 vccd1 vccd1 _09030_/X sky130_fd_sc_hd__buf_4
XFILLER_164_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18228_ _18412_/CLK _18228_/D vssd1 vssd1 vccd1 vccd1 _18228_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_248_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_57_HCLK_A clkbuf_4_12_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17396__S _17565_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18159_ _18198_/CLK _18159_/D vssd1 vssd1 vccd1 vccd1 _18159_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10747__B1 _10418_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold302 HWDATA[20] vssd1 vssd1 vccd1 vccd1 input50/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold313 MSI_S3 vssd1 vssd1 vccd1 vccd1 input72/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold324 hold324/A vssd1 vssd1 vccd1 vccd1 hold324/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16478__A2 _16597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold335 hold335/A vssd1 vssd1 vccd1 vccd1 hold335/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold346 hold346/A vssd1 vssd1 vccd1 vccd1 hold346/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold357 hold357/A vssd1 vssd1 vccd1 vccd1 hold357/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20121_ _20122_/CLK _20121_/D repeater234/X vssd1 vssd1 vccd1 vccd1 _20121_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17770__S1 _19646_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold368 hold368/A vssd1 vssd1 vccd1 vccd1 hold368/X sky130_fd_sc_hd__dlygate4sd3_1
X_09932_ _19951_/Q _09930_/Y _19959_/Q _16621_/A vssd1 vssd1 vccd1 vccd1 _09932_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_89_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15150__A2 _15146_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20052_ _20055_/CLK _20052_/D repeater207/X vssd1 vssd1 vccd1 vccd1 _20052_/Q sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_48_HCLK clkbuf_opt_2_HCLK/A vssd1 vssd1 vccd1 vccd1 _19825_/CLK sky130_fd_sc_hd__clkbuf_16
X_09863_ _09863_/A _09863_/B vssd1 vssd1 vccd1 vccd1 _09975_/A sky130_fd_sc_hd__or2_1
XFILLER_58_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09794_ _09794_/A _09794_/B vssd1 vssd1 vccd1 vccd1 _09794_/Y sky130_fd_sc_hd__nor2_2
XFILLER_245_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrepeater152 _17385_/S vssd1 vssd1 vccd1 vccd1 _17535_/S sky130_fd_sc_hd__buf_8
XFILLER_27_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater163 _17042_/S vssd1 vssd1 vccd1 vccd1 _17512_/S sky130_fd_sc_hd__buf_6
Xrepeater174 _17474_/S vssd1 vssd1 vccd1 vccd1 _17318_/S sky130_fd_sc_hd__buf_8
XPHY_4306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater185 hold371/X vssd1 vssd1 vccd1 vccd1 repeater185/X sky130_fd_sc_hd__buf_6
XPHY_4317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater196 repeater197/X vssd1 vssd1 vccd1 vccd1 repeater196/X sky130_fd_sc_hd__buf_6
XANTENNA__12672__B1 hold303/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12424__B1 _12223_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19902__CLK _20123_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17363__A0 _15768_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09228_ _15709_/A _09226_/X _18646_/Q _09227_/Y vssd1 vssd1 vccd1 vccd1 _15711_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_194_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09159_ _15321_/A _15322_/B _09146_/A vssd1 vssd1 vccd1 vccd1 _09159_/X sky130_fd_sc_hd__o21a_1
XANTENNA__19549__RESET_B repeater269/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17115__A0 _17473_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16504__A _16504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12170_ _19269_/Q _12164_/X _11975_/X _12165_/X vssd1 vssd1 vccd1 vccd1 _19269_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11121_ _11094_/Y _19635_/Q _11094_/Y _19635_/Q vssd1 vssd1 vccd1 vccd1 _19635_/D
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__18037__CLK _19851_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11052_ _11147_/A _14301_/B vssd1 vssd1 vccd1 vccd1 _11053_/B sky130_fd_sc_hd__or2_1
XFILLER_89_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10003_ _19939_/Q _09734_/A _10001_/A _09964_/X vssd1 vssd1 vccd1 vccd1 _19939_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_131_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15860_ _15851_/X _15857_/X _15859_/X vssd1 vssd1 vccd1 vccd1 _15860_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__10910__B1 _17936_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input21_A HADDR[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14811_ _18166_/Q _14801_/X _14810_/X _14804_/X vssd1 vssd1 vccd1 vccd1 _18166_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_218_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15791_ _18010_/Q vssd1 vssd1 vccd1 vccd1 _15791_/Y sky130_fd_sc_hd__inv_2
XFILLER_190_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17530_ _17529_/X _09465_/A _17530_/S vssd1 vssd1 vccd1 vccd1 _17530_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_233_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11954_ _11954_/A1 _11948_/X _09039_/X _11949_/X vssd1 vssd1 vccd1 vccd1 _19388_/D
+ sky130_fd_sc_hd__a22o_1
X_14742_ _18202_/Q _14733_/A _14693_/X _14734_/A vssd1 vssd1 vccd1 vccd1 _18202_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_123_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10905_ _15208_/B vssd1 vssd1 vccd1 vccd1 _15215_/B sky130_fd_sc_hd__buf_1
XFILLER_60_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17461_ _16046_/X _20042_/Q _19498_/Q vssd1 vssd1 vccd1 vccd1 _17461_/X sky130_fd_sc_hd__mux2_1
X_14673_ _18240_/Q _14669_/X _09171_/X _14671_/X vssd1 vssd1 vccd1 vccd1 _18240_/D
+ sky130_fd_sc_hd__a22o_1
X_11885_ _11892_/A vssd1 vssd1 vccd1 vccd1 _11885_/X sky130_fd_sc_hd__buf_1
XFILLER_33_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output108_A _16465_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19200_ _19585_/CLK _19200_/D hold367/X vssd1 vssd1 vccd1 vccd1 _19200_/Q sky130_fd_sc_hd__dfrtp_1
X_16412_ _18473_/Q vssd1 vssd1 vccd1 vccd1 _16412_/Y sky130_fd_sc_hd__inv_2
X_13624_ _18803_/Q _13623_/X _18803_/Q _13623_/X vssd1 vssd1 vccd1 vccd1 _18803_/D
+ sky130_fd_sc_hd__o2bb2a_1
X_10836_ _10836_/A vssd1 vssd1 vccd1 vccd1 _19719_/D sky130_fd_sc_hd__inv_2
XANTENNA__12415__B1 _12413_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17392_ _17391_/X _19130_/Q _17548_/S vssd1 vssd1 vccd1 vccd1 _17392_/X sky130_fd_sc_hd__mux2_2
XFILLER_186_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19131_ _19970_/CLK _19131_/D repeater249/X vssd1 vssd1 vccd1 vccd1 _19131_/Q sky130_fd_sc_hd__dfrtp_4
X_13555_ _13555_/A _13555_/B vssd1 vssd1 vccd1 vccd1 _13563_/A sky130_fd_sc_hd__or2_1
XANTENNA__17354__A0 _15963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16343_ _18048_/Q vssd1 vssd1 vccd1 vccd1 _16343_/Y sky130_fd_sc_hd__inv_2
XANTENNA_repeater160_A _17493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10767_ _19751_/Q _10767_/B vssd1 vssd1 vccd1 vccd1 _10767_/Y sky130_fd_sc_hd__nand2_1
XFILLER_185_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12506_ _12506_/A vssd1 vssd1 vccd1 vccd1 _12506_/X sky130_fd_sc_hd__clkbuf_2
X_19062_ _19608_/CLK _19062_/D hold355/X vssd1 vssd1 vccd1 vccd1 _19062_/Q sky130_fd_sc_hd__dfrtp_4
X_16274_ _17378_/X _16415_/B vssd1 vssd1 vccd1 vccd1 _16274_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__19972__RESET_B hold371/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13486_ _13486_/A vssd1 vssd1 vccd1 vccd1 _13489_/A sky130_fd_sc_hd__inv_2
X_10698_ _14791_/A vssd1 vssd1 vccd1 vccd1 _10698_/X sky130_fd_sc_hd__buf_4
X_15225_ _18635_/Q vssd1 vssd1 vccd1 vccd1 _15278_/B sky130_fd_sc_hd__inv_2
X_18013_ _18165_/CLK _18013_/D vssd1 vssd1 vccd1 vccd1 _18013_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12437_ _12487_/B _15863_/B vssd1 vssd1 vccd1 vccd1 _12438_/S sky130_fd_sc_hd__or2_1
XANTENNA__19901__RESET_B repeater195/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10729__B1 _10425_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15156_ _17953_/Q _15147_/A _14949_/X _15148_/A vssd1 vssd1 vccd1 vccd1 _17953_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_114_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12368_ _19159_/Q _12334_/A _12238_/X _12335_/A vssd1 vssd1 vccd1 vccd1 _19159_/D
+ sky130_fd_sc_hd__a22o_1
X_14107_ _14028_/A _14107_/A2 _14106_/X _14104_/Y vssd1 vssd1 vccd1 vccd1 _18698_/D
+ sky130_fd_sc_hd__a211oi_2
X_11319_ _19580_/Q _11316_/Y _11461_/A _18962_/Q _11318_/X vssd1 vssd1 vccd1 vccd1
+ _11319_/X sky130_fd_sc_hd__a221o_1
XFILLER_180_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15087_ _18000_/Q _15083_/X hold236/X _15085_/X vssd1 vssd1 vccd1 vccd1 _18000_/D
+ sky130_fd_sc_hd__a22o_1
X_19964_ _19964_/CLK _19964_/D repeater185/X vssd1 vssd1 vccd1 vccd1 _19964_/Q sky130_fd_sc_hd__dfrtp_4
X_12299_ _14277_/A vssd1 vssd1 vccd1 vccd1 _12299_/X sky130_fd_sc_hd__buf_2
XFILLER_234_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13143__A1 _19168_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14038_ _19079_/Q vssd1 vssd1 vccd1 vccd1 _14038_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14340__B1 _14277_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18915_ _19222_/CLK _18915_/D repeater186/X vssd1 vssd1 vccd1 vccd1 _18915_/Q sky130_fd_sc_hd__dfrtp_1
X_19895_ _20055_/CLK _19895_/D repeater205/X vssd1 vssd1 vccd1 vccd1 _19895_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_68_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11154__B1 _11153_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18846_ _18866_/CLK _18846_/D repeater233/X vssd1 vssd1 vccd1 vccd1 _18846_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_227_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10901__B1 _10866_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13492__B _15858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18854__RESET_B repeater231/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18777_ _19847_/CLK _18777_/D repeater264/X vssd1 vssd1 vccd1 vccd1 _18777_/Q sky130_fd_sc_hd__dfrtp_1
X_15989_ _15980_/Y _15864_/B _15982_/X _15988_/X vssd1 vssd1 vccd1 vccd1 _15989_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12389__A hold303/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_243_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17728_ _17936_/Q _19685_/Q _18510_/Q vssd1 vssd1 vccd1 vccd1 _17728_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12654__B1 _12533_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17659_ _15599_/X _19030_/Q _17664_/S vssd1 vssd1 vccd1 vccd1 _18593_/D sky130_fd_sc_hd__mux2_1
XANTENNA__16396__A1 _11742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19329_ _19513_/CLK _19329_/D repeater259/X vssd1 vssd1 vccd1 vccd1 _19329_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_148_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09013_ _12187_/A _12659_/A vssd1 vssd1 vccd1 vccd1 _09084_/A sky130_fd_sc_hd__or2_4
XANTENNA__19642__RESET_B repeater261/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold132 hold132/A vssd1 vssd1 vccd1 vccd1 hold132/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold143 HADDR[20] vssd1 vssd1 vccd1 vccd1 input13/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_160_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold154 HADDR[17] vssd1 vssd1 vccd1 vccd1 input9/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 input5/X vssd1 vssd1 vccd1 vccd1 hold165/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 hold176/A vssd1 vssd1 vccd1 vccd1 hold176/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09338__B1 _20038_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold187 HADDR[7] vssd1 vssd1 vccd1 vccd1 input30/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_120_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20104_ _20107_/CLK _20104_/D repeater233/X vssd1 vssd1 vccd1 vccd1 _20104_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__14331__B1 _14312_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold198 hold198/A vssd1 vssd1 vccd1 vccd1 hold198/X sky130_fd_sc_hd__dlygate4sd3_1
X_09915_ _09862_/A _19346_/Q _19954_/Q _09914_/Y vssd1 vssd1 vccd1 vccd1 _09915_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_58_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20035_ _20035_/CLK _20035_/D repeater216/X vssd1 vssd1 vccd1 vccd1 _20035_/Q sky130_fd_sc_hd__dfrtp_1
X_09846_ _19940_/Q vssd1 vssd1 vccd1 vccd1 _09849_/A sky130_fd_sc_hd__inv_2
XFILLER_59_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18595__RESET_B repeater269/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09777_ _09746_/A _09746_/B _09767_/X _09775_/Y vssd1 vssd1 vccd1 vccd1 _19990_/D
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__12299__A _14277_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12645__B1 hold239/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11931__A _11933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11670_ _19543_/Q _11668_/X _11651_/A _11669_/X vssd1 vssd1 vccd1 vccd1 _19543_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10621_ _19809_/Q vssd1 vssd1 vccd1 vccd1 _10939_/B sky130_fd_sc_hd__inv_2
XPHY_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17336__A0 _15768_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16933__S _16946_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13340_ _13429_/D _13340_/B vssd1 vssd1 vccd1 vccd1 _13453_/A sky130_fd_sc_hd__or2_1
XFILLER_10_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10552_ _10583_/A _10552_/B vssd1 vssd1 vccd1 vccd1 _10553_/A sky130_fd_sc_hd__or2_2
XFILLER_183_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13271_ _13256_/X _13262_/B _13737_/B vssd1 vssd1 vccd1 vccd1 _13271_/Y sky130_fd_sc_hd__o21ai_1
X_10483_ _10734_/A vssd1 vssd1 vccd1 vccd1 _11655_/A sky130_fd_sc_hd__buf_1
XANTENNA_clkbuf_leaf_40_HCLK_A clkbuf_opt_1_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15010_ _15011_/A vssd1 vssd1 vccd1 vccd1 _15010_/X sky130_fd_sc_hd__clkbuf_2
X_12222_ _19237_/Q _12219_/X _12038_/X _12220_/X vssd1 vssd1 vccd1 vccd1 _19237_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_182_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14570__B1 hold320/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12153_ _19282_/Q _12150_/X _12098_/X _12151_/X vssd1 vssd1 vccd1 vccd1 _19282_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_162_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11104_ _11093_/Y _17755_/X _11091_/X _11103_/X vssd1 vssd1 vccd1 vccd1 _19639_/D
+ sky130_fd_sc_hd__o22ai_1
XANTENNA__14322__B1 _14277_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16961_ _16960_/X _13362_/Y _17535_/S vssd1 vssd1 vccd1 vccd1 _16961_/X sky130_fd_sc_hd__mux2_1
X_12084_ _12096_/A vssd1 vssd1 vccd1 vccd1 _12084_/X sky130_fd_sc_hd__buf_1
X_18700_ _18701_/CLK _18700_/D hold359/X vssd1 vssd1 vccd1 vccd1 _18700_/Q sky130_fd_sc_hd__dfrtp_1
X_11035_ _19649_/Q _11025_/B _11026_/A _11029_/Y vssd1 vssd1 vccd1 vccd1 _11035_/X
+ sky130_fd_sc_hd__o211a_1
X_15912_ _16509_/A vssd1 vssd1 vccd1 vccd1 _16683_/A sky130_fd_sc_hd__clkbuf_4
X_19680_ _19795_/CLK _19680_/D repeater218/X vssd1 vssd1 vccd1 vccd1 _19680_/Q sky130_fd_sc_hd__dfrtp_2
X_16892_ _17486_/A0 _13114_/Y _17543_/S vssd1 vssd1 vccd1 vccd1 _16892_/X sky130_fd_sc_hd__mux2_1
XFILLER_209_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19948__CLK _19976_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16075__B1 _17451_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18631_ _19780_/CLK _18631_/D repeater225/X vssd1 vssd1 vccd1 vccd1 _18631_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_94_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15843_ _15735_/A _15840_/X _15841_/Y _15842_/X vssd1 vssd1 vccd1 vccd1 _15843_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_225_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18562_ _20058_/CLK _18562_/D repeater194/X vssd1 vssd1 vccd1 vccd1 _18562_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_218_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12986_ _12986_/A vssd1 vssd1 vccd1 vccd1 _12986_/X sky130_fd_sc_hd__buf_2
X_15774_ _15774_/A vssd1 vssd1 vccd1 vccd1 _17548_/S sky130_fd_sc_hd__inv_16
XFILLER_205_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17513_ _17512_/X _15581_/B _17513_/S vssd1 vssd1 vccd1 vccd1 _17513_/X sky130_fd_sc_hd__mux2_2
X_14725_ _14793_/A vssd1 vssd1 vccd1 vccd1 _14725_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_233_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18493_ _20057_/CLK _18493_/D repeater202/X vssd1 vssd1 vccd1 vccd1 _18493_/Q sky130_fd_sc_hd__dfrtp_1
X_11937_ _15772_/A _12066_/A vssd1 vssd1 vccd1 vccd1 _11977_/A sky130_fd_sc_hd__or2_4
XANTENNA__17004__S _17318_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11841__A _12313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17444_ _17443_/X _09691_/Y _17517_/S vssd1 vssd1 vccd1 vccd1 _17444_/X sky130_fd_sc_hd__mux2_1
XFILLER_220_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11868_ _11851_/A _11867_/X _11865_/X vssd1 vssd1 vccd1 vccd1 _19434_/D sky130_fd_sc_hd__a21boi_1
X_14656_ _14657_/A vssd1 vssd1 vccd1 vccd1 _14656_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_221_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13607_ _13607_/A vssd1 vssd1 vccd1 vccd1 _13607_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17327__A0 _15963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10819_ _10819_/A _12370_/B _12130_/C vssd1 vssd1 vccd1 vccd1 _15845_/D sky130_fd_sc_hd__or3_4
XFILLER_20_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17375_ _16274_/Y _10203_/Y _17566_/S vssd1 vssd1 vccd1 vccd1 _17375_/X sky130_fd_sc_hd__mux2_1
XFILLER_220_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14587_ _14588_/A vssd1 vssd1 vccd1 vccd1 _14587_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__16843__S _17493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11799_ _19461_/Q _11793_/X _09039_/X _11794_/X vssd1 vssd1 vccd1 vccd1 _19461_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_229_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19114_ _19115_/CLK _19114_/D hold353/X vssd1 vssd1 vccd1 vccd1 _19114_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_201_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16326_ _15749_/B _16320_/X _16322_/X _16324_/X _16325_/X vssd1 vssd1 vccd1 vccd1
+ _16326_/X sky130_fd_sc_hd__o2111a_1
X_13538_ _13538_/A _13538_/B vssd1 vssd1 vccd1 vccd1 _13539_/B sky130_fd_sc_hd__or2_2
X_19045_ _19566_/CLK _19045_/D repeater255/X vssd1 vssd1 vccd1 vccd1 _19045_/Q sky130_fd_sc_hd__dfrtp_1
X_13469_ _13469_/A _13473_/A vssd1 vssd1 vccd1 vccd1 _13470_/B sky130_fd_sc_hd__or2_2
X_16257_ _18071_/Q vssd1 vssd1 vccd1 vccd1 _16257_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15208_ _15208_/A _15208_/B vssd1 vssd1 vccd1 vccd1 _15208_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__19053__RESET_B repeater267/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16188_ _17981_/Q vssd1 vssd1 vccd1 vccd1 _16188_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17674__S _17683_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15139_ _17966_/Q _15134_/X hold244/X _15136_/X vssd1 vssd1 vccd1 vccd1 _17966_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_126_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14313__B1 _14312_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19947_ _19956_/CLK _19947_/D hold371/X vssd1 vssd1 vccd1 vccd1 _19947_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09700_ _19408_/Q vssd1 vssd1 vccd1 vccd1 _09700_/Y sky130_fd_sc_hd__inv_2
XFILLER_229_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19878_ _20059_/CLK _19878_/D repeater199/X vssd1 vssd1 vccd1 vccd1 _19878_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_95_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16605__A2 _15889_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09631_ _19976_/Q vssd1 vssd1 vccd1 vccd1 _09788_/A sky130_fd_sc_hd__inv_2
X_18829_ _19255_/CLK _18829_/D repeater237/X vssd1 vssd1 vccd1 vccd1 _18829_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_228_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09562_ _20035_/Q _09560_/Y _20028_/Q _16670_/A vssd1 vssd1 vccd1 vccd1 _09562_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12627__B1 _12396_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14092__A2 _18673_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09493_ _09493_/A _09571_/A vssd1 vssd1 vccd1 vccd1 _09494_/B sky130_fd_sc_hd__or2_2
XFILLER_36_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11751__A _11772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19894__RESET_B repeater205/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13678__A _13678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16541__A1 _15199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_191_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14552__B1 _14509_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17584__S _17584_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18845__CLK _18866_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18705__RESET_B repeater253/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20018_ _20091_/CLK _20018_/D repeater236/X vssd1 vssd1 vccd1 vccd1 _20018_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_247_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09829_ _19957_/Q vssd1 vssd1 vccd1 vccd1 _09865_/A sky130_fd_sc_hd__inv_2
XFILLER_207_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16928__S _16946_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12840_ _18944_/Q vssd1 vssd1 vccd1 vccd1 _12887_/A sky130_fd_sc_hd__inv_2
XANTENNA__12618__B1 _12380_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12771_ _18804_/Q vssd1 vssd1 vccd1 vccd1 _13528_/A sky130_fd_sc_hd__inv_2
XPHY_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11722_ _19511_/Q _11716_/X _16943_/X _11717_/X vssd1 vssd1 vccd1 vccd1 hold220/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_54_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14510_ _18334_/Q _14503_/X _14509_/X _14505_/X vssd1 vssd1 vccd1 vccd1 _18334_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__15133__A _15169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15490_ _15490_/A vssd1 vssd1 vccd1 vccd1 _15490_/Y sky130_fd_sc_hd__inv_2
XFILLER_242_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_203_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11653_ _11653_/A _11653_/B vssd1 vssd1 vccd1 vccd1 _15389_/C sky130_fd_sc_hd__or2_1
X_14441_ _14749_/A vssd1 vssd1 vccd1 vccd1 _14441_/X sky130_fd_sc_hd__clkbuf_2
XPHY_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16780__A1 _19395_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10604_ _10618_/A vssd1 vssd1 vccd1 vccd1 _10617_/A sky130_fd_sc_hd__inv_2
XFILLER_168_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17160_ _17159_/X _09442_/Y _17529_/S vssd1 vssd1 vccd1 vccd1 _17160_/X sky130_fd_sc_hd__mux2_1
X_14372_ _18415_/Q _14367_/X _14359_/X _14369_/X vssd1 vssd1 vccd1 vccd1 _18415_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11584_ _11584_/A _11597_/A _11584_/C vssd1 vssd1 vccd1 vccd1 _11594_/A sky130_fd_sc_hd__or3_4
XPHY_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13323_ _18844_/Q vssd1 vssd1 vccd1 vccd1 _13467_/A sky130_fd_sc_hd__inv_1
XPHY_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16111_ _18101_/Q vssd1 vssd1 vccd1 vccd1 _16111_/Y sky130_fd_sc_hd__inv_2
X_10535_ _15289_/A vssd1 vssd1 vccd1 vccd1 _11648_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_13_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19620__CLK _19920_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17091_ _17090_/X _12913_/Y _17487_/S vssd1 vssd1 vccd1 vccd1 _17091_/X sky130_fd_sc_hd__mux2_1
XANTENNA__16532__A1 _17161_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14543__B1 _14474_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16042_ _18769_/Q vssd1 vssd1 vccd1 vccd1 _16042_/Y sky130_fd_sc_hd__inv_2
X_13254_ _18870_/Q vssd1 vssd1 vccd1 vccd1 _13254_/Y sky130_fd_sc_hd__inv_2
X_10466_ _19823_/Q _10472_/A vssd1 vssd1 vccd1 vccd1 _10466_/X sky130_fd_sc_hd__or2_1
XFILLER_142_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12205_ _12205_/A vssd1 vssd1 vccd1 vccd1 _12205_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__17494__S _17548_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13185_ _18906_/Q _13184_/Y _13180_/X _13185_/C1 vssd1 vssd1 vccd1 vccd1 _18906_/D
+ sky130_fd_sc_hd__o211a_1
X_10397_ _19851_/Q vssd1 vssd1 vccd1 vccd1 _14990_/A sky130_fd_sc_hd__buf_1
XFILLER_123_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19801_ _19812_/CLK _19801_/D repeater222/X vssd1 vssd1 vccd1 vccd1 _19801_/Q sky130_fd_sc_hd__dfrtp_4
X_12136_ _12172_/A vssd1 vssd1 vccd1 vccd1 _12151_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_150_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17993_ _18169_/CLK _17993_/D vssd1 vssd1 vccd1 vccd1 _17993_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_215_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19732_ _20057_/CLK _19732_/D repeater202/X vssd1 vssd1 vccd1 vccd1 _19732_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__11836__A _11996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12067_ _12121_/A vssd1 vssd1 vccd1 vccd1 _12094_/A sky130_fd_sc_hd__clkbuf_2
X_16944_ _19488_/Q hold153/X _16946_/S vssd1 vssd1 vccd1 vccd1 _16944_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10740__A _15826_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11018_ _10408_/X _10956_/C _10973_/B _11017_/X vssd1 vssd1 vccd1 vccd1 _19655_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_49_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19663_ _19668_/CLK _19663_/D repeater270/X vssd1 vssd1 vccd1 vccd1 _19663_/Q sky130_fd_sc_hd__dfrtp_1
X_16875_ _16874_/X _13080_/A _17542_/S vssd1 vssd1 vccd1 vccd1 _16875_/X sky130_fd_sc_hd__mux2_2
XANTENNA__16838__S _17547_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_237_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18614_ _19157_/CLK _18614_/D repeater266/X vssd1 vssd1 vccd1 vccd1 _18614_/Q sky130_fd_sc_hd__dfrtp_1
X_15826_ _15826_/A vssd1 vssd1 vccd1 vccd1 _15866_/A sky130_fd_sc_hd__clkbuf_2
X_19594_ _19595_/CLK _19594_/D hold346/A vssd1 vssd1 vccd1 vccd1 _19594_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__17891__S0 _17913_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_237_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18545_ _18545_/CLK _18545_/D repeater232/X vssd1 vssd1 vccd1 vccd1 _18545_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_18_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15757_ _18883_/Q _18881_/Q _18882_/Q _15756_/X vssd1 vssd1 vccd1 vccd1 _18524_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17548__A0 _17547_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12969_ _12967_/X _18943_/Q _18944_/Q _12969_/D vssd1 vssd1 vccd1 vccd1 _12970_/C
+ sky130_fd_sc_hd__and4b_1
XFILLER_205_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14708_ _18222_/Q _14698_/X _14707_/X _14701_/X vssd1 vssd1 vccd1 vccd1 _18222_/D
+ sky130_fd_sc_hd__a22o_1
X_18476_ _20064_/CLK _18476_/D repeater198/X vssd1 vssd1 vccd1 vccd1 _18476_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_205_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15688_ _15688_/A _15688_/B vssd1 vssd1 vccd1 vccd1 _15688_/Y sky130_fd_sc_hd__nor2_1
XFILLER_60_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17669__S _17683_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17427_ _16118_/X _20043_/Q _19498_/Q vssd1 vssd1 vccd1 vccd1 _17427_/X sky130_fd_sc_hd__mux2_1
X_14639_ _18259_/Q _14631_/A _09185_/X _14632_/A vssd1 vssd1 vccd1 vccd1 _18259_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_147_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17358_ _17357_/X _13406_/Y _17529_/S vssd1 vssd1 vccd1 vccd1 _17358_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_186_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16309_ _16305_/Y _15971_/X _16306_/Y _15973_/X _16308_/X vssd1 vssd1 vccd1 vccd1
+ _16309_/X sky130_fd_sc_hd__o221a_1
XANTENNA__13498__A _15195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17289_ _17288_/X _09424_/Y _17413_/S vssd1 vssd1 vccd1 vccd1 _17289_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19028_ _19667_/CLK _19028_/D repeater269/X vssd1 vssd1 vccd1 vccd1 _19028_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_126_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08993_ _19515_/Q vssd1 vssd1 vccd1 vccd1 _09259_/B sky130_fd_sc_hd__inv_2
XFILLER_130_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_229_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09614_ _09469_/A _09616_/C1 _09612_/Y _09607_/X vssd1 vssd1 vccd1 vccd1 _20008_/D
+ sky130_fd_sc_hd__a211oi_4
XANTENNA__18248__CLK _19847_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17882__S0 _17913_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_232_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09545_ _09545_/A _09545_/B _09545_/C _09545_/D vssd1 vssd1 vccd1 vccd1 _09565_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_52_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09476_ _09476_/A _09476_/B vssd1 vssd1 vccd1 vccd1 _09598_/A sky130_fd_sc_hd__or2_1
XFILLER_240_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17579__S _17584_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10320_ _10368_/A vssd1 vssd1 vccd1 vccd1 _10320_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__14525__B1 hold330/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18957__RESET_B repeater257/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10251_ _10819_/A _11935_/B _12130_/C vssd1 vssd1 vccd1 vccd1 _15899_/A sky130_fd_sc_hd__or3_4
XFILLER_117_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16512__A _16512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10182_ _19752_/Q _19751_/Q _19753_/Q _19750_/Q _19754_/Q vssd1 vssd1 vccd1 vccd1
+ _10759_/C sky130_fd_sc_hd__a41o_1
XFILLER_121_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14990_ _14990_/A _15094_/B _15009_/C vssd1 vssd1 vccd1 vccd1 _14993_/A sky130_fd_sc_hd__or3_4
XANTENNA__09126__A _17605_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13941_ _13941_/A vssd1 vssd1 vccd1 vccd1 _13941_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_247_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16660_ _16974_/X _16633_/X _16999_/X _16634_/X vssd1 vssd1 vccd1 vccd1 _16660_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_219_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13872_ _19199_/Q vssd1 vssd1 vccd1 vccd1 _13872_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17873__S0 _17913_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_216_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15611_ _18597_/Q vssd1 vssd1 vccd1 vccd1 _15611_/Y sky130_fd_sc_hd__inv_2
X_12823_ _18812_/Q vssd1 vssd1 vccd1 vccd1 _13536_/A sky130_fd_sc_hd__clkinv_1
XANTENNA__19745__RESET_B repeater205/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16591_ _16688_/A vssd1 vssd1 vccd1 vccd1 _16591_/X sky130_fd_sc_hd__buf_4
XFILLER_222_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12487__A _12659_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10078__B1 _10026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18330_ _18333_/CLK _18330_/D vssd1 vssd1 vccd1 vccd1 _18330_/Q sky130_fd_sc_hd__dfxtp_1
X_15542_ _19399_/Q vssd1 vssd1 vccd1 vccd1 _15542_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_188_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12754_ _19256_/Q vssd1 vssd1 vccd1 vccd1 _16719_/A sky130_fd_sc_hd__inv_2
XPHY_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10719__B _13252_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17489__S _17546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11705_ _11703_/A _18621_/Q hold210/X _10950_/A vssd1 vssd1 vccd1 vccd1 hold213/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_70_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18261_ _20076_/CLK _18261_/D vssd1 vssd1 vccd1 vccd1 _18261_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12685_ _12699_/A vssd1 vssd1 vccd1 vccd1 _12685_/X sky130_fd_sc_hd__clkbuf_2
X_15473_ _18563_/Q vssd1 vssd1 vccd1 vccd1 _15475_/A sky130_fd_sc_hd__inv_2
XFILLER_203_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17212_ _17473_/A0 _09880_/Y _17522_/S vssd1 vssd1 vccd1 vccd1 _17212_/X sky130_fd_sc_hd__mux2_1
XPHY_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14424_ _14425_/A vssd1 vssd1 vccd1 vccd1 _14424_/X sky130_fd_sc_hd__clkbuf_2
X_11636_ _19551_/Q _11635_/Y _11622_/B _11563_/X vssd1 vssd1 vccd1 vccd1 _19551_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__14764__B1 _14751_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18192_ _18216_/CLK _18192_/D vssd1 vssd1 vccd1 vccd1 _18192_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17143_ _17142_/X _11418_/Y _17548_/S vssd1 vssd1 vccd1 vccd1 _17143_/X sky130_fd_sc_hd__mux2_1
XPHY_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_repeater240_A repeater241/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11567_ _11567_/A vssd1 vssd1 vccd1 vccd1 _11590_/B sky130_fd_sc_hd__inv_2
XFILLER_11_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14355_ hold237/X vssd1 vssd1 vccd1 vccd1 _14749_/A sky130_fd_sc_hd__clkbuf_2
XPHY_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10518_ _19544_/Q vssd1 vssd1 vccd1 vccd1 _10530_/A sky130_fd_sc_hd__inv_2
X_13306_ _18859_/Q vssd1 vssd1 vccd1 vccd1 _13431_/D sky130_fd_sc_hd__clkinv_2
XANTENNA__14516__B1 _14474_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17074_ _17073_/X _18824_/Q _17386_/S vssd1 vssd1 vccd1 vccd1 _17074_/X sky130_fd_sc_hd__mux2_2
XFILLER_155_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14286_ _18754_/Q _14286_/B _15192_/A vssd1 vssd1 vccd1 vccd1 _15082_/C sky130_fd_sc_hd__or3_4
XFILLER_170_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11498_ _19605_/Q _11497_/Y _11490_/X _11486_/B vssd1 vssd1 vccd1 vccd1 _19605_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__18698__RESET_B hold359/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13237_ _18881_/Q _13231_/A _18543_/Q _13230_/A vssd1 vssd1 vccd1 vccd1 _18881_/D
+ sky130_fd_sc_hd__a22o_1
X_16025_ _18244_/Q _16096_/B vssd1 vssd1 vccd1 vccd1 _16025_/Y sky130_fd_sc_hd__nor2_1
XFILLER_226_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10449_ _19832_/Q _10441_/X _10448_/X _10442_/X vssd1 vssd1 vccd1 vccd1 _19832_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18627__RESET_B repeater221/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13168_ _13087_/A _13168_/A2 _13166_/Y _13199_/B vssd1 vssd1 vccd1 vccd1 _18915_/D
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__11566__A _19024_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12119_ _19302_/Q _12114_/X _11911_/X _12115_/X vssd1 vssd1 vccd1 vccd1 _19302_/D
+ sky130_fd_sc_hd__a22o_1
X_17976_ _20090_/CLK _17976_/D vssd1 vssd1 vccd1 vccd1 _17976_/Q sky130_fd_sc_hd__dfxtp_1
X_13099_ _19177_/Q _13078_/A _16544_/A _18901_/Q vssd1 vssd1 vccd1 vccd1 _13099_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_242_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19715_ _19795_/CLK _19715_/D repeater218/X vssd1 vssd1 vccd1 vccd1 _19715_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_78_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16927_ _19471_/Q hold193/X _16950_/S vssd1 vssd1 vccd1 vccd1 _16927_/X sky130_fd_sc_hd__mux2_1
XFILLER_66_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_81_HCLK clkbuf_4_13_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19283_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_226_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19646_ _19859_/CLK _19646_/D repeater262/X vssd1 vssd1 vccd1 vccd1 _19646_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_65_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16858_ _16857_/X _09401_/Y _17529_/S vssd1 vssd1 vccd1 vccd1 _16858_/X sky130_fd_sc_hd__mux2_1
XANTENNA__17864__S0 _19633_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14047__A2 _18701_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_214_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19486__RESET_B repeater260/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15809_ _18218_/Q vssd1 vssd1 vccd1 vccd1 _15809_/Y sky130_fd_sc_hd__inv_2
X_19577_ _19577_/CLK _19577_/D repeater268/X vssd1 vssd1 vccd1 vccd1 _19577_/Q sky130_fd_sc_hd__dfrtp_1
X_16789_ _16716_/Y _18989_/Q _17459_/S vssd1 vssd1 vccd1 vccd1 _16789_/X sky130_fd_sc_hd__mux2_1
XFILLER_46_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09330_ _20046_/Q _15724_/A _20046_/Q _15724_/A vssd1 vssd1 vccd1 vccd1 _09330_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_18528_ _19771_/CLK _18528_/D repeater189/X vssd1 vssd1 vccd1 vccd1 _18528_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__19415__RESET_B repeater193/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17399__S _17568_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09261_ _12257_/A _15914_/A vssd1 vssd1 vccd1 vccd1 _09340_/B sky130_fd_sc_hd__or2_2
XFILLER_179_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18459_ _18869_/CLK _18459_/D vssd1 vssd1 vccd1 vccd1 _18459_/Q sky130_fd_sc_hd__dfxtp_1
X_09192_ _09192_/A _09192_/B vssd1 vssd1 vccd1 vccd1 _09192_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__15858__D _15858_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17919__S1 _18752_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12230__A1 _19233_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14507__B1 _14441_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13021__A _13021_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15180__B1 _09255_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20023__CLK _20091_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11741__B1 _16930_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18070__CLK _18169_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08976_ _20069_/Q vssd1 vssd1 vccd1 vccd1 _08977_/C sky130_fd_sc_hd__inv_2
XFILLER_248_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17855__S0 _17908_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold166_A HADDR[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13246__B1 _12602_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09528_ _09516_/X _09528_/B _09528_/C _09528_/D vssd1 vssd1 vccd1 vccd1 _09565_/B
+ sky130_fd_sc_hd__and4b_1
XPHY_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold333_A HWDATA[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12100__A hold318/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09459_ _19929_/Q vssd1 vssd1 vccd1 vccd1 _10045_/A sky130_fd_sc_hd__inv_2
XPHY_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11272__A2 _19013_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15411__A _15413_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17102__S _17459_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12470_ _19105_/Q _12464_/X hold270/X _12465_/X vssd1 vssd1 vccd1 vccd1 _19105_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_131_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11421_ _11581_/A _19148_/Q _19547_/Q _11420_/Y vssd1 vssd1 vccd1 vccd1 _11421_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__16941__S _16946_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14140_ _18679_/Q _14139_/Y _14112_/A _14140_/C1 vssd1 vssd1 vccd1 vccd1 _18679_/D
+ sky130_fd_sc_hd__o211a_1
X_11352_ _19579_/Q _11351_/Y _19605_/Q _11300_/Y vssd1 vssd1 vccd1 vccd1 _11352_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_152_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18791__RESET_B repeater261/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11980__B1 _11978_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10303_ _18599_/Q _15617_/A vssd1 vssd1 vccd1 vccd1 _15621_/A sky130_fd_sc_hd__or2_2
XFILLER_180_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14071_ _14068_/Y _18677_/Q _19064_/Q _14006_/A _14070_/X vssd1 vssd1 vccd1 vccd1
+ _14080_/B sky130_fd_sc_hd__o221a_1
X_11283_ _19018_/Q vssd1 vssd1 vccd1 vccd1 _11283_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18720__RESET_B repeater253/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13022_ _12859_/B _13024_/A _12859_/A vssd1 vssd1 vccd1 vccd1 _13023_/B sky130_fd_sc_hd__o21a_1
X_10234_ _19839_/Q vssd1 vssd1 vccd1 vccd1 _10234_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11386__A _19147_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17830_ _18336_/Q _18216_/Q _18208_/Q _18200_/Q _17918_/S0 _18750_/Q vssd1 vssd1
+ vccd1 vccd1 _17830_/X sky130_fd_sc_hd__mux4_1
X_10165_ _19499_/Q _14245_/A _11842_/B _10186_/B vssd1 vssd1 vccd1 vccd1 _10174_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_86_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_158_HCLK_A clkbuf_4_0_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17761_ _15195_/Y _15194_/Y _17761_/S vssd1 vssd1 vccd1 vccd1 _17761_/X sky130_fd_sc_hd__mux2_2
X_10096_ _10084_/A _10084_/B _10094_/Y _10107_/C vssd1 vssd1 vccd1 vccd1 _19912_/D
+ sky130_fd_sc_hd__a211oi_2
X_14973_ _18067_/Q _14965_/A _14816_/X _14966_/A vssd1 vssd1 vccd1 vccd1 _18067_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_208_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19500_ _19859_/CLK hold222/X repeater262/X vssd1 vssd1 vccd1 vccd1 _19500_/Q sky130_fd_sc_hd__dfrtp_2
X_16712_ _16850_/X _16683_/X _16847_/X _16684_/X _16711_/X vssd1 vssd1 vccd1 vccd1
+ _16715_/B sky130_fd_sc_hd__o221a_4
XANTENNA__10838__A2 _10831_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13924_ _13924_/A vssd1 vssd1 vccd1 vccd1 _13924_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17846__S0 _17908_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17692_ _15464_/X _19443_/Q _17696_/S vssd1 vssd1 vccd1 vccd1 _18560_/D sky130_fd_sc_hd__mux2_1
XFILLER_47_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19431_ _20003_/CLK _19431_/D repeater185/X vssd1 vssd1 vccd1 vccd1 _19431_/Q sky130_fd_sc_hd__dfrtp_1
X_16643_ _16643_/A _16647_/B vssd1 vssd1 vccd1 vccd1 _16643_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__11833__B _12309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13855_ _19201_/Q vssd1 vssd1 vccd1 vccd1 _13855_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12806_ _19249_/Q _13549_/A _16646_/A _18826_/Q vssd1 vssd1 vccd1 vccd1 _12806_/X
+ sky130_fd_sc_hd__o22a_1
X_19362_ _19968_/CLK _19362_/D hold370/X vssd1 vssd1 vccd1 vccd1 _19362_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_16_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14985__B1 _14791_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16574_ _16684_/A vssd1 vssd1 vccd1 vccd1 _16574_/X sky130_fd_sc_hd__buf_2
XANTENNA__12010__A _12017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10998_ _10998_/A vssd1 vssd1 vccd1 vccd1 _19661_/D sky130_fd_sc_hd__inv_2
X_13786_ _18726_/Q vssd1 vssd1 vccd1 vccd1 _13912_/D sky130_fd_sc_hd__inv_4
XFILLER_222_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11799__B1 _09039_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18313_ _18416_/CLK _18313_/D vssd1 vssd1 vccd1 vccd1 _18313_/Q sky130_fd_sc_hd__dfxtp_1
X_15525_ _15530_/B vssd1 vssd1 vccd1 vccd1 _15525_/Y sky130_fd_sc_hd__inv_2
X_12737_ _19244_/Q vssd1 vssd1 vccd1 vccd1 _16586_/A sky130_fd_sc_hd__inv_2
XANTENNA__12460__A1 _19113_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19293_ _19293_/CLK _19293_/D repeater211/X vssd1 vssd1 vccd1 vccd1 _19293_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_148_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17012__S _17522_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18244_ _19847_/CLK _18244_/D vssd1 vssd1 vccd1 vccd1 _18244_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14737__B1 _14606_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_230_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15456_ _18559_/Q vssd1 vssd1 vccd1 vccd1 _15456_/Y sky130_fd_sc_hd__inv_2
XPHY_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12668_ _18988_/Q _12661_/X hold279/X _12664_/X vssd1 vssd1 vccd1 vccd1 _18988_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14407_ _19642_/Q _19641_/Q _15296_/B vssd1 vssd1 vccd1 vccd1 _14571_/C sky130_fd_sc_hd__or3_4
X_11619_ _11639_/A _11639_/B _11619_/C vssd1 vssd1 vccd1 vccd1 _11637_/A sky130_fd_sc_hd__or3_1
X_18175_ _18198_/CLK _18175_/D vssd1 vssd1 vccd1 vccd1 _18175_/Q sky130_fd_sc_hd__dfxtp_1
X_15387_ _15208_/Y _15386_/Y _15384_/A vssd1 vssd1 vccd1 vccd1 _18510_/D sky130_fd_sc_hd__o21a_1
XFILLER_191_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16851__S _17534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18808__RESET_B repeater217/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12599_ _14277_/A vssd1 vssd1 vccd1 vccd1 _12599_/X sky130_fd_sc_hd__buf_4
XFILLER_237_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17126_ _17125_/X _15624_/Y _17318_/S vssd1 vssd1 vccd1 vccd1 _17126_/X sky130_fd_sc_hd__mux2_2
X_14338_ _14338_/A vssd1 vssd1 vccd1 vccd1 _14338_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__11971__B1 _09071_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17057_ _17473_/A0 _16681_/Y _17547_/S vssd1 vssd1 vccd1 vccd1 _17057_/X sky130_fd_sc_hd__mux2_1
X_14269_ _18466_/Q _14259_/A _14268_/X _14260_/A vssd1 vssd1 vccd1 vccd1 _18466_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_98_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16008_ _18020_/Q vssd1 vssd1 vccd1 vccd1 _16008_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17682__S _17683_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17959_ _20079_/CLK _17959_/D vssd1 vssd1 vccd1 vccd1 _17959_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__19667__RESET_B repeater270/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_17_HCLK_A clkbuf_4_3_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17837__S0 _17908_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19629_ _19630_/CLK _19629_/D repeater257/X vssd1 vssd1 vccd1 vccd1 _19629_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_5_HCLK_A clkbuf_4_2_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09313_ _20047_/Q vssd1 vssd1 vccd1 vccd1 _09313_/Y sky130_fd_sc_hd__inv_2
XFILLER_222_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17914__A0 _17910_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09244_ _19872_/Q _10181_/A _19877_/Q _19750_/Q vssd1 vssd1 vccd1 vccd1 _09253_/S
+ sky130_fd_sc_hd__or4_4
XFILLER_166_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12203__A1 _19250_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09175_ _14707_/A _09163_/X _09174_/X _09165_/X vssd1 vssd1 vccd1 vccd1 _20078_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_147_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09080__B1 _09079_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12590__A _12598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11714__B1 _16949_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17592__S _17600_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_hold283_A HWDATA[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08959_ _18776_/Q vssd1 vssd1 vccd1 vccd1 _08959_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17828__S0 _17918_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11970_ _11979_/A vssd1 vssd1 vccd1 vccd1 _11970_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_56_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19981__CLK _19992_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10921_ _19681_/Q _18511_/Q _10920_/Y _10912_/C vssd1 vssd1 vccd1 vccd1 _10922_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_205_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16936__S _16946_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10852_ _19710_/Q _10844_/A _10425_/X _10845_/A vssd1 vssd1 vccd1 vccd1 _19710_/D
+ sky130_fd_sc_hd__a22o_1
X_13640_ _13637_/A _13630_/X _13637_/Y vssd1 vssd1 vccd1 vccd1 _18796_/D sky130_fd_sc_hd__a21oi_1
XANTENNA__14967__B1 _14802_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09438__A2 _09436_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13571_ _13588_/A vssd1 vssd1 vccd1 vccd1 _13571_/X sky130_fd_sc_hd__clkbuf_4
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10783_ _20036_/Q vssd1 vssd1 vccd1 vccd1 _10805_/A sky130_fd_sc_hd__inv_2
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16237__A _17386_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15310_ _15309_/Y _15307_/X _15268_/X vssd1 vssd1 vccd1 vccd1 _18628_/D sky130_fd_sc_hd__o21ai_1
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10453__B1 _10451_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12522_ _19071_/Q _12519_/X _12356_/X _12520_/X vssd1 vssd1 vccd1 vccd1 _19071_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16290_ _18111_/Q vssd1 vssd1 vccd1 vccd1 _16290_/Y sky130_fd_sc_hd__inv_2
XFILLER_197_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20069__CLK _20070_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17381__A1 _19405_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15241_ _15259_/A vssd1 vssd1 vccd1 vccd1 _15285_/A sky130_fd_sc_hd__buf_1
X_12453_ _19118_/Q _12450_/X _12392_/X _12451_/X vssd1 vssd1 vccd1 vccd1 _19118_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_184_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18901__RESET_B repeater188/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11404_ _11575_/A _19142_/Q _11580_/A _19147_/Q vssd1 vssd1 vccd1 vccd1 _11404_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08949__B2 _08945_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12384_ hold279/X vssd1 vssd1 vccd1 vccd1 _12384_/X sky130_fd_sc_hd__buf_2
X_15172_ _15172_/A vssd1 vssd1 vccd1 vccd1 _15172_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_181_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11953__B1 _09037_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11335_ _11473_/A _18975_/Q _19593_/Q _11334_/Y vssd1 vssd1 vccd1 vccd1 _11335_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_21_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14123_ _14123_/A vssd1 vssd1 vccd1 vccd1 _14123_/Y sky130_fd_sc_hd__clkinv_1
XANTENNA__15144__B1 _09255_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19980_ _19992_/CLK _19980_/D repeater192/X vssd1 vssd1 vccd1 vccd1 _19980_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_180_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16892__A0 _17486_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18931_ _19282_/CLK _18931_/D repeater215/X vssd1 vssd1 vccd1 vccd1 _18931_/Q sky130_fd_sc_hd__dfrtp_1
X_14054_ _19074_/Q vssd1 vssd1 vccd1 vccd1 _14054_/Y sky130_fd_sc_hd__inv_2
X_11266_ _19584_/Q _11264_/Y _11463_/A _18996_/Q vssd1 vssd1 vccd1 vccd1 _11266_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_180_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11705__B1 hold210/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10217_ _19666_/Q vssd1 vssd1 vccd1 vccd1 _10966_/A sky130_fd_sc_hd__inv_2
X_13005_ _13005_/A _13014_/A vssd1 vssd1 vccd1 vccd1 _13006_/B sky130_fd_sc_hd__or2_2
X_18862_ _18866_/CLK _18862_/D repeater232/X vssd1 vssd1 vccd1 vccd1 _18862_/Q sky130_fd_sc_hd__dfrtp_1
X_11197_ _17719_/X _11191_/X _19612_/Q _11192_/X vssd1 vssd1 vccd1 vccd1 _19612_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_repeater203_A repeater204/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17813_ _17930_/Q _18452_/Q _18460_/Q _18060_/Q _17918_/S0 _18750_/Q vssd1 vssd1
+ vccd1 vccd1 _17813_/X sky130_fd_sc_hd__mux4_2
X_10148_ _10148_/A _19515_/Q _10250_/C vssd1 vssd1 vccd1 vccd1 _12370_/C sky130_fd_sc_hd__or3_4
XFILLER_94_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18793_ _18795_/CLK _18793_/D repeater261/X vssd1 vssd1 vccd1 vccd1 _18793_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_223_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17007__S _17547_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11844__A _15867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17744_ _15365_/Y _19701_/Q _18508_/D vssd1 vssd1 vccd1 vccd1 _17744_/X sky130_fd_sc_hd__mux2_1
XANTENNA__17819__S0 _18751_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10079_ _10079_/A vssd1 vssd1 vccd1 vccd1 _10107_/C sky130_fd_sc_hd__buf_2
X_14956_ _18080_/Q _14952_/X _14925_/X _14954_/X vssd1 vssd1 vccd1 vccd1 _18080_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_35_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19007__RESET_B hold346/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13907_ _13925_/A vssd1 vssd1 vccd1 vccd1 _13907_/X sky130_fd_sc_hd__clkbuf_2
X_17675_ _15535_/Y _19460_/Q _17683_/S vssd1 vssd1 vccd1 vccd1 _18577_/D sky130_fd_sc_hd__mux2_1
X_14887_ _18120_/Q _14883_/X _14806_/X _14885_/X vssd1 vssd1 vccd1 vccd1 _18120_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16846__S _17487_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19414_ _19905_/CLK _19414_/D repeater210/X vssd1 vssd1 vccd1 vccd1 _19414_/Q sky130_fd_sc_hd__dfrtp_1
X_16626_ _17068_/X _16555_/X _17065_/X _16556_/X vssd1 vssd1 vccd1 vccd1 _16629_/B
+ sky130_fd_sc_hd__a22o_1
X_13838_ _19219_/Q vssd1 vssd1 vccd1 vccd1 _13838_/Y sky130_fd_sc_hd__inv_2
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_111_HCLK clkbuf_opt_0_HCLK/A vssd1 vssd1 vccd1 vccd1 _18686_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_50_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19345_ _19952_/CLK _19345_/D repeater245/X vssd1 vssd1 vccd1 vccd1 _19345_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_16_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12433__A1 _19128_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16557_ _17118_/X _16597_/A _17108_/X _16598_/A vssd1 vssd1 vccd1 vccd1 _16557_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_15_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13769_ _18742_/Q _18743_/Q _13772_/S vssd1 vssd1 vccd1 vccd1 _18743_/D sky130_fd_sc_hd__mux2_1
XFILLER_204_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15508_ _18572_/Q vssd1 vssd1 vccd1 vccd1 _15511_/A sky130_fd_sc_hd__inv_2
XANTENNA__10444__B1 _09077_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19276_ _19282_/CLK _19276_/D repeater216/X vssd1 vssd1 vccd1 vccd1 _19276_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_176_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16488_ _17568_/S _17567_/S vssd1 vssd1 vccd1 vccd1 _16504_/A sky130_fd_sc_hd__or2_4
XFILLER_31_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18227_ _18412_/CLK _18227_/D vssd1 vssd1 vccd1 vccd1 _18227_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17677__S _17683_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15439_ _15439_/A _17569_/X vssd1 vssd1 vccd1 vccd1 _18550_/D sky130_fd_sc_hd__and2_1
XANTENNA__16580__C1 _16579_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12197__B1 _12080_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18158_ _18198_/CLK _18158_/D vssd1 vssd1 vccd1 vccd1 _18158_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09062__B1 _09061_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11944__B1 _09021_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold303 input56/X vssd1 vssd1 vccd1 vccd1 hold303/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold314 hold314/A vssd1 vssd1 vccd1 vccd1 hold314/X sky130_fd_sc_hd__dlygate4sd3_1
X_17109_ _17486_/A0 _13153_/Y _17543_/S vssd1 vssd1 vccd1 vccd1 _17109_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold325 hold325/A vssd1 vssd1 vccd1 vccd1 hold325/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18089_ _20079_/CLK _18089_/D vssd1 vssd1 vccd1 vccd1 _18089_/Q sky130_fd_sc_hd__dfxtp_1
Xhold336 input49/X vssd1 vssd1 vccd1 vccd1 hold336/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold347 hold364/X vssd1 vssd1 vccd1 vccd1 hold363/A sky130_fd_sc_hd__dlygate4sd3_1
X_20120_ _20120_/CLK _20120_/D repeater234/X vssd1 vssd1 vccd1 vccd1 _20120_/Q sky130_fd_sc_hd__dfrtp_4
Xhold358 hold358/A vssd1 vssd1 vccd1 vccd1 hold358/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold369 scl_i_S4 vssd1 vssd1 vccd1 vccd1 hold369/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09931_ _19351_/Q vssd1 vssd1 vccd1 vccd1 _16621_/A sky130_fd_sc_hd__inv_2
XANTENNA__19848__RESET_B repeater257/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20051_ _20051_/CLK _20051_/D repeater206/X vssd1 vssd1 vccd1 vccd1 _20051_/Q sky130_fd_sc_hd__dfrtp_1
X_09862_ _09862_/A _09978_/A vssd1 vssd1 vccd1 vccd1 _09863_/B sky130_fd_sc_hd__or2_2
XFILLER_140_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09793_ _09793_/A _09797_/A vssd1 vssd1 vccd1 vccd1 _09794_/B sky130_fd_sc_hd__or2_2
XFILLER_133_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_141_HCLK_A clkbuf_4_3_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater153 _17529_/S vssd1 vssd1 vccd1 vccd1 _17385_/S sky130_fd_sc_hd__buf_6
Xrepeater164 _17042_/S vssd1 vssd1 vccd1 vccd1 _17473_/S sky130_fd_sc_hd__buf_6
XFILLER_85_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater175 _17513_/S vssd1 vssd1 vccd1 vccd1 _17474_/S sky130_fd_sc_hd__buf_8
XPHY_4307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater186 repeater188/X vssd1 vssd1 vccd1 vccd1 repeater186/X sky130_fd_sc_hd__clkbuf_8
XPHY_4318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater197 repeater199/X vssd1 vssd1 vccd1 vccd1 repeater197/X sky130_fd_sc_hd__buf_6
XPHY_4329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12672__A1 _18986_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_213_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_210_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17587__S _17600_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09227_ _18644_/Q _09226_/X _18646_/Q vssd1 vssd1 vccd1 vccd1 _09227_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_139_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16571__C1 _16504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09158_ _20083_/Q _09156_/Y _09156_/B _09157_/X vssd1 vssd1 vccd1 vccd1 _20083_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_181_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09089_ hold245/X vssd1 vssd1 vccd1 vccd1 _10451_/A sky130_fd_sc_hd__buf_4
X_11120_ _17755_/X _11108_/Y _11119_/X _11094_/Y _19636_/Q vssd1 vssd1 vccd1 vccd1
+ _19636_/D sky130_fd_sc_hd__a32o_1
XFILLER_162_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13688__B1 _13676_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11051_ _19643_/Q vssd1 vssd1 vccd1 vccd1 _11147_/A sky130_fd_sc_hd__inv_2
XFILLER_107_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12360__B1 _12296_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10002_ _19940_/Q _10001_/Y _10002_/B1 _09964_/X vssd1 vssd1 vccd1 vccd1 _19940_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_77_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_237_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18486__SET_B repeater222/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14810_ _14810_/A vssd1 vssd1 vccd1 vccd1 _14810_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__19171__RESET_B hold370/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15790_ _18162_/Q vssd1 vssd1 vccd1 vccd1 _15790_/Y sky130_fd_sc_hd__inv_2
XFILLER_92_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12112__B1 _12030_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_217_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_134_HCLK clkbuf_4_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19462_/CLK sky130_fd_sc_hd__clkbuf_16
X_14741_ _18203_/Q _14733_/A _14691_/X _14734_/A vssd1 vssd1 vccd1 vccd1 _18203_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_91_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11953_ _19389_/Q _11948_/X _09037_/X _11949_/X vssd1 vssd1 vccd1 vccd1 _19389_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16929__A1 hold199/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_63_HCLK_A clkbuf_opt_3_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20076__RESET_B repeater196/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10904_ _18481_/Q vssd1 vssd1 vccd1 vccd1 _15208_/B sky130_fd_sc_hd__inv_2
X_17460_ _17459_/X _11444_/Y _17548_/S vssd1 vssd1 vccd1 vccd1 _17460_/X sky130_fd_sc_hd__mux2_1
XFILLER_233_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14672_ _18241_/Q _14669_/X _09168_/X _14671_/X vssd1 vssd1 vccd1 vccd1 _18241_/D
+ sky130_fd_sc_hd__a22o_1
X_11884_ _11891_/A vssd1 vssd1 vccd1 vccd1 _11884_/X sky130_fd_sc_hd__buf_1
XFILLER_45_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14404__A2 _14395_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16411_ _18409_/Q vssd1 vssd1 vccd1 vccd1 _16411_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13623_ _13499_/X _13617_/Y _17762_/S _13621_/X _13622_/X vssd1 vssd1 vccd1 vccd1
+ _13623_/X sky130_fd_sc_hd__o221a_1
X_10835_ _15349_/A _10831_/B _10834_/Y _10708_/Y _10840_/S vssd1 vssd1 vccd1 vccd1
+ _10836_/A sky130_fd_sc_hd__o32a_1
X_17391_ _16208_/Y _18964_/Q _17459_/S vssd1 vssd1 vccd1 vccd1 _17391_/X sky130_fd_sc_hd__mux2_1
XFILLER_198_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10426__B1 _10425_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19130_ _19970_/CLK _19130_/D repeater249/X vssd1 vssd1 vccd1 vccd1 _19130_/Q sky130_fd_sc_hd__dfrtp_2
X_16342_ _18472_/Q vssd1 vssd1 vccd1 vccd1 _16342_/Y sky130_fd_sc_hd__inv_2
XFILLER_186_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13554_ _13554_/A _13566_/A vssd1 vssd1 vccd1 vccd1 _13555_/B sky130_fd_sc_hd__or2_2
XFILLER_13_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10766_ _19750_/Q _10766_/B vssd1 vssd1 vccd1 vccd1 _10767_/B sky130_fd_sc_hd__and2_1
XANTENNA__09292__B1 _09090_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19061_ _19610_/CLK _19061_/D hold343/X vssd1 vssd1 vccd1 vccd1 _19061_/Q sky130_fd_sc_hd__dfrtp_1
X_12505_ _12505_/A vssd1 vssd1 vccd1 vccd1 _12505_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__17497__S _19498_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16273_ _16434_/B vssd1 vssd1 vccd1 vccd1 _16415_/B sky130_fd_sc_hd__buf_1
XANTENNA__18751__CLK _19900_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13485_ _13485_/A _13485_/B _13489_/C vssd1 vssd1 vccd1 vccd1 _18840_/D sky130_fd_sc_hd__nor3_1
X_10697_ _10451_/A _17749_/X _17749_/S _10694_/Y _19778_/Q vssd1 vssd1 vccd1 vccd1
+ _19778_/D sky130_fd_sc_hd__a32o_1
XANTENNA_repeater153_A _17529_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12179__B1 _11926_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18012_ _18954_/CLK _18012_/D vssd1 vssd1 vccd1 vccd1 _18012_/Q sky130_fd_sc_hd__dfxtp_1
X_15224_ _15224_/A vssd1 vssd1 vccd1 vccd1 _15334_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__09044__B1 hold314/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12436_ _15867_/A _15858_/C _12436_/C _19500_/Q vssd1 vssd1 vccd1 vccd1 _15863_/B
+ sky130_fd_sc_hd__or4b_4
XFILLER_154_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11839__A _12558_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15155_ _17954_/Q _15147_/A _14713_/A _15148_/A vssd1 vssd1 vccd1 vccd1 _17954_/D
+ sky130_fd_sc_hd__a22o_1
X_12367_ _19160_/Q _12361_/X _12236_/X _12362_/X vssd1 vssd1 vccd1 vccd1 _19160_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_154_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output82_A _16533_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14106_ _14118_/A vssd1 vssd1 vccd1 vccd1 _14106_/X sky130_fd_sc_hd__clkbuf_4
X_11318_ _19591_/Q _18973_/Q _11471_/A _11317_/Y vssd1 vssd1 vccd1 vccd1 _11318_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_126_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15086_ _18001_/Q _15083_/X hold247/X _15085_/X vssd1 vssd1 vccd1 vccd1 _18001_/D
+ sky130_fd_sc_hd__a22o_1
X_12298_ _12298_/A vssd1 vssd1 vccd1 vccd1 _12298_/X sky130_fd_sc_hd__clkbuf_2
X_19963_ _19968_/CLK _19963_/D hold370/X vssd1 vssd1 vccd1 vccd1 _19963_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_113_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13679__B1 _13678_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11249_ _19594_/Q vssd1 vssd1 vccd1 vccd1 _11474_/A sky130_fd_sc_hd__inv_2
X_14037_ _19092_/Q _14034_/Y _14035_/Y _18681_/Q _14036_/X vssd1 vssd1 vccd1 vccd1
+ _14049_/A sky130_fd_sc_hd__a221o_1
X_18914_ _19222_/CLK _18914_/D repeater188/X vssd1 vssd1 vccd1 vccd1 _18914_/Q sky130_fd_sc_hd__dfrtp_1
X_19894_ _20055_/CLK _19894_/D repeater205/X vssd1 vssd1 vccd1 vccd1 _19894_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12351__B1 hold270/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18845_ _18866_/CLK _18845_/D repeater233/X vssd1 vssd1 vccd1 vccd1 _18845_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_79_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18131__CLK _18198_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_227_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18776_ _19855_/CLK _18776_/D repeater264/X vssd1 vssd1 vccd1 vccd1 _18776_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_67_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13492__C _15190_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15988_ _15983_/Y _15836_/A _15984_/Y _15838_/X _15987_/X vssd1 vssd1 vccd1 vccd1
+ _15988_/X sky130_fd_sc_hd__o221a_1
XANTENNA__12103__B1 _12102_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17727_ _19673_/Q _19686_/Q _18510_/Q vssd1 vssd1 vccd1 vccd1 _17727_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14939_ _14940_/A vssd1 vssd1 vccd1 vccd1 _14939_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__17042__A0 _17473_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18281__CLK _19847_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17658_ _15603_/X _19031_/Q _17664_/S vssd1 vssd1 vccd1 vccd1 _18594_/D sky130_fd_sc_hd__mux2_1
X_16609_ _19044_/Q vssd1 vssd1 vccd1 vccd1 _16609_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18507__D _18507_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17589_ _15359_/X _19714_/Q _17600_/S vssd1 vssd1 vccd1 vccd1 _17589_/X sky130_fd_sc_hd__mux2_1
XANTENNA__18823__RESET_B repeater217/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19328_ _19971_/CLK _19328_/D repeater241/X vssd1 vssd1 vccd1 vccd1 _19328_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_204_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17345__A1 _19832_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19259_ _20035_/CLK _19259_/D repeater242/X vssd1 vssd1 vccd1 vccd1 _19259_/Q sky130_fd_sc_hd__dfrtp_1
X_09012_ _10842_/A _11996_/A vssd1 vssd1 vccd1 vccd1 _12659_/A sky130_fd_sc_hd__or2_4
XANTENNA__17200__S _17534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_15_HCLK clkbuf_4_2_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _18216_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__11917__B1 _10885_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold133 input10/X vssd1 vssd1 vccd1 vccd1 hold133/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 hold144/A vssd1 vssd1 vccd1 vccd1 hold144/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__19682__RESET_B repeater219/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold155 hold155/A vssd1 vssd1 vccd1 vccd1 hold155/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold166 HADDR[13] vssd1 vssd1 vccd1 vccd1 input5/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 input32/X vssd1 vssd1 vccd1 vccd1 hold177/X sky130_fd_sc_hd__dlygate4sd3_1
X_20103_ _20107_/CLK _20103_/D repeater233/X vssd1 vssd1 vccd1 vccd1 _20103_/Q sky130_fd_sc_hd__dfrtp_2
Xhold188 hold188/A vssd1 vssd1 vccd1 vccd1 hold188/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold199 input23/X vssd1 vssd1 vccd1 vccd1 hold199/X sky130_fd_sc_hd__dlygate4sd3_1
X_09914_ _19346_/Q vssd1 vssd1 vccd1 vccd1 _09914_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20034_ _20035_/CLK _20034_/D repeater240/X vssd1 vssd1 vccd1 vccd1 _20034_/Q sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_157_HCLK clkbuf_4_0_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19637_/CLK sky130_fd_sc_hd__clkbuf_16
X_09845_ _19941_/Q vssd1 vssd1 vccd1 vccd1 _09850_/A sky130_fd_sc_hd__inv_2
XFILLER_247_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09776_ _19991_/Q _09775_/Y _09763_/X _09748_/B vssd1 vssd1 vccd1 vccd1 _19991_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_160_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12645__A1 _19003_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14795__A hold264/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17033__A0 _17486_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold246_A HWDATA[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_214_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10620_ _10620_/A vssd1 vssd1 vccd1 vccd1 _19810_/D sky130_fd_sc_hd__inv_2
XFILLER_168_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09274__B1 _09090_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10551_ _10551_/A vssd1 vssd1 vccd1 vccd1 _10552_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_195_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17110__S _17487_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10482_ _19545_/Q vssd1 vssd1 vccd1 vccd1 _10734_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__09026__B1 _09025_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13270_ _18755_/Q vssd1 vssd1 vccd1 vccd1 _14366_/B sky130_fd_sc_hd__buf_1
XFILLER_211_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11908__B1 _09075_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12221_ _19238_/Q _12219_/X _12035_/X _12220_/X vssd1 vssd1 vccd1 vccd1 _19238_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_136_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12581__B1 _12408_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12152_ _19283_/Q _12150_/X _12095_/X _12151_/X vssd1 vssd1 vccd1 vccd1 _19283_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18154__CLK _19900_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11103_ _11103_/A _11103_/B _11103_/C _11103_/D vssd1 vssd1 vccd1 vccd1 _11103_/X
+ sky130_fd_sc_hd__or4_4
XANTENNA_clkbuf_2_2_0_HCLK_A clkbuf_2_3_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16960_ _15963_/X _12798_/Y _17534_/S vssd1 vssd1 vccd1 vccd1 _16960_/X sky130_fd_sc_hd__mux2_1
X_12083_ hold303/X vssd1 vssd1 vccd1 vccd1 _12083_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_2_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12333__B1 _12092_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11034_ _11031_/X _11030_/X _11031_/X _11030_/X vssd1 vssd1 vccd1 vccd1 _19651_/D
+ sky130_fd_sc_hd__o2bb2ai_1
X_15911_ _15911_/A vssd1 vssd1 vccd1 vccd1 _16509_/A sky130_fd_sc_hd__clkbuf_2
X_16891_ _16890_/X _13840_/Y _17545_/S vssd1 vssd1 vccd1 vccd1 _16891_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18630_ _18633_/CLK _18630_/D repeater225/X vssd1 vssd1 vccd1 vccd1 _18630_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__16075__B2 _16003_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15842_ _16055_/A vssd1 vssd1 vccd1 vccd1 _15842_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_92_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18561_ _19992_/CLK _18561_/D repeater198/X vssd1 vssd1 vccd1 vccd1 _18561_/Q sky130_fd_sc_hd__dfrtp_1
X_15773_ _16723_/B vssd1 vssd1 vccd1 vccd1 _17042_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA_output120_A _16751_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12985_ _12985_/A vssd1 vssd1 vccd1 vccd1 _12986_/A sky130_fd_sc_hd__buf_6
X_17512_ _17511_/X _15879_/Y _17512_/S vssd1 vssd1 vccd1 vccd1 _17512_/X sky130_fd_sc_hd__mux2_1
XFILLER_205_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14724_ _18214_/Q _14717_/X _14723_/X _14719_/X vssd1 vssd1 vccd1 vccd1 _18214_/D
+ sky130_fd_sc_hd__a22o_1
X_18492_ _20057_/CLK _18492_/D repeater202/X vssd1 vssd1 vccd1 vccd1 _18492_/Q sky130_fd_sc_hd__dfrtp_1
X_11936_ _11936_/A _15897_/A vssd1 vssd1 vccd1 vccd1 _12066_/A sky130_fd_sc_hd__or2_2
XFILLER_18_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17443_ _17486_/A0 _09896_/Y _17543_/S vssd1 vssd1 vccd1 vccd1 _17443_/X sky130_fd_sc_hd__mux2_1
X_14655_ _14681_/A _16115_/A vssd1 vssd1 vccd1 vccd1 _14657_/A sky130_fd_sc_hd__or2_4
XANTENNA_repeater270_A repeater272/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11867_ _11867_/A _11869_/B vssd1 vssd1 vccd1 vccd1 _11867_/X sky130_fd_sc_hd__or2_1
XFILLER_14_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13606_ _13532_/A _13606_/A2 _13588_/X _13604_/Y vssd1 vssd1 vccd1 vccd1 _18808_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_177_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09265__A0 _09255_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17374_ _16295_/X _17966_/Q _17564_/S vssd1 vssd1 vccd1 vccd1 _17374_/X sky130_fd_sc_hd__mux2_1
X_10818_ _20036_/Q _10788_/Y _20050_/Q _19725_/Q _10810_/X vssd1 vssd1 vccd1 vccd1
+ _19725_/D sky130_fd_sc_hd__a32o_1
XPHY_3992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14586_ _14598_/A _14598_/B _15070_/C vssd1 vssd1 vccd1 vccd1 _14588_/A sky130_fd_sc_hd__or3_4
X_11798_ _19462_/Q _11793_/X _09037_/X _11794_/X vssd1 vssd1 vccd1 vccd1 _19462_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_201_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19113_ _19115_/CLK _19113_/D hold353/X vssd1 vssd1 vccd1 vccd1 _19113_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_119_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16325_ _17350_/X _16148_/X _17359_/X _16003_/X vssd1 vssd1 vccd1 vccd1 _16325_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_229_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13537_ _13537_/A _13537_/B _13537_/C vssd1 vssd1 vccd1 vccd1 _13538_/B sky130_fd_sc_hd__or3_1
X_10749_ _19758_/Q _10742_/A _10423_/X _10743_/A vssd1 vssd1 vccd1 vccd1 _19758_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17020__S _17413_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19044_ _19597_/CLK _19044_/D repeater255/X vssd1 vssd1 vccd1 vccd1 _19044_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_118_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16256_ _17991_/Q vssd1 vssd1 vccd1 vccd1 _16256_/Y sky130_fd_sc_hd__inv_2
X_13468_ _13468_/A _13468_/B vssd1 vssd1 vccd1 vccd1 _13473_/A sky130_fd_sc_hd__or2_1
XFILLER_173_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15207_ _18640_/Q vssd1 vssd1 vccd1 vccd1 _15208_/A sky130_fd_sc_hd__inv_2
XFILLER_127_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12419_ _19138_/Q _12412_/X hold270/X _12414_/X vssd1 vssd1 vccd1 vccd1 _19138_/D
+ sky130_fd_sc_hd__a22o_1
X_16187_ _18262_/Q vssd1 vssd1 vccd1 vccd1 _16187_/Y sky130_fd_sc_hd__inv_2
X_13399_ _20121_/Q vssd1 vssd1 vccd1 vccd1 _13399_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16838__A0 _17473_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12572__B1 _12392_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09039__A hold298/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15138_ _17967_/Q _15134_/X hold236/X _15136_/X vssd1 vssd1 vccd1 vccd1 _17967_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_142_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15069_ _18010_/Q _15060_/A _15020_/X _15061_/A vssd1 vssd1 vccd1 vccd1 _18010_/D
+ sky130_fd_sc_hd__a22o_1
X_19946_ _19976_/CLK _19946_/D repeater244/X vssd1 vssd1 vccd1 vccd1 _19946_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_229_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12324__B1 _12076_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19877_ _20050_/CLK _19877_/D repeater197/X vssd1 vssd1 vccd1 vccd1 _19877_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_68_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17690__S _17696_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10886__B1 _10885_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09630_ _20001_/Q vssd1 vssd1 vccd1 vccd1 _09667_/C sky130_fd_sc_hd__inv_2
X_18828_ _19255_/CLK _18828_/D repeater239/X vssd1 vssd1 vccd1 vccd1 _18828_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_56_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09561_ _19318_/Q vssd1 vssd1 vccd1 vccd1 _16670_/A sky130_fd_sc_hd__inv_2
XFILLER_67_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18759_ _20123_/CLK _18759_/D repeater195/X vssd1 vssd1 vccd1 vccd1 _18759_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__17015__A0 _15768_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09492_ _09492_/A _09492_/B vssd1 vssd1 vccd1 vccd1 _09571_/A sky130_fd_sc_hd__or2_1
XFILLER_70_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_196_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19863__RESET_B repeater267/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13107__A2 _18916_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16070__A _16637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12315__A0 _12313_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20017_ _20091_/CLK _20017_/D repeater235/X vssd1 vssd1 vccd1 vccd1 _20017_/Q sky130_fd_sc_hd__dfrtp_1
X_09828_ _19958_/Q vssd1 vssd1 vccd1 vccd1 _09866_/A sky130_fd_sc_hd__inv_2
XFILLER_171_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09759_ _09848_/B vssd1 vssd1 vccd1 vccd1 _09759_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__17105__S _17545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_199_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12770_ _12765_/Y _18834_/Q _19257_/Q _13557_/A _12769_/X vssd1 vssd1 vccd1 vccd1
+ _12783_/B sky130_fd_sc_hd__o221a_1
XPHY_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ _19512_/Q _11716_/X _16944_/X _11717_/X vssd1 vssd1 vccd1 vccd1 hold225/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_70_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16944__S _16946_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14440_ _18377_/Q _14436_/X _14437_/X _14439_/X vssd1 vssd1 vccd1 vccd1 _18377_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11652_ _18520_/Q _11652_/B vssd1 vssd1 vccd1 vccd1 _15271_/A sky130_fd_sc_hd__or2_1
XPHY_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10603_ _10553_/A _10600_/Y _10601_/X vssd1 vssd1 vccd1 vccd1 _10618_/A sky130_fd_sc_hd__o21ai_4
XPHY_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14371_ _18416_/Q _14367_/X _14356_/X _14369_/X vssd1 vssd1 vccd1 vccd1 _18416_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11583_ _11583_/A _11583_/B vssd1 vssd1 vccd1 vccd1 _11597_/A sky130_fd_sc_hd__or2_2
XFILLER_80_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16110_ _18085_/Q vssd1 vssd1 vccd1 vccd1 _16110_/Y sky130_fd_sc_hd__inv_2
X_13322_ _13322_/A _13322_/B _13483_/C vssd1 vssd1 vccd1 vccd1 _13463_/C sky130_fd_sc_hd__or3_1
XFILLER_196_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10534_ _18520_/Q vssd1 vssd1 vccd1 vccd1 _15289_/A sky130_fd_sc_hd__buf_1
X_17090_ _17486_/A0 _13105_/Y _17543_/S vssd1 vssd1 vccd1 vccd1 _17090_/X sky130_fd_sc_hd__mux2_1
XPHY_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16041_ _18108_/Q vssd1 vssd1 vccd1 vccd1 _16041_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19533__RESET_B repeater221/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10465_ _10471_/A vssd1 vssd1 vccd1 vccd1 _10472_/A sky130_fd_sc_hd__inv_2
X_13253_ _12313_/X _18871_/Q _13253_/S vssd1 vssd1 vccd1 vccd1 _18871_/D sky130_fd_sc_hd__mux2_1
XFILLER_129_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12204_ _19249_/Q _12198_/X _12092_/X _12199_/X vssd1 vssd1 vccd1 vccd1 _19249_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_123_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10396_ _10396_/A vssd1 vssd1 vccd1 vccd1 _10396_/Y sky130_fd_sc_hd__inv_2
X_13184_ _13184_/A vssd1 vssd1 vccd1 vccd1 _13184_/Y sky130_fd_sc_hd__inv_2
X_19800_ _19808_/CLK _19800_/D repeater222/X vssd1 vssd1 vccd1 vccd1 _19800_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_123_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12135_ _12171_/A vssd1 vssd1 vccd1 vccd1 _12172_/A sky130_fd_sc_hd__inv_2
X_17992_ _18169_/CLK _17992_/D vssd1 vssd1 vccd1 vccd1 _17992_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12306__B1 _12236_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19731_ _20055_/CLK _19731_/D repeater202/X vssd1 vssd1 vccd1 vccd1 _19731_/Q sky130_fd_sc_hd__dfrtp_1
X_16943_ _19487_/Q hold159/X _16946_/S vssd1 vssd1 vccd1 vccd1 _16943_/X sky130_fd_sc_hd__mux2_1
XFILLER_78_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12066_ _12066_/A _12187_/B vssd1 vssd1 vccd1 vccd1 _12121_/A sky130_fd_sc_hd__or2_4
XANTENNA__10740__B _13252_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11017_ _19654_/Q _19653_/Q _19655_/Q _11016_/X vssd1 vssd1 vccd1 vccd1 _11017_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__09722__B2 _19422_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19662_ _19846_/CLK _19662_/D repeater270/X vssd1 vssd1 vccd1 vccd1 _19662_/Q sky130_fd_sc_hd__dfrtp_1
X_16874_ _16873_/X _16630_/Y _17541_/S vssd1 vssd1 vccd1 vccd1 _16874_/X sky130_fd_sc_hd__mux2_1
XANTENNA__14059__B1 _14039_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15825_ _19685_/Q vssd1 vssd1 vccd1 vccd1 _15825_/Y sky130_fd_sc_hd__inv_2
X_18613_ _19041_/CLK _18613_/D repeater255/X vssd1 vssd1 vccd1 vccd1 _18613_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_237_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19593_ _19595_/CLK _19593_/D repeater282/X vssd1 vssd1 vccd1 vccd1 _19593_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_231_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17891__S1 _19632_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17015__S _17546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18544_ _18852_/CLK hold338/X repeater232/X vssd1 vssd1 vccd1 vccd1 _18545_/D sky130_fd_sc_hd__dfrtp_1
X_15756_ _18883_/Q _18881_/Q vssd1 vssd1 vccd1 vccd1 _15756_/X sky130_fd_sc_hd__or2_1
XFILLER_52_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_206_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12968_ _19191_/Q _12968_/B vssd1 vssd1 vccd1 vccd1 _12969_/D sky130_fd_sc_hd__or2_1
XFILLER_33_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14707_ _14707_/A vssd1 vssd1 vccd1 vccd1 _14707_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_205_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18475_ _19842_/CLK _18475_/D vssd1 vssd1 vccd1 vccd1 _18475_/Q sky130_fd_sc_hd__dfxtp_1
X_11919_ _19405_/Q _11914_/X _11918_/X _11915_/X vssd1 vssd1 vccd1 vccd1 _19405_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_206_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15687_ _15687_/A vssd1 vssd1 vccd1 vccd1 _15687_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16854__S _17522_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12899_ _12898_/Y _18950_/Q _19293_/Q _12893_/Y vssd1 vssd1 vccd1 vccd1 _12899_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_220_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17426_ _17425_/X _11366_/Y _17548_/S vssd1 vssd1 vccd1 vccd1 _17426_/X sky130_fd_sc_hd__mux2_1
X_14638_ _18260_/Q _14631_/A _09183_/X _14632_/A vssd1 vssd1 vccd1 vccd1 _18260_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_221_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17357_ _15963_/X _12790_/Y _17534_/S vssd1 vssd1 vccd1 vccd1 _17357_/X sky130_fd_sc_hd__mux2_1
X_14569_ hold321/X vssd1 vssd1 vccd1 vccd1 hold320/A sky130_fd_sc_hd__clkbuf_2
XFILLER_174_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16308_ _15219_/Y _15854_/A _16307_/Y _15976_/X vssd1 vssd1 vccd1 vccd1 _16308_/X
+ sky130_fd_sc_hd__o22a_1
X_17288_ _15963_/X _09518_/Y _17534_/S vssd1 vssd1 vccd1 vccd1 _17288_/X sky130_fd_sc_hd__mux2_1
X_19027_ _19437_/CLK _19027_/D repeater269/X vssd1 vssd1 vccd1 vccd1 _19027_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17685__S _17696_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15994__A _16637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16239_ _16634_/A vssd1 vssd1 vccd1 vccd1 _16555_/A sky130_fd_sc_hd__inv_2
XFILLER_115_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14298__B1 _13682_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08992_ _11935_/B vssd1 vssd1 vccd1 vccd1 _12130_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_141_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20108__RESET_B repeater217/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19929_ _19933_/CLK _19929_/D repeater235/X vssd1 vssd1 vccd1 vccd1 _19929_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_205_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10859__B1 _10448_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09613_ _20009_/Q _09612_/Y _09471_/B _09581_/X vssd1 vssd1 vccd1 vccd1 _20009_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_56_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_244_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17882__S1 _19632_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09544_ _20014_/Q _09541_/Y _09469_/A _19298_/Q _09543_/X vssd1 vssd1 vccd1 vccd1
+ _09545_/D sky130_fd_sc_hd__o221a_1
XFILLER_24_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14470__B1 _14417_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09475_ _09475_/A _09601_/A vssd1 vssd1 vccd1 vccd1 _09476_/B sky130_fd_sc_hd__or2_2
XPHY_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16764__S _17535_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18812__CLK _20115_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16514__A2 _15896_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19938__CLK _20013_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17595__S _17600_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10250_ _19516_/Q _19515_/Q _10250_/C vssd1 vssd1 vccd1 vccd1 _12130_/C sky130_fd_sc_hd__or3_4
XFILLER_105_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17475__A0 _17486_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11937__A _15772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15409__A _15413_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10181_ _10181_/A vssd1 vssd1 vccd1 vccd1 _15715_/B sky130_fd_sc_hd__inv_2
XFILLER_132_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10841__A _10841_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16939__S _16946_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13940_ _13911_/B _13817_/B _13938_/Y _13927_/X vssd1 vssd1 vccd1 vccd1 _18718_/D
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__09704__B2 _19429_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13871_ _19216_/Q vssd1 vssd1 vccd1 vccd1 _13871_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17873__S1 _19632_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_234_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15610_ _15610_/A _15610_/B vssd1 vssd1 vccd1 vccd1 _15610_/Y sky130_fd_sc_hd__nor2_1
X_12822_ _19243_/Q vssd1 vssd1 vccd1 vccd1 _12822_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16590_ _19042_/Q _16622_/B vssd1 vssd1 vccd1 vccd1 _16590_/Y sky130_fd_sc_hd__nand2_1
XFILLER_234_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14461__B1 _14405_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12487__B _12487_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15541_ _18579_/Q vssd1 vssd1 vccd1 vccd1 _15541_/Y sky130_fd_sc_hd__inv_2
X_12753_ _18809_/Q vssd1 vssd1 vccd1 vccd1 _13533_/A sky130_fd_sc_hd__inv_2
XPHY_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_199_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14983__A hold245/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11704_ _11704_/A vssd1 vssd1 vccd1 vccd1 _18622_/D sky130_fd_sc_hd__buf_1
X_18260_ _18260_/CLK _18260_/D vssd1 vssd1 vccd1 vccd1 _18260_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19785__RESET_B repeater203/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15472_ _15475_/B _15471_/Y _15459_/X vssd1 vssd1 vccd1 vccd1 _15472_/X sky130_fd_sc_hd__o21a_1
XFILLER_202_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12684_ _12698_/A vssd1 vssd1 vccd1 vccd1 _12684_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_42_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17211_ _17210_/X _11419_/Y _17548_/S vssd1 vssd1 vccd1 vccd1 _17211_/X sky130_fd_sc_hd__mux2_1
XPHY_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14423_ _14450_/A _14450_/B _15070_/C vssd1 vssd1 vccd1 vccd1 _14425_/A sky130_fd_sc_hd__or3_4
XPHY_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11635_ _11635_/A vssd1 vssd1 vccd1 vccd1 _11635_/Y sky130_fd_sc_hd__inv_2
X_18191_ _18198_/CLK _18191_/D vssd1 vssd1 vccd1 vccd1 _18191_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_118_HCLK_A clkbuf_opt_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17142_ _17141_/X _11348_/Y _17493_/S vssd1 vssd1 vccd1 vccd1 _17142_/X sky130_fd_sc_hd__mux2_1
X_14354_ _18425_/Q _14349_/X _14351_/X _14353_/X vssd1 vssd1 vccd1 vccd1 _18425_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11566_ _19024_/Q _11566_/B vssd1 vssd1 vccd1 vccd1 _11567_/A sky130_fd_sc_hd__or2_2
XFILLER_10_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13305_ _18860_/Q vssd1 vssd1 vccd1 vccd1 _13431_/C sky130_fd_sc_hd__inv_2
X_10517_ _10517_/A _11654_/B vssd1 vssd1 vccd1 vccd1 _10530_/C sky130_fd_sc_hd__or2_1
X_17073_ _16619_/Y _20111_/Q _17385_/S vssd1 vssd1 vccd1 vccd1 _17073_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14285_ _18458_/Q _14274_/A _13682_/X _14275_/A vssd1 vssd1 vccd1 vccd1 _18458_/D
+ sky130_fd_sc_hd__a22o_1
X_11497_ _11497_/A vssd1 vssd1 vccd1 vccd1 _11497_/Y sky130_fd_sc_hd__inv_2
XFILLER_170_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12527__B1 _12296_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16024_ _18228_/Q vssd1 vssd1 vccd1 vccd1 _16024_/Y sky130_fd_sc_hd__inv_2
X_13236_ _18882_/Q _13231_/X _18881_/Q _13230_/A vssd1 vssd1 vccd1 vccd1 _18882_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_40_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10448_ _10448_/A vssd1 vssd1 vccd1 vccd1 _10448_/X sky130_fd_sc_hd__buf_4
XFILLER_152_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13167_ _18916_/Q _13166_/Y _13162_/X _13167_/C1 vssd1 vssd1 vccd1 vccd1 _18916_/D
+ sky130_fd_sc_hd__o211a_1
X_10379_ _08921_/X _08964_/X _10321_/C _10321_/D vssd1 vssd1 vccd1 vccd1 _10379_/X
+ sky130_fd_sc_hd__o31a_1
X_12118_ _19303_/Q _12114_/X _11909_/X _12115_/X vssd1 vssd1 vccd1 vccd1 _19303_/D
+ sky130_fd_sc_hd__a22o_1
X_17975_ _20090_/CLK _17975_/D vssd1 vssd1 vccd1 vccd1 _17975_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13098_ _19172_/Q vssd1 vssd1 vccd1 vccd1 _16544_/A sky130_fd_sc_hd__inv_2
XFILLER_112_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16849__S _17490_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_0_0_HCLK clkbuf_3_1_0_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_1_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_242_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19714_ _19795_/CLK _19714_/D repeater218/X vssd1 vssd1 vccd1 vccd1 _19714_/Q sky130_fd_sc_hd__dfstp_1
X_16926_ _11708_/X _16926_/A1 _18624_/D vssd1 vssd1 vccd1 vccd1 _18623_/D sky130_fd_sc_hd__mux2_4
X_12049_ _19333_/Q _12043_/X _11922_/X _12044_/X vssd1 vssd1 vccd1 vccd1 _19333_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_65_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19645_ _19873_/CLK _19645_/D repeater262/X vssd1 vssd1 vccd1 vccd1 _19645_/Q sky130_fd_sc_hd__dfrtp_2
X_16857_ _15963_/X _09501_/Y _17534_/S vssd1 vssd1 vccd1 vccd1 _16857_/X sky130_fd_sc_hd__mux2_1
XANTENNA__17864__S1 _19634_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15808_ _18234_/Q vssd1 vssd1 vccd1 vccd1 _15808_/Y sky130_fd_sc_hd__inv_2
X_19576_ _19576_/CLK _19576_/D repeater268/X vssd1 vssd1 vccd1 vccd1 _19576_/Q sky130_fd_sc_hd__dfrtp_1
X_16788_ _16787_/X _15700_/Y _17474_/S vssd1 vssd1 vccd1 vccd1 _16788_/X sky130_fd_sc_hd__mux2_1
XFILLER_93_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15739_ _18667_/Q _18665_/Q _18666_/Q _15738_/X vssd1 vssd1 vccd1 vccd1 _18486_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_222_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18527_ _19825_/CLK _18527_/D repeater223/X vssd1 vssd1 vccd1 vccd1 _18527_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_34_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09260_ _12370_/A _12130_/B _12256_/C vssd1 vssd1 vccd1 vccd1 _15914_/A sky130_fd_sc_hd__or3_4
XFILLER_34_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18458_ _19842_/CLK _18458_/D vssd1 vssd1 vccd1 vccd1 _18458_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_221_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_3_5_0_HCLK_A clkbuf_3_5_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17409_ _17486_/A0 _09917_/Y _17543_/S vssd1 vssd1 vccd1 vccd1 _17409_/X sky130_fd_sc_hd__mux2_1
X_09191_ _20072_/Q _20071_/Q _20073_/Q _10133_/B _08983_/B vssd1 vssd1 vccd1 vccd1
+ _09192_/B sky130_fd_sc_hd__a41o_1
XFILLER_147_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18389_ _18441_/CLK _18389_/D vssd1 vssd1 vccd1 vccd1 _18389_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__19455__RESET_B repeater272/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_221_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12518__B1 hold270/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11757__A _11771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10661__A _10676_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11741__B2 _11738_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08975_ _20067_/Q vssd1 vssd1 vccd1 vccd1 _09205_/A sky130_fd_sc_hd__inv_2
XANTENNA__17209__A0 _15768_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17855__S1 _18759_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09527_ _09482_/A _19312_/Q _20010_/Q _09525_/Y _09526_/X vssd1 vssd1 vccd1 vccd1
+ _09528_/D sky130_fd_sc_hd__o221a_1
XFILLER_25_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09458_ _19379_/Q vssd1 vssd1 vccd1 vccd1 _09458_/Y sky130_fd_sc_hd__inv_2
XFILLER_169_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19196__RESET_B repeater188/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09389_ _19907_/Q vssd1 vssd1 vccd1 vccd1 _10101_/C sky130_fd_sc_hd__inv_1
X_11420_ _19127_/Q vssd1 vssd1 vccd1 vccd1 _11420_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19125__RESET_B hold370/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16499__A1 _16487_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11351_ _18961_/Q vssd1 vssd1 vccd1 vccd1 _11351_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17791__S0 _17923_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12509__B1 _12406_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10302_ _18598_/Q _15612_/A vssd1 vssd1 vccd1 vccd1 _15617_/A sky130_fd_sc_hd__or2_1
X_14070_ _19084_/Q _14025_/A _14069_/Y _18684_/Q vssd1 vssd1 vccd1 vccd1 _14070_/X
+ sky130_fd_sc_hd__o22a_1
X_11282_ _19003_/Q vssd1 vssd1 vccd1 vccd1 _11282_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13021_ _13021_/A _13021_/B _13021_/C vssd1 vssd1 vccd1 vccd1 _13024_/A sky130_fd_sc_hd__or3_4
X_10233_ _10230_/Y _19659_/Q _19832_/Q _10959_/A _10232_/X vssd1 vssd1 vccd1 vccd1
+ _10246_/B sky130_fd_sc_hd__o221a_1
XFILLER_140_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10164_ _19888_/Q _10155_/A _09108_/X _10156_/A vssd1 vssd1 vccd1 vccd1 _19888_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_79_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18760__RESET_B repeater196/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_239_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10095_ _19913_/Q _10094_/Y _10026_/A _10086_/B vssd1 vssd1 vccd1 vccd1 _19913_/D
+ sky130_fd_sc_hd__o211a_1
X_14972_ _18068_/Q _14965_/A _14814_/X _14966_/A vssd1 vssd1 vccd1 vccd1 _18068_/D
+ sky130_fd_sc_hd__a22o_1
X_17760_ _15195_/Y _13491_/Y _17762_/S vssd1 vssd1 vccd1 vccd1 _17760_/X sky130_fd_sc_hd__mux2_2
XFILLER_86_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13923_ _13914_/B _13827_/B _13921_/Y _13970_/C vssd1 vssd1 vccd1 vccd1 _18728_/D
+ sky130_fd_sc_hd__a211oi_2
X_16711_ _16798_/X _16493_/A _16803_/X _16512_/A vssd1 vssd1 vccd1 vccd1 _16711_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_19_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17691_ _15468_/X _19444_/Q _17696_/S vssd1 vssd1 vccd1 vccd1 _18561_/D sky130_fd_sc_hd__mux2_1
XANTENNA__17846__S1 _18759_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19430_ _19997_/CLK _19430_/D repeater185/X vssd1 vssd1 vccd1 vccd1 _19430_/Q sky130_fd_sc_hd__dfrtp_1
X_16642_ _16669_/A vssd1 vssd1 vccd1 vccd1 _16647_/B sky130_fd_sc_hd__buf_6
XFILLER_63_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13854_ _13851_/Y _18717_/Q _19206_/Q _13909_/C _13853_/X vssd1 vssd1 vccd1 vccd1
+ _13867_/A sky130_fd_sc_hd__o221a_1
XANTENNA__18858__CLK _18866_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14434__B1 _14405_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12805_ _19249_/Q vssd1 vssd1 vccd1 vccd1 _16646_/A sky130_fd_sc_hd__inv_2
XFILLER_34_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19361_ _19970_/CLK _19361_/D hold370/X vssd1 vssd1 vccd1 vccd1 _19361_/Q sky130_fd_sc_hd__dfrtp_1
X_16573_ _16683_/A vssd1 vssd1 vccd1 vccd1 _16573_/X sky130_fd_sc_hd__buf_2
X_13785_ _18727_/Q vssd1 vssd1 vccd1 vccd1 _13912_/C sky130_fd_sc_hd__inv_2
XFILLER_15_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10997_ _10993_/B _10978_/A _10996_/X _10989_/X _10996_/A vssd1 vssd1 vccd1 vccd1
+ _10998_/A sky130_fd_sc_hd__o32a_1
XFILLER_16_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18312_ _19847_/CLK _18312_/D vssd1 vssd1 vccd1 vccd1 _18312_/Q sky130_fd_sc_hd__dfxtp_1
X_15524_ _15537_/B vssd1 vssd1 vccd1 vccd1 _15530_/B sky130_fd_sc_hd__clkbuf_2
X_12736_ _19235_/Q vssd1 vssd1 vccd1 vccd1 _16469_/A sky130_fd_sc_hd__inv_2
XFILLER_16_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19292_ _19293_/CLK _19292_/D repeater187/X vssd1 vssd1 vccd1 vccd1 _19292_/Q sky130_fd_sc_hd__dfrtp_1
X_18243_ _19847_/CLK _18243_/D vssd1 vssd1 vccd1 vccd1 _18243_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15455_ _15479_/A _15455_/B vssd1 vssd1 vccd1 vccd1 _15455_/Y sky130_fd_sc_hd__nor2_1
XPHY_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12667_ _18989_/Q _12661_/X hold289/X _12664_/X vssd1 vssd1 vccd1 vccd1 _18989_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14406_ _18394_/Q _14395_/A _14405_/X _14396_/A vssd1 vssd1 vccd1 vccd1 _18394_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11618_ _11571_/A _11571_/B _11615_/Y _11645_/C vssd1 vssd1 vccd1 vccd1 _19558_/D
+ sky130_fd_sc_hd__a211oi_2
X_18174_ _18198_/CLK _18174_/D vssd1 vssd1 vccd1 vccd1 _18174_/Q sky130_fd_sc_hd__dfxtp_1
X_15386_ _15386_/A vssd1 vssd1 vccd1 vccd1 _15386_/Y sky130_fd_sc_hd__inv_2
XFILLER_156_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12598_ _12598_/A vssd1 vssd1 vccd1 vccd1 _12598_/X sky130_fd_sc_hd__clkbuf_2
XPHY_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17125_ _17473_/A0 _16526_/Y _17547_/S vssd1 vssd1 vccd1 vccd1 _17125_/X sky130_fd_sc_hd__mux2_1
XPHY_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08967__A2 _18778_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14337_ _14337_/A vssd1 vssd1 vccd1 vccd1 _14338_/A sky130_fd_sc_hd__inv_2
XFILLER_156_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11549_ _11549_/A vssd1 vssd1 vccd1 vccd1 _11639_/A sky130_fd_sc_hd__buf_1
XFILLER_171_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_183_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17782__S0 _17923_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17056_ _17055_/X _18911_/Q _17542_/S vssd1 vssd1 vccd1 vccd1 _17056_/X sky130_fd_sc_hd__mux2_1
XANTENNA__15162__B2 _15160_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14268_ _18952_/Q vssd1 vssd1 vccd1 vccd1 _14268_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_132_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18848__RESET_B repeater232/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17439__A0 _17473_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16007_ _18140_/Q vssd1 vssd1 vccd1 vccd1 _16007_/Y sky130_fd_sc_hd__inv_2
X_13219_ _18532_/Q _13219_/B vssd1 vssd1 vccd1 vccd1 _13220_/B sky130_fd_sc_hd__or2_1
X_14199_ _19119_/Q vssd1 vssd1 vccd1 vccd1 _14199_/Y sky130_fd_sc_hd__inv_2
XANTENNA__09392__A2 _09391_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09047__A hold318/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19633__CLK _19851_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16662__A1 _17014_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17958_ _20079_/CLK _17958_/D vssd1 vssd1 vccd1 vccd1 _17958_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16909_ _16908_/X _18909_/Q _17542_/S vssd1 vssd1 vccd1 vccd1 _16909_/X sky130_fd_sc_hd__mux2_1
XANTENNA__17837__S1 _18759_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17889_ _17885_/X _17886_/X _17887_/X _17888_/X _18760_/Q _18761_/Q vssd1 vssd1 vccd1
+ vccd1 _17889_/X sky130_fd_sc_hd__mux4_2
XFILLER_38_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19628_ _19630_/CLK _19628_/D repeater257/X vssd1 vssd1 vccd1 vccd1 _19628_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_226_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19636__RESET_B repeater258/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19559_ _19561_/CLK _19559_/D hold348/A vssd1 vssd1 vccd1 vccd1 _19559_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17203__S _17534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09312_ _18660_/Q _09305_/B _09311_/Y _18661_/Q _09305_/Y vssd1 vssd1 vccd1 vccd1
+ _18661_/D sky130_fd_sc_hd__a32o_1
XFILLER_15_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15512__A _15512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09243_ _10759_/B vssd1 vssd1 vccd1 vccd1 _10181_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__10656__A _19672_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09174_ _14705_/A vssd1 vssd1 vccd1 vccd1 _09174_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__13400__A1 _13399_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_101_HCLK_A clkbuf_4_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09080__A1 _20099_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_164_HCLK_A clkbuf_4_0_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17773__S0 _17923_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20123__RESET_B repeater196/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15153__B2 _15148_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18589__RESET_B repeater269/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11487__A _11487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18518__RESET_B repeater208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11714__A1 _12130_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11714__B2 _16950_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14113__C1 _14112_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16653__A1 _16964_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08958_ _19856_/Q vssd1 vssd1 vccd1 vccd1 _10322_/A sky130_fd_sc_hd__inv_2
XFILLER_243_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14664__B1 _14582_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17828__S1 _18750_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10920_ _19681_/Q vssd1 vssd1 vccd1 vccd1 _10920_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14416__B1 _14415_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10851_ _19711_/Q _10844_/A _10423_/X _10845_/A vssd1 vssd1 vccd1 vccd1 _19711_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17113__S _17318_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13570_ _18829_/Q _13569_/Y _13560_/X _13553_/B vssd1 vssd1 vccd1 vccd1 _18829_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_241_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10782_ _19888_/Q _10771_/A _19742_/Q _10774_/A vssd1 vssd1 vccd1 vccd1 _19742_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_201_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12521_ _19072_/Q _12519_/X _12353_/X _12520_/X vssd1 vssd1 vccd1 vccd1 _19072_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14038__A _19079_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15240_ _15304_/A vssd1 vssd1 vccd1 vccd1 _15259_/A sky130_fd_sc_hd__buf_1
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12452_ _19119_/Q _12450_/X _12389_/X _12451_/X vssd1 vssd1 vccd1 vccd1 _19119_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_184_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11403_ _19567_/Q vssd1 vssd1 vccd1 vccd1 _11580_/A sky130_fd_sc_hd__inv_2
X_15171_ _15171_/A vssd1 vssd1 vccd1 vccd1 _15172_/A sky130_fd_sc_hd__inv_2
XFILLER_126_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12383_ _19155_/Q _12374_/X _12382_/X _12378_/X vssd1 vssd1 vccd1 vccd1 _19155_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_153_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14122_ _14020_/A _14122_/A2 _14120_/Y _14118_/X vssd1 vssd1 vccd1 vccd1 _18690_/D
+ sky130_fd_sc_hd__a211oi_2
X_11334_ _18975_/Q vssd1 vssd1 vccd1 vccd1 _11334_/Y sky130_fd_sc_hd__inv_2
XFILLER_114_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_23_HCLK_A clkbuf_4_9_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_86_HCLK_A clkbuf_4_13_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14053_ _19063_/Q vssd1 vssd1 vccd1 vccd1 _14053_/Y sky130_fd_sc_hd__inv_2
X_18930_ _18947_/CLK _18930_/D repeater213/X vssd1 vssd1 vccd1 vccd1 _18930_/Q sky130_fd_sc_hd__dfrtp_1
X_11265_ _19582_/Q vssd1 vssd1 vccd1 vccd1 _11463_/A sky130_fd_sc_hd__inv_2
XFILLER_137_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13004_ _13004_/A _13004_/B vssd1 vssd1 vccd1 vccd1 _13014_/A sky130_fd_sc_hd__or2_1
X_10216_ _19826_/Q _10211_/X _10212_/Y _19653_/Q _10215_/X vssd1 vssd1 vccd1 vccd1
+ _10247_/B sky130_fd_sc_hd__o221a_1
X_18861_ _18866_/CLK _18861_/D repeater231/X vssd1 vssd1 vccd1 vccd1 _18861_/Q sky130_fd_sc_hd__dfrtp_1
X_11196_ _17718_/X _11191_/X _19613_/Q _11192_/X vssd1 vssd1 vccd1 vccd1 _19613_/D
+ sky130_fd_sc_hd__a22o_1
X_17812_ _18356_/Q _17996_/Q _18412_/Q _18396_/Q _17918_/S0 _18750_/Q vssd1 vssd1
+ vccd1 vccd1 _17812_/X sky130_fd_sc_hd__mux4_2
XFILLER_121_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10147_ hold321/X vssd1 vssd1 vccd1 vccd1 _10147_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_67_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18792_ _19647_/CLK _18792_/D repeater261/X vssd1 vssd1 vccd1 vccd1 _18792_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_153_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17743_ _15366_/X _19702_/Q _18508_/D vssd1 vssd1 vccd1 vccd1 _17743_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11844__B _16055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14955_ _18081_/Q _14952_/X _14921_/X _14954_/X vssd1 vssd1 vccd1 vccd1 _18081_/D
+ sky130_fd_sc_hd__a22o_1
X_10078_ _19919_/Q _10077_/Y _10026_/A _10036_/B vssd1 vssd1 vccd1 vccd1 _19919_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__17819__S1 _18752_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13906_ _13906_/A vssd1 vssd1 vccd1 vccd1 _13916_/A sky130_fd_sc_hd__inv_2
XFILLER_236_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14886_ _18121_/Q _14883_/X _14802_/X _14885_/X vssd1 vssd1 vccd1 vccd1 _18121_/D
+ sky130_fd_sc_hd__a22o_1
X_17674_ _15540_/X _19461_/Q _17683_/S vssd1 vssd1 vccd1 vccd1 _18578_/D sky130_fd_sc_hd__mux2_1
XFILLER_90_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19413_ _19905_/CLK _19413_/D repeater193/X vssd1 vssd1 vccd1 vccd1 _19413_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_223_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16625_ _17066_/X _16563_/X _17038_/X _16591_/X vssd1 vssd1 vccd1 vccd1 _16629_/A
+ sky130_fd_sc_hd__o22ai_4
X_13837_ _19213_/Q _13909_/B _19222_/Q _13831_/A vssd1 vssd1 vccd1 vccd1 _13837_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__15080__B1 _14780_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17023__S _17541_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16556_ _16556_/A vssd1 vssd1 vccd1 vccd1 _16556_/X sky130_fd_sc_hd__clkbuf_2
X_19344_ _19952_/CLK _19344_/D repeater244/X vssd1 vssd1 vccd1 vccd1 _19344_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13768_ _18743_/Q _18744_/Q _13772_/S vssd1 vssd1 vccd1 vccd1 _18744_/D sky130_fd_sc_hd__mux2_1
XANTENNA__20013__CLK _20013_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15507_ _15511_/B _15506_/X _15483_/X vssd1 vssd1 vccd1 vccd1 _15507_/X sky130_fd_sc_hd__o21a_1
X_12719_ _18956_/Q vssd1 vssd1 vccd1 vccd1 _14810_/A sky130_fd_sc_hd__clkbuf_2
X_16487_ _17230_/X _16505_/A _17308_/X _16506_/A vssd1 vssd1 vccd1 vccd1 _16487_/X
+ sky130_fd_sc_hd__o22a_2
X_19275_ _19282_/CLK _19275_/D repeater216/X vssd1 vssd1 vccd1 vccd1 _19275_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__16862__S _17547_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13699_ _17760_/X _13523_/Y _13698_/X vssd1 vssd1 vccd1 vccd1 _18764_/D sky130_fd_sc_hd__a21oi_1
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15438_ _18633_/Q _17570_/X _15436_/A _15437_/X vssd1 vssd1 vccd1 vccd1 _15438_/X
+ sky130_fd_sc_hd__a22o_1
X_18226_ _18412_/CLK _18226_/D vssd1 vssd1 vccd1 vccd1 _18226_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_248_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09062__A1 _20105_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15369_ _19785_/Q _10645_/B _10646_/B vssd1 vssd1 vccd1 vccd1 _15369_/X sky130_fd_sc_hd__a21bo_1
XFILLER_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18157_ _18460_/CLK _18157_/D vssd1 vssd1 vccd1 vccd1 _18157_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12691__A _12698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17108_ _17107_/X _18818_/Q _17536_/S vssd1 vssd1 vccd1 vccd1 _17108_/X sky130_fd_sc_hd__mux2_2
Xhold304 HWDATA[26] vssd1 vssd1 vccd1 vccd1 input56/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold315 input51/X vssd1 vssd1 vccd1 vccd1 hold315/X sky130_fd_sc_hd__dlygate4sd3_1
X_18088_ _18137_/CLK _18088_/D vssd1 vssd1 vccd1 vccd1 _18088_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold326 input64/X vssd1 vssd1 vccd1 vccd1 hold326/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__18682__RESET_B repeater252/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold337 HWDATA[1] vssd1 vssd1 vccd1 vccd1 input49/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold348 hold348/A vssd1 vssd1 vccd1 vccd1 hold348/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17693__S _17696_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17039_ _15768_/Y _11217_/Y _17546_/S vssd1 vssd1 vccd1 vccd1 _17039_/X sky130_fd_sc_hd__mux2_1
X_09930_ _19343_/Q vssd1 vssd1 vccd1 vccd1 _09930_/Y sky130_fd_sc_hd__inv_2
XFILLER_172_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold359 hold359/A vssd1 vssd1 vccd1 vccd1 hold359/X sky130_fd_sc_hd__dlygate4sd3_1
X_20050_ _20050_/CLK _20050_/D repeater206/X vssd1 vssd1 vccd1 vccd1 _20050_/Q sky130_fd_sc_hd__dfrtp_1
X_09861_ _09861_/A _09861_/B vssd1 vssd1 vccd1 vccd1 _09978_/A sky130_fd_sc_hd__or2_1
XFILLER_86_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09792_ _09792_/A _09792_/B vssd1 vssd1 vccd1 vccd1 _09797_/A sky130_fd_sc_hd__or2_1
XFILLER_39_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13525__A1_N _18761_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09505__A _19323_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater154 _17413_/S vssd1 vssd1 vccd1 vccd1 _17529_/S sky130_fd_sc_hd__buf_8
XFILLER_38_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater165 _17543_/S vssd1 vssd1 vccd1 vccd1 _17546_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_227_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrepeater176 _17524_/S vssd1 vssd1 vccd1 vccd1 _17513_/S sky130_fd_sc_hd__buf_8
XPHY_4308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater187 repeater188/X vssd1 vssd1 vccd1 vccd1 repeater187/X sky130_fd_sc_hd__buf_4
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrepeater198 repeater199/X vssd1 vssd1 vccd1 vccd1 repeater198/X sky130_fd_sc_hd__clkbuf_8
XPHY_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19470__RESET_B repeater274/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11880__B1 _09021_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_94_HCLK clkbuf_4_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19956_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_42_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16772__S _17534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09226_ _18645_/Q vssd1 vssd1 vccd1 vccd1 _09226_/X sky130_fd_sc_hd__buf_1
XFILLER_166_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16571__B1 _17566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09157_ _09154_/A _09156_/A _15321_/A _15322_/B vssd1 vssd1 vccd1 vccd1 _09157_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_108_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09088_ _20097_/Q _09084_/X _09086_/X _09087_/X vssd1 vssd1 vccd1 vccd1 _20097_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16323__B1 _17373_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_0_HCLK clkbuf_4_0_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _18142_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__12106__A _12121_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11699__B1 _10868_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11050_ _19644_/Q vssd1 vssd1 vccd1 vccd1 _14335_/A sky130_fd_sc_hd__buf_1
XFILLER_77_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10001_ _10001_/A vssd1 vssd1 vccd1 vccd1 _10001_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16626__A1 _17068_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15417__A _15419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17108__S _17536_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_237_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_4_8_0_HCLK_A clkbuf_4_9_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19558__RESET_B hold348/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16947__S _16950_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14740_ _18204_/Q _14733_/A _14727_/X _14734_/A vssd1 vssd1 vccd1 vccd1 _18204_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_218_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11952_ _19390_/Q _11948_/X hold305/X _11949_/X vssd1 vssd1 vccd1 vccd1 _19390_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_17_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10903_ _19685_/Q _10894_/A _10870_/X _10895_/A vssd1 vssd1 vccd1 vccd1 _19685_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_17_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14671_ _14671_/A vssd1 vssd1 vccd1 vccd1 _14671_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_72_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11883_ _19428_/Q _11875_/X _09027_/X _11878_/X vssd1 vssd1 vccd1 vccd1 _19428_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_45_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_233_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16410_ _18345_/Q vssd1 vssd1 vccd1 vccd1 _16410_/Y sky130_fd_sc_hd__inv_2
X_13622_ _18802_/Q _13499_/X _18802_/Q _13620_/A vssd1 vssd1 vccd1 vccd1 _13622_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_10834_ _19719_/Q vssd1 vssd1 vccd1 vccd1 _10834_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19140__RESET_B hold348/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17390_ _17389_/X _19197_/Q _17545_/S vssd1 vssd1 vccd1 vccd1 _17390_/X sky130_fd_sc_hd__mux2_1
X_16341_ _18408_/Q vssd1 vssd1 vccd1 vccd1 _16341_/Y sky130_fd_sc_hd__inv_2
XFILLER_198_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13553_ _13553_/A _13553_/B vssd1 vssd1 vccd1 vccd1 _13566_/A sky130_fd_sc_hd__or2_1
X_10765_ _18643_/Q _10765_/B vssd1 vssd1 vccd1 vccd1 _10766_/B sky130_fd_sc_hd__nand2_1
XFILLER_185_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12504_ _19083_/Q _12498_/X _12398_/X _12499_/X vssd1 vssd1 vccd1 vccd1 _19083_/D
+ sky130_fd_sc_hd__a22o_1
X_19060_ _19630_/CLK _19060_/D repeater257/X vssd1 vssd1 vccd1 vccd1 _19060_/Q sky130_fd_sc_hd__dfrtp_1
X_16272_ _18247_/Q _16433_/B vssd1 vssd1 vccd1 vccd1 _16272_/X sky130_fd_sc_hd__or2_1
X_13484_ _13322_/B _13486_/A _13322_/A vssd1 vssd1 vccd1 vccd1 _13485_/B sky130_fd_sc_hd__o21a_1
XFILLER_9_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10696_ _10448_/A _17749_/X _17749_/S _10694_/Y _19779_/Q vssd1 vssd1 vccd1 vccd1
+ _19779_/D sky130_fd_sc_hd__a32o_1
XFILLER_12_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18011_ _18959_/CLK _18011_/D vssd1 vssd1 vccd1 vccd1 _18011_/Q sky130_fd_sc_hd__dfxtp_1
X_15223_ _15223_/A vssd1 vssd1 vccd1 vccd1 _15223_/Y sky130_fd_sc_hd__inv_2
XFILLER_185_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12435_ _19126_/Q _12400_/A _12241_/X _12402_/A vssd1 vssd1 vccd1 vccd1 _19126_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_166_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15154_ _17955_/Q _15147_/A _14711_/A _15148_/A vssd1 vssd1 vccd1 vccd1 _17955_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_5_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11839__B _15776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12366_ _19161_/Q _12361_/X _12234_/X _12362_/X vssd1 vssd1 vccd1 vccd1 _19161_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_154_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14105_ _18699_/Q _14104_/Y _14096_/X _14030_/B vssd1 vssd1 vccd1 vccd1 _18699_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_141_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11317_ _18973_/Q vssd1 vssd1 vccd1 vccd1 _11317_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15085_ _15085_/A vssd1 vssd1 vccd1 vccd1 _15085_/X sky130_fd_sc_hd__clkbuf_2
X_19962_ _19964_/CLK _19962_/D hold371/X vssd1 vssd1 vccd1 vccd1 _19962_/Q sky130_fd_sc_hd__dfrtp_2
X_12297_ _19200_/Q _12290_/X _12296_/X _12291_/X vssd1 vssd1 vccd1 vccd1 _19200_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12016__A _12016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14036_ _19069_/Q _14011_/A _19078_/Q _14019_/A vssd1 vssd1 vccd1 vccd1 _14036_/X
+ sky130_fd_sc_hd__a22o_1
X_18913_ _19222_/CLK _18913_/D repeater188/X vssd1 vssd1 vccd1 vccd1 _18913_/Q sky130_fd_sc_hd__dfrtp_1
X_11248_ _11248_/A _11248_/B _11248_/C _11248_/D vssd1 vssd1 vccd1 vccd1 _11248_/X
+ sky130_fd_sc_hd__and4_1
X_19893_ _20055_/CLK _19893_/D repeater205/X vssd1 vssd1 vccd1 vccd1 _19893_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12351__A1 _19170_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17018__S _17318_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18844_ _18866_/CLK _18844_/D repeater232/X vssd1 vssd1 vccd1 vccd1 _18844_/Q sky130_fd_sc_hd__dfrtp_1
X_11179_ _17705_/X _11176_/X _19626_/Q _11178_/X vssd1 vssd1 vccd1 vccd1 _19626_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_68_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19981__RESET_B repeater192/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18775_ _19855_/CLK _18775_/D repeater265/X vssd1 vssd1 vccd1 vccd1 _18775_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__19299__RESET_B repeater241/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_227_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15987_ _15985_/Y _15831_/A _15986_/Y _15842_/X vssd1 vssd1 vccd1 vccd1 _15987_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__16857__S _17534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17726_ _19674_/Q _19687_/Q _18510_/Q vssd1 vssd1 vccd1 vccd1 _17726_/X sky130_fd_sc_hd__mux2_1
XFILLER_35_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14938_ _15109_/A _15145_/B _14951_/C vssd1 vssd1 vccd1 vccd1 _14940_/A sky130_fd_sc_hd__or3_4
XFILLER_235_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17657_ _15607_/X _19032_/Q _17664_/S vssd1 vssd1 vccd1 vccd1 _18595_/D sky130_fd_sc_hd__mux2_1
XANTENNA__15053__B1 _15000_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14869_ _18130_/Q _14859_/A _14868_/X _14860_/A vssd1 vssd1 vccd1 vccd1 _18130_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_35_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16608_ _19458_/Q vssd1 vssd1 vccd1 vccd1 _16608_/Y sky130_fd_sc_hd__inv_2
X_17588_ _15361_/X _19715_/Q _17600_/S vssd1 vssd1 vccd1 vccd1 _17588_/X sky130_fd_sc_hd__mux2_1
XFILLER_195_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19327_ _19905_/CLK _19327_/D repeater191/X vssd1 vssd1 vccd1 vccd1 _19327_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__11614__B1 _11617_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17688__S _17696_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16539_ _17178_/X _16684_/A _17166_/X _16493_/X vssd1 vssd1 vccd1 vccd1 _16539_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_188_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19258_ _19324_/CLK _19258_/D repeater237/X vssd1 vssd1 vccd1 vccd1 _19258_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18863__RESET_B repeater231/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09011_ _19503_/Q _11832_/B _11832_/C vssd1 vssd1 vccd1 vccd1 _11996_/A sky130_fd_sc_hd__or3_4
XFILLER_136_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18209_ _19630_/CLK _18209_/D vssd1 vssd1 vccd1 vccd1 _18209_/Q sky130_fd_sc_hd__dfxtp_1
X_19189_ _19293_/CLK _19189_/D repeater186/X vssd1 vssd1 vccd1 vccd1 _19189_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_163_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold134 HADDR[18] vssd1 vssd1 vccd1 vccd1 input10/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold145 input7/X vssd1 vssd1 vccd1 vccd1 hold145/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 input6/X vssd1 vssd1 vccd1 vccd1 hold156/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold167 hold167/A vssd1 vssd1 vccd1 vccd1 hold167/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_160_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20102_ _20107_/CLK _20102_/D repeater234/X vssd1 vssd1 vccd1 vccd1 _20102_/Q sky130_fd_sc_hd__dfrtp_1
Xhold178 HADDR[9] vssd1 vssd1 vccd1 vccd1 input32/A sky130_fd_sc_hd__dlygate4sd3_1
X_09913_ _19348_/Q vssd1 vssd1 vccd1 vccd1 _16588_/A sky130_fd_sc_hd__inv_2
Xhold189 hold356/X vssd1 vssd1 vccd1 vccd1 hold355/A sky130_fd_sc_hd__dlygate4sd3_1
X_20033_ _20035_/CLK _20033_/D repeater240/X vssd1 vssd1 vccd1 vccd1 _20033_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__11765__A _11772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09844_ _19942_/Q vssd1 vssd1 vccd1 vccd1 _09851_/A sky130_fd_sc_hd__inv_2
XFILLER_219_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17900__S0 _17913_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19651__RESET_B repeater261/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09775_ _09775_/A vssd1 vssd1 vccd1 vccd1 _09775_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16767__S _17385_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_227_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09510__A2 _19323_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_214_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12596__A _14273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_215_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15044__B1 _15006_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17598__S _17600_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10550_ _10582_/A _19811_/Q _19812_/Q vssd1 vssd1 vccd1 vccd1 _10551_/A sky130_fd_sc_hd__or3b_2
XFILLER_183_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09209_ _18644_/Q _18645_/Q _18646_/Q _18647_/Q vssd1 vssd1 vccd1 vccd1 _09238_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_167_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10481_ _18546_/Q vssd1 vssd1 vccd1 vccd1 _15389_/A sky130_fd_sc_hd__clkbuf_2
X_12220_ _12229_/A vssd1 vssd1 vccd1 vccd1 _12220_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_204_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12151_ _12151_/A vssd1 vssd1 vccd1 vccd1 _12151_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_136_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11102_ _19634_/Q _11101_/X _19634_/Q _11101_/X vssd1 vssd1 vccd1 vccd1 _11103_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_118_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12082_ _12094_/A vssd1 vssd1 vccd1 vccd1 _12082_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_101_HCLK clkbuf_4_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _18908_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_111_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11033_ _19652_/Q _11032_/X _19652_/Q _11032_/X vssd1 vssd1 vccd1 vccd1 _19652_/D
+ sky130_fd_sc_hd__o2bb2a_1
X_15910_ _15999_/A vssd1 vssd1 vccd1 vccd1 _16505_/A sky130_fd_sc_hd__clkbuf_2
X_16890_ _16889_/X _14060_/Y _17544_/S vssd1 vssd1 vccd1 vccd1 _16890_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16075__A2 _16002_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15841_ _19673_/Q vssd1 vssd1 vccd1 vccd1 _15841_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14086__B2 _18681_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16480__C1 _16479_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12097__B1 _12095_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18560_ _19992_/CLK _18560_/D repeater193/X vssd1 vssd1 vccd1 vccd1 _18560_/Q sky130_fd_sc_hd__dfrtp_1
X_12984_ _18940_/Q _12983_/Y _12980_/A _12883_/B vssd1 vssd1 vccd1 vccd1 _18940_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_45_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15772_ _15772_/A vssd1 vssd1 vccd1 vccd1 _16723_/B sky130_fd_sc_hd__inv_2
XFILLER_94_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17511_ _17510_/X _15880_/Y _17539_/S vssd1 vssd1 vccd1 vccd1 _17511_/X sky130_fd_sc_hd__mux2_2
XFILLER_245_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11935_ _12130_/A _11935_/B _12370_/C vssd1 vssd1 vccd1 vccd1 _15897_/A sky130_fd_sc_hd__or3_4
X_14723_ _14791_/A vssd1 vssd1 vccd1 vccd1 _14723_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_output113_A _15780_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18491_ _19720_/CLK _18491_/D repeater201/X vssd1 vssd1 vccd1 vccd1 _18491_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_33_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14654_ _14680_/A _15839_/A vssd1 vssd1 vccd1 vccd1 _16115_/A sky130_fd_sc_hd__or2_2
X_17442_ _17441_/X _15452_/Y _17518_/S vssd1 vssd1 vccd1 vccd1 _17442_/X sky130_fd_sc_hd__mux2_1
XFILLER_233_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11866_ _11848_/Y _11856_/Y _11862_/Y _19435_/Q _11865_/X vssd1 vssd1 vccd1 vccd1
+ _19435_/D sky130_fd_sc_hd__a32o_1
XFILLER_220_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13605_ _18809_/Q _13604_/Y _13591_/X _13534_/B vssd1 vssd1 vccd1 vccd1 _18809_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_3971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10817_ _17621_/X _10809_/A _19726_/Q _10810_/A vssd1 vssd1 vccd1 vccd1 _19726_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_32_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14585_ _18290_/Q _14573_/A hold320/X _14574_/A vssd1 vssd1 vccd1 vccd1 _18290_/D
+ sky130_fd_sc_hd__a22o_1
X_17373_ _17372_/X _17859_/X _17568_/S vssd1 vssd1 vccd1 vccd1 _17373_/X sky130_fd_sc_hd__mux2_2
XPHY_3993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11797_ _19463_/Q _11793_/X hold305/X _11794_/X vssd1 vssd1 vccd1 vccd1 _19463_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_220_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17301__S _17386_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19112_ _19115_/CLK _19112_/D hold353/X vssd1 vssd1 vccd1 vccd1 _19112_/Q sky130_fd_sc_hd__dfrtp_2
X_13536_ _13536_/A _13536_/B vssd1 vssd1 vccd1 vccd1 _13537_/C sky130_fd_sc_hd__or2_2
XANTENNA__15610__A _15610_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16324_ _17362_/X _15997_/X _17365_/X _15998_/X _16323_/X vssd1 vssd1 vccd1 vccd1
+ _16324_/X sky130_fd_sc_hd__o221a_2
XFILLER_201_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10748_ _19759_/Q _10741_/X _10421_/X _10743_/X vssd1 vssd1 vccd1 vccd1 _19759_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_185_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16255_ _18119_/Q vssd1 vssd1 vccd1 vccd1 _16255_/Y sky130_fd_sc_hd__inv_2
X_19043_ _19597_/CLK _19043_/D repeater255/X vssd1 vssd1 vccd1 vccd1 _19043_/Q sky130_fd_sc_hd__dfrtp_1
X_13467_ _13467_/A _13476_/A vssd1 vssd1 vccd1 vccd1 _13468_/B sky130_fd_sc_hd__or2_1
X_10679_ _17740_/X _10676_/X _19785_/Q _10677_/X vssd1 vssd1 vccd1 vccd1 _19785_/D
+ sky130_fd_sc_hd__a22o_1
X_15206_ _18513_/Q vssd1 vssd1 vccd1 vccd1 _15206_/Y sky130_fd_sc_hd__inv_2
X_12418_ _19139_/Q _12412_/X hold256/X _12414_/X vssd1 vssd1 vccd1 vccd1 _19139_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12021__B1 _09049_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16186_ _18078_/Q vssd1 vssd1 vccd1 vccd1 _16186_/Y sky130_fd_sc_hd__inv_2
X_13398_ _20092_/Q vssd1 vssd1 vccd1 vccd1 _13398_/Y sky130_fd_sc_hd__inv_4
XFILLER_142_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15137_ _17968_/Q _15134_/X hold247/X _15136_/X vssd1 vssd1 vccd1 vccd1 _17968_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_245_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12349_ _19171_/Q _12341_/X hold256/X _12342_/X vssd1 vssd1 vccd1 vccd1 _19171_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_126_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15068_ _18011_/Q _15060_/A _14816_/A _15061_/A vssd1 vssd1 vccd1 vccd1 _18011_/D
+ sky130_fd_sc_hd__a22o_1
X_19945_ _19976_/CLK _19945_/D repeater244/X vssd1 vssd1 vccd1 vccd1 _19945_/Q sky130_fd_sc_hd__dfrtp_1
X_14019_ _14019_/A _14123_/A vssd1 vssd1 vccd1 vccd1 _14020_/B sky130_fd_sc_hd__or2_2
XFILLER_96_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19876_ _19900_/CLK _19876_/D repeater197/X vssd1 vssd1 vccd1 vccd1 _19876_/Q sky130_fd_sc_hd__dfstp_4
XFILLER_229_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18827_ _18827_/CLK _18827_/D repeater217/X vssd1 vssd1 vccd1 vccd1 _18827_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_67_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09560_ _19325_/Q vssd1 vssd1 vccd1 vccd1 _09560_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18758_ _20123_/CLK _18758_/D repeater195/X vssd1 vssd1 vccd1 vccd1 _18758_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_243_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17709_ _15431_/X _19768_/Q _18546_/D vssd1 vssd1 vccd1 vccd1 _17709_/X sky130_fd_sc_hd__mux2_1
X_09491_ _09491_/A _09574_/A vssd1 vssd1 vccd1 vccd1 _09492_/B sky130_fd_sc_hd__or2_1
X_18689_ _18701_/CLK _18689_/D hold359/X vssd1 vssd1 vccd1 vccd1 _18689_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__15026__B1 _14992_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17211__S _17548_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12012__B1 _09033_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_124_HCLK clkbuf_4_4_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19566_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_219_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20016_ _20091_/CLK _20016_/D repeater236/X vssd1 vssd1 vccd1 vccd1 _20016_/Q sky130_fd_sc_hd__dfrtp_1
X_09827_ _19959_/Q vssd1 vssd1 vccd1 vccd1 _09867_/A sky130_fd_sc_hd__inv_2
XFILLER_104_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12079__B1 _12078_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09758_ _19999_/Q _19998_/Q _09758_/C vssd1 vssd1 vccd1 vccd1 _09758_/X sky130_fd_sc_hd__and3_1
XANTENNA__11826__B1 _10863_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09689_ _09689_/A _09689_/B _09689_/C _09689_/D vssd1 vssd1 vccd1 vccd1 _09728_/A
+ sky130_fd_sc_hd__and4_1
XPHY_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15017__B1 _15002_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ _19513_/Q _11716_/X _16945_/X _11717_/X vssd1 vssd1 vccd1 vccd1 hold224/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_64_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11651_ _11651_/A _11651_/B vssd1 vssd1 vccd1 vccd1 _11656_/A sky130_fd_sc_hd__or2_1
XPHY_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18714__RESET_B repeater252/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10602_ _18508_/Q _10909_/A _10616_/C _10583_/A _10601_/X vssd1 vssd1 vccd1 vccd1
+ _19813_/D sky130_fd_sc_hd__a32o_1
XANTENNA__17121__S _17546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14370_ _18417_/Q _14367_/X _14351_/X _14369_/X vssd1 vssd1 vccd1 vccd1 _18417_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11582_ _11582_/A _11600_/A vssd1 vssd1 vccd1 vccd1 _11583_/B sky130_fd_sc_hd__or2_1
XPHY_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13321_ _18838_/Q vssd1 vssd1 vccd1 vccd1 _13483_/C sky130_fd_sc_hd__clkinvlp_4
XFILLER_80_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10533_ _15389_/A _11672_/C vssd1 vssd1 vccd1 vccd1 _10537_/B sky130_fd_sc_hd__nand2_1
XPHY_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16960__S _17534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16040_ _18100_/Q vssd1 vssd1 vccd1 vccd1 _16040_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13252_ _14245_/A _15821_/B _14245_/C _13252_/D vssd1 vssd1 vccd1 vccd1 _13253_/S
+ sky130_fd_sc_hd__or4_4
XANTENNA_input74_A RsRx_S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10464_ _18549_/Q _18548_/Q vssd1 vssd1 vccd1 vccd1 _10471_/A sky130_fd_sc_hd__or2_2
XFILLER_170_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12203_ _19250_/Q _12198_/X _12090_/X _12199_/X vssd1 vssd1 vccd1 vccd1 _19250_/D
+ sky130_fd_sc_hd__a22o_1
X_13183_ _13079_/A _13183_/A2 _13179_/Y _13182_/X vssd1 vssd1 vccd1 vccd1 _18907_/D
+ sky130_fd_sc_hd__a211oi_2
X_10395_ _10404_/A _14476_/A vssd1 vssd1 vccd1 vccd1 _10396_/A sky130_fd_sc_hd__or2_1
XANTENNA__19397__CLK _20091_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08979__A _17605_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12134_ _12150_/A vssd1 vssd1 vccd1 vccd1 _12134_/X sky130_fd_sc_hd__clkbuf_2
X_17991_ _18169_/CLK _17991_/D vssd1 vssd1 vccd1 vccd1 _17991_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19730_ _20055_/CLK _19730_/D repeater202/X vssd1 vssd1 vccd1 vccd1 _19730_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_111_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16942_ _19486_/Q hold145/X _16946_/S vssd1 vssd1 vccd1 vccd1 _16942_/X sky130_fd_sc_hd__mux2_1
X_12065_ _11991_/X _19326_/Q _12065_/S vssd1 vssd1 vccd1 vccd1 _19326_/D sky130_fd_sc_hd__mux2_1
XANTENNA__17245__A1 _18821_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11016_ _10224_/X _10211_/X _10956_/C vssd1 vssd1 vccd1 vccd1 _11016_/X sky130_fd_sc_hd__o21a_1
X_19661_ _19846_/CLK _19661_/D repeater270/X vssd1 vssd1 vccd1 vccd1 _19661_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_93_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16873_ _17486_/A0 _13148_/Y _17543_/S vssd1 vssd1 vccd1 vccd1 _16873_/X sky130_fd_sc_hd__mux2_1
X_18612_ _19041_/CLK _18612_/D repeater266/X vssd1 vssd1 vccd1 vccd1 _18612_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_64_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15824_ _16303_/A vssd1 vssd1 vccd1 vccd1 _15864_/B sky130_fd_sc_hd__clkbuf_4
X_19592_ _19595_/CLK _19592_/D hold346/A vssd1 vssd1 vccd1 vccd1 _19592_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_161_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18543_ _18886_/CLK _18543_/D repeater221/X vssd1 vssd1 vccd1 vccd1 _18543_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__11817__B1 _09075_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15755_ _18526_/D _15755_/B vssd1 vssd1 vccd1 vccd1 _18547_/D sky130_fd_sc_hd__nor2_1
X_12967_ _12967_/A _12967_/B _12967_/C _12966_/X vssd1 vssd1 vccd1 vccd1 _12967_/X
+ sky130_fd_sc_hd__or4b_4
X_11918_ _12232_/A vssd1 vssd1 vccd1 vccd1 _11918_/X sky130_fd_sc_hd__buf_2
X_14706_ _18223_/Q _14698_/X _14705_/X _14701_/X vssd1 vssd1 vccd1 vccd1 _18223_/D
+ sky130_fd_sc_hd__a22o_1
X_18474_ _19842_/CLK _18474_/D vssd1 vssd1 vccd1 vccd1 _18474_/Q sky130_fd_sc_hd__dfxtp_1
X_15686_ _18614_/Q _15686_/B vssd1 vssd1 vccd1 vccd1 _15687_/A sky130_fd_sc_hd__or2_1
XFILLER_61_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12898_ _19293_/Q vssd1 vssd1 vccd1 vccd1 _12898_/Y sky130_fd_sc_hd__inv_2
XPHY_4480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17425_ _17424_/X _11337_/Y _17459_/S vssd1 vssd1 vccd1 vccd1 _17425_/X sky130_fd_sc_hd__mux2_1
XFILLER_220_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11849_ _19434_/Q vssd1 vssd1 vccd1 vccd1 _11851_/A sky130_fd_sc_hd__inv_2
X_14637_ _18261_/Q _14630_/X _09180_/X _14632_/X vssd1 vssd1 vccd1 vccd1 _18261_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_221_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12242__B1 _12241_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17356_ _17355_/X _09470_/A _17530_/S vssd1 vssd1 vccd1 vccd1 _17356_/X sky130_fd_sc_hd__mux2_1
XFILLER_147_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14568_ _18299_/Q _14559_/A _14567_/X _14560_/A vssd1 vssd1 vccd1 vccd1 _18299_/D
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_147_HCLK clkbuf_4_1_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19855_/CLK sky130_fd_sc_hd__clkbuf_16
X_16307_ _19678_/Q vssd1 vssd1 vccd1 vccd1 _16307_/Y sky130_fd_sc_hd__inv_2
XFILLER_159_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13519_ _18765_/Q vssd1 vssd1 vccd1 vccd1 _14642_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__16870__S _17534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17287_ _17286_/X _13883_/Y _17545_/S vssd1 vssd1 vccd1 vccd1 _17287_/X sky130_fd_sc_hd__mux2_1
X_14499_ _18340_/Q _14492_/A _12729_/X _14493_/A vssd1 vssd1 vccd1 vccd1 _18340_/D
+ sky130_fd_sc_hd__a22o_1
X_19026_ _19157_/CLK _19026_/D repeater266/X vssd1 vssd1 vccd1 vccd1 _19026_/Q sky130_fd_sc_hd__dfrtp_4
X_16238_ _16238_/A vssd1 vssd1 vccd1 vccd1 _16638_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_133_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16169_ _11023_/Y _18227_/Q _16168_/X vssd1 vssd1 vccd1 vccd1 _16169_/Y sky130_fd_sc_hd__o21ai_1
X_08991_ _19517_/Q vssd1 vssd1 vccd1 vccd1 _11935_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_69_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19928_ _19933_/CLK _19928_/D repeater230/X vssd1 vssd1 vccd1 vccd1 _19928_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_102_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19859_ _19859_/CLK _19859_/D repeater262/X vssd1 vssd1 vccd1 vccd1 _19859_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_244_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09612_ _09612_/A vssd1 vssd1 vccd1 vccd1 _09612_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17206__S _17543_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16995__A0 _16994_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09543_ _20026_/Q _16647_/A _09486_/A _19316_/Q vssd1 vssd1 vccd1 vccd1 _09543_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_37_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09474_ _09474_/A _09474_/B _09605_/A vssd1 vssd1 vccd1 vccd1 _09601_/A sky130_fd_sc_hd__or3_1
XFILLER_169_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12481__B1 _12302_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_240_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18144__CLK _18169_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_200_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12233__B1 _12232_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16780__S _17413_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18294__CLK _19847_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10180_ _19878_/Q _10174_/X _09108_/X _10175_/X vssd1 vssd1 vccd1 vccd1 _19878_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_59_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12114__A _12121_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09704__A2 _19405_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_28_HCLK clkbuf_4_9_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20057_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_120_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17116__S _17513_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13870_ _19196_/Q _13802_/A _13868_/Y _18732_/Q _13869_/X vssd1 vssd1 vccd1 vccd1
+ _13882_/A sky130_fd_sc_hd__o221a_1
XANTENNA__16986__A0 _17834_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18966__RESET_B hold370/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12821_ _19233_/Q vssd1 vssd1 vccd1 vccd1 _12821_/Y sky130_fd_sc_hd__inv_2
XFILLER_234_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12752_ _19234_/Q vssd1 vssd1 vccd1 vccd1 _12752_/Y sky130_fd_sc_hd__inv_2
X_15540_ _15538_/Y _15539_/X _15512_/X vssd1 vssd1 vccd1 vccd1 _15540_/X sky130_fd_sc_hd__o21a_1
XFILLER_188_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11703_ _11703_/A _18621_/Q vssd1 vssd1 vccd1 vccd1 _11704_/A sky130_fd_sc_hd__and2_1
XFILLER_42_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15471_ _15471_/A _15471_/B vssd1 vssd1 vccd1 vccd1 _15471_/Y sky130_fd_sc_hd__nor2_1
XFILLER_202_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12683_ _18977_/Q _12677_/X hold294/X _12678_/X vssd1 vssd1 vccd1 vccd1 _18977_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_199_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14422_ _18386_/Q _14410_/A _14405_/X _14411_/A vssd1 vssd1 vccd1 vccd1 _18386_/D
+ sky130_fd_sc_hd__a22o_1
X_17210_ _17209_/X _11344_/Y _17459_/S vssd1 vssd1 vccd1 vccd1 _17210_/X sky130_fd_sc_hd__mux2_1
XPHY_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12224__B1 _12223_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11634_ _11622_/A _11622_/B _11632_/Y _11645_/C vssd1 vssd1 vccd1 vccd1 _19552_/D
+ sky130_fd_sc_hd__a211oi_2
XPHY_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18190_ _18198_/CLK _18190_/D vssd1 vssd1 vccd1 vccd1 _18190_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17141_ _15768_/Y _11250_/Y _17546_/S vssd1 vssd1 vccd1 vccd1 _17141_/X sky130_fd_sc_hd__mux2_1
X_14353_ _14353_/A vssd1 vssd1 vccd1 vccd1 _14353_/X sky130_fd_sc_hd__clkbuf_2
XPHY_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11565_ _11565_/A vssd1 vssd1 vccd1 vccd1 _11569_/A sky130_fd_sc_hd__buf_2
XFILLER_11_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13304_ _18861_/Q vssd1 vssd1 vccd1 vccd1 _13433_/B sky130_fd_sc_hd__inv_2
XPHY_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10516_ _10516_/A _10516_/B vssd1 vssd1 vccd1 vccd1 _11649_/B sky130_fd_sc_hd__nand2_1
XFILLER_156_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17072_ _17071_/X _19150_/Q _17548_/S vssd1 vssd1 vccd1 vccd1 _17072_/X sky130_fd_sc_hd__mux2_1
XFILLER_155_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14284_ _18459_/Q _14274_/A _13680_/X _14275_/A vssd1 vssd1 vccd1 vccd1 _18459_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16910__A0 _17473_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11496_ _11486_/A _11486_/B _11528_/A _11494_/Y vssd1 vssd1 vccd1 vccd1 _19606_/D
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__19754__RESET_B repeater196/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13235_ _18883_/Q _13231_/X _18882_/Q _13230_/A vssd1 vssd1 vccd1 vccd1 _18883_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_7_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16023_ _19844_/Q vssd1 vssd1 vccd1 vccd1 _16023_/Y sky130_fd_sc_hd__inv_2
XFILLER_170_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10447_ _19833_/Q _10441_/X _10446_/X _10442_/X vssd1 vssd1 vccd1 vccd1 _19833_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_170_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17466__A1 _13491_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13166_ _13166_/A vssd1 vssd1 vccd1 vccd1 _13166_/Y sky130_fd_sc_hd__inv_2
X_10378_ _10378_/A vssd1 vssd1 vccd1 vccd1 _19856_/D sky130_fd_sc_hd__inv_2
XFILLER_151_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12117_ _19304_/Q _12114_/X _12038_/X _12115_/X vssd1 vssd1 vccd1 vccd1 _19304_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_2_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17974_ _20090_/CLK _17974_/D vssd1 vssd1 vccd1 vccd1 _17974_/Q sky130_fd_sc_hd__dfxtp_1
X_13097_ _19181_/Q vssd1 vssd1 vccd1 vccd1 _13097_/Y sky130_fd_sc_hd__inv_2
X_19713_ _19794_/CLK _19713_/D repeater219/X vssd1 vssd1 vccd1 vccd1 _19713_/Q sky130_fd_sc_hd__dfstp_1
X_16925_ _19669_/Q hold148/X _16950_/S vssd1 vssd1 vccd1 vccd1 _16925_/X sky130_fd_sc_hd__mux2_1
X_12048_ _19334_/Q _12043_/X _11920_/X _12044_/X vssd1 vssd1 vccd1 vccd1 _19334_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_238_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17026__S _17414_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19644_ _19647_/CLK _19644_/D repeater261/X vssd1 vssd1 vccd1 vccd1 _19644_/Q sky130_fd_sc_hd__dfrtp_4
X_16856_ _16855_/X _09865_/A _17524_/S vssd1 vssd1 vccd1 vccd1 _16856_/X sky130_fd_sc_hd__mux2_1
XFILLER_226_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18167__CLK _18169_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_219_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15807_ _18250_/Q vssd1 vssd1 vccd1 vccd1 _15807_/Y sky130_fd_sc_hd__inv_2
X_19575_ _19595_/CLK _19575_/D hold346/A vssd1 vssd1 vccd1 vccd1 _19575_/Q sky130_fd_sc_hd__dfrtp_1
X_16787_ _17473_/A0 _16730_/Y _17473_/S vssd1 vssd1 vccd1 vccd1 _16787_/X sky130_fd_sc_hd__mux2_1
XANTENNA__16865__S _17523_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19412__CLK _19984_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13999_ _18675_/Q vssd1 vssd1 vccd1 vccd1 _14006_/A sky130_fd_sc_hd__inv_2
XFILLER_81_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18526_ _19825_/CLK _18526_/D repeater223/X vssd1 vssd1 vccd1 vccd1 _18526_/Q sky130_fd_sc_hd__dfstp_1
X_15738_ _18667_/Q _18665_/Q vssd1 vssd1 vccd1 vccd1 _15738_/X sky130_fd_sc_hd__or2_1
XFILLER_234_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12463__B1 _12410_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18457_ _18465_/CLK _18457_/D vssd1 vssd1 vccd1 vccd1 _18457_/Q sky130_fd_sc_hd__dfxtp_1
X_15669_ _15669_/A vssd1 vssd1 vccd1 vccd1 _15669_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17408_ _17407_/X _15456_/Y _17518_/S vssd1 vssd1 vccd1 vccd1 _17408_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12215__B1 _12026_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09190_ _20071_/Q vssd1 vssd1 vccd1 vccd1 _09192_/A sky130_fd_sc_hd__inv_2
X_18388_ _19515_/CLK _18388_/D vssd1 vssd1 vccd1 vccd1 _18388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17696__S _17696_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17339_ _16367_/Y _15300_/Y _19498_/Q vssd1 vssd1 vccd1 vccd1 _17339_/X sky130_fd_sc_hd__mux2_1
XANTENNA__19495__RESET_B repeater260/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19009_ _19597_/CLK _19009_/D repeater281/X vssd1 vssd1 vccd1 vccd1 _19009_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__19424__RESET_B repeater271/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11741__A2 _11737_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08974_ _20068_/Q vssd1 vssd1 vccd1 vccd1 _09203_/A sky130_fd_sc_hd__inv_2
XFILLER_29_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09698__B2 _19409_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_217_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_124_HCLK_A clkbuf_4_4_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16775__S _17534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09526_ _09474_/A _19304_/Q _09484_/A _19314_/Q vssd1 vssd1 vccd1 vccd1 _09526_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12454__B1 _12394_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_231_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09457_ _19919_/Q vssd1 vssd1 vccd1 vccd1 _10035_/A sky130_fd_sc_hd__inv_2
XFILLER_196_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09388_ _10088_/A _19376_/Q _10044_/A _09388_/B2 _09387_/X vssd1 vssd1 vccd1 vccd1
+ _09394_/C sky130_fd_sc_hd__o221a_1
XFILLER_184_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_hold319_A HWDATA[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11350_ _19584_/Q _11328_/Y _19594_/Q _11348_/Y _11349_/X vssd1 vssd1 vccd1 vccd1
+ _11350_/X sky130_fd_sc_hd__a221o_1
XANTENNA__16499__A2 _16504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10301_ _18597_/Q _18596_/Q _15605_/A vssd1 vssd1 vccd1 vccd1 _15612_/A sky130_fd_sc_hd__or3_1
XFILLER_153_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17791__S1 _19646_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11281_ _19012_/Q vssd1 vssd1 vccd1 vccd1 _16615_/A sky130_fd_sc_hd__inv_2
XANTENNA__19165__RESET_B hold370/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14324__A hold325/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13020_ _18923_/Q _13023_/A _13017_/A _12958_/X vssd1 vssd1 vccd1 vccd1 _18923_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_4_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10232_ _19833_/Q _19660_/Q _19833_/Q _19660_/Q vssd1 vssd1 vccd1 vccd1 _10232_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_133_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10163_ _19889_/Q _10155_/A _09105_/X _10156_/A vssd1 vssd1 vccd1 vccd1 _19889_/D
+ sky130_fd_sc_hd__a22o_1
X_10094_ _10094_/A vssd1 vssd1 vccd1 vccd1 _10094_/Y sky130_fd_sc_hd__inv_2
X_14971_ _18069_/Q _14964_/X _14812_/X _14966_/X vssd1 vssd1 vccd1 vccd1 _18069_/D
+ sky130_fd_sc_hd__a22o_1
X_16710_ _19053_/Q vssd1 vssd1 vccd1 vccd1 _16710_/Y sky130_fd_sc_hd__inv_2
XFILLER_120_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13922_ _18729_/Q _13921_/Y _13907_/X _13829_/B vssd1 vssd1 vccd1 vccd1 _18729_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12693__B1 hold239/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17690_ _15472_/X _19445_/Q _17696_/S vssd1 vssd1 vccd1 vccd1 _18562_/D sky130_fd_sc_hd__mux2_1
XFILLER_208_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16641_ _16572_/X _16641_/B _16641_/C vssd1 vssd1 vccd1 vccd1 _16641_/Y sky130_fd_sc_hd__nand3b_4
X_13853_ _13852_/Y _18713_/Q _19202_/Q _13950_/A vssd1 vssd1 vccd1 vccd1 _13853_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_142_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12804_ _18826_/Q vssd1 vssd1 vccd1 vccd1 _13549_/A sky130_fd_sc_hd__inv_6
XFILLER_16_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19360_ _19970_/CLK _19360_/D repeater249/X vssd1 vssd1 vccd1 vccd1 _19360_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__12445__B1 _12375_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16572_ _16682_/A vssd1 vssd1 vccd1 vccd1 _16572_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_leaf_46_HCLK_A clkbuf_opt_2_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10996_ _10996_/A _10996_/B vssd1 vssd1 vccd1 vccd1 _10996_/X sky130_fd_sc_hd__and2_1
X_13784_ _18728_/Q vssd1 vssd1 vccd1 vccd1 _13914_/B sky130_fd_sc_hd__inv_2
XFILLER_204_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18311_ _18431_/CLK _18311_/D vssd1 vssd1 vccd1 vccd1 _18311_/Q sky130_fd_sc_hd__dfxtp_1
X_15523_ _18575_/Q _15523_/B vssd1 vssd1 vccd1 vccd1 _15537_/B sky130_fd_sc_hd__or2_1
X_12735_ _18813_/Q vssd1 vssd1 vccd1 vccd1 _13537_/B sky130_fd_sc_hd__inv_2
X_19291_ _19293_/CLK _19291_/D repeater187/X vssd1 vssd1 vccd1 vccd1 _19291_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_15_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_repeater176_A _17524_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18242_ _19847_/CLK _18242_/D vssd1 vssd1 vccd1 vccd1 _18242_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12666_ _18990_/Q _12661_/X hold291/X _12664_/X vssd1 vssd1 vccd1 vccd1 _18990_/D
+ sky130_fd_sc_hd__a22o_1
X_15454_ _18558_/Q _15453_/A _15452_/Y _15453_/Y vssd1 vssd1 vccd1 vccd1 _15455_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_188_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11617_ _11617_/A vssd1 vssd1 vccd1 vccd1 _11645_/C sky130_fd_sc_hd__buf_2
X_14405_ _14405_/A vssd1 vssd1 vccd1 vccd1 _14405_/X sky130_fd_sc_hd__buf_2
XANTENNA__17136__A0 _17473_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18173_ _18216_/CLK _18173_/D vssd1 vssd1 vccd1 vccd1 _18173_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15385_ _15211_/Y _15217_/A _15384_/A vssd1 vssd1 vccd1 vccd1 _18511_/D sky130_fd_sc_hd__o21a_1
X_12597_ _19032_/Q _12590_/X _12596_/X _12591_/X vssd1 vssd1 vccd1 vccd1 _19032_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_184_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17124_ _16484_/X _10242_/Y _17566_/S vssd1 vssd1 vccd1 vccd1 _17124_/X sky130_fd_sc_hd__mux2_1
XPHY_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14336_ _14337_/A vssd1 vssd1 vccd1 vccd1 _14336_/X sky130_fd_sc_hd__clkbuf_2
X_11548_ _11548_/A _11548_/B _11639_/C vssd1 vssd1 vccd1 vccd1 _11619_/C sky130_fd_sc_hd__or3_1
XFILLER_237_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17782__S1 _19646_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14267_ _18467_/Q _14259_/A _12731_/X _14260_/A vssd1 vssd1 vccd1 vccd1 _18467_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_116_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17055_ _16667_/Y _17055_/A1 _17541_/S vssd1 vssd1 vccd1 vccd1 _17055_/X sky130_fd_sc_hd__mux2_1
XANTENNA__15162__A2 _15158_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11479_ _11479_/A _11508_/A vssd1 vssd1 vccd1 vccd1 _11480_/B sky130_fd_sc_hd__or2_2
XANTENNA__14234__A _14236_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13218_ _18531_/Q _13218_/B vssd1 vssd1 vccd1 vccd1 _13219_/B sky130_fd_sc_hd__or2_1
X_16006_ _15846_/X _15979_/X _15859_/X _15989_/X _16005_/X vssd1 vssd1 vccd1 vccd1
+ _16006_/Y sky130_fd_sc_hd__o221ai_4
XANTENNA__14370__B1 _14351_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14198_ _14194_/Y _18683_/Q _14195_/Y _18678_/Q _14197_/X vssd1 vssd1 vccd1 vccd1
+ _14219_/B sky130_fd_sc_hd__o221a_1
XFILLER_97_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13149_ _19167_/Q vssd1 vssd1 vccd1 vccd1 _13149_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18757__SET_B repeater196/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18888__RESET_B repeater188/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17957_ _20077_/CLK _17957_/D vssd1 vssd1 vccd1 vccd1 _17957_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18817__RESET_B repeater231/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16908_ _16645_/Y _19284_/Q _17541_/S vssd1 vssd1 vccd1 vccd1 _16908_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17888_ _16038_/Y _16039_/Y _16040_/Y _16041_/Y _17908_/S0 _18759_/Q vssd1 vssd1
+ vccd1 vccd1 _17888_/X sky130_fd_sc_hd__mux4_2
XFILLER_238_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19627_ _19873_/CLK _19627_/D repeater261/X vssd1 vssd1 vccd1 vccd1 _19627_/Q sky130_fd_sc_hd__dfrtp_2
X_16839_ _16838_/X _15690_/Y _17318_/S vssd1 vssd1 vccd1 vccd1 _16839_/X sky130_fd_sc_hd__mux2_1
XFILLER_81_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19558_ _19582_/CLK _19558_/D hold348/A vssd1 vssd1 vccd1 vccd1 _19558_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_241_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09311_ _18661_/Q vssd1 vssd1 vccd1 vccd1 _09311_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18509_ _19544_/CLK _18509_/D repeater222/X vssd1 vssd1 vccd1 vccd1 _18509_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_178_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19489_ _19515_/CLK hold135/X repeater259/X vssd1 vssd1 vccd1 vccd1 _19489_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_61_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09242_ _09242_/A _09242_/B _18651_/D _09241_/X vssd1 vssd1 vccd1 vccd1 _10759_/B
+ sky130_fd_sc_hd__or4b_4
X_09173_ _20078_/Q vssd1 vssd1 vccd1 vccd1 _14707_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__17127__A0 _17486_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19605__RESET_B hold359/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15689__B1 _15673_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17773__S1 _19646_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15153__A2 _15146_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14361__B1 hold324/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_227_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08957_ _19864_/Q vssd1 vssd1 vccd1 vccd1 _10330_/A sky130_fd_sc_hd__inv_2
XFILLER_88_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12599__A _14277_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18558__RESET_B repeater193/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12675__B1 hold296/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold269_A HWDATA[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10850_ _19712_/Q _10843_/X _10421_/X _10845_/X vssd1 vssd1 vccd1 vccd1 _19712_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_112_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09509_ _19301_/Q vssd1 vssd1 vccd1 vccd1 _09509_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16169__A1 _11023_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17366__A0 _15768_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10781_ _17630_/X _10773_/A _19743_/Q _10774_/A vssd1 vssd1 vccd1 vccd1 _19743_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_12_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12520_ _12529_/A vssd1 vssd1 vccd1 vccd1 _12520_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_201_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15916__A1 _17545_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_234_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15916__B2 _15915_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12451_ _12458_/A vssd1 vssd1 vccd1 vccd1 _12451_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_200_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19346__RESET_B repeater245/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11402_ _19562_/Q vssd1 vssd1 vccd1 vccd1 _11575_/A sky130_fd_sc_hd__inv_2
XFILLER_21_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15170_ _15171_/A vssd1 vssd1 vccd1 vccd1 _15170_/X sky130_fd_sc_hd__clkbuf_2
X_12382_ hold289/X vssd1 vssd1 vccd1 vccd1 _12382_/X sky130_fd_sc_hd__buf_2
XFILLER_126_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14121_ _18691_/Q _14120_/Y _14116_/X _14121_/C1 vssd1 vssd1 vccd1 vccd1 _18691_/D
+ sky130_fd_sc_hd__o211a_1
X_11333_ _18977_/Q vssd1 vssd1 vccd1 vccd1 _11333_/Y sky130_fd_sc_hd__inv_2
XFILLER_192_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14052_ _19079_/Q _14020_/A _14050_/Y _18678_/Q _14051_/X vssd1 vssd1 vccd1 vccd1
+ _14064_/A sky130_fd_sc_hd__a221o_1
XFILLER_113_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11264_ _18998_/Q vssd1 vssd1 vccd1 vccd1 _11264_/Y sky130_fd_sc_hd__inv_2
XFILLER_122_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13003_ _13003_/A _13017_/A vssd1 vssd1 vccd1 vccd1 _13004_/B sky130_fd_sc_hd__or2_1
X_10215_ _10213_/Y _19664_/Q _19837_/Q _10964_/A vssd1 vssd1 vccd1 vccd1 _10215_/X
+ sky130_fd_sc_hd__o22a_1
X_18860_ _18866_/CLK _18860_/D repeater232/X vssd1 vssd1 vccd1 vccd1 _18860_/Q sky130_fd_sc_hd__dfrtp_1
X_11195_ _17717_/X _11191_/X _19614_/Q _11192_/X vssd1 vssd1 vccd1 vccd1 _19614_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_239_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17811_ _18188_/Q _18180_/Q _18172_/Q _18156_/Q _17918_/S0 _18750_/Q vssd1 vssd1
+ vccd1 vccd1 _17811_/X sky130_fd_sc_hd__mux4_1
X_10146_ hold322/X vssd1 vssd1 vccd1 vccd1 hold321/A sky130_fd_sc_hd__clkbuf_2
XFILLER_79_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18791_ _19647_/CLK _18791_/D repeater261/X vssd1 vssd1 vccd1 vccd1 _18791_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18910__RESET_B repeater188/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17742_ _15367_/X _19703_/Q _18508_/D vssd1 vssd1 vccd1 vccd1 _17742_/X sky130_fd_sc_hd__mux2_1
XFILLER_153_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10077_ _10077_/A vssd1 vssd1 vccd1 vccd1 _10077_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12666__B1 hold291/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14954_ _14954_/A vssd1 vssd1 vccd1 vccd1 _14954_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__12302__A _14279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13905_ _13832_/A _13832_/B _13833_/Y _13970_/C vssd1 vssd1 vccd1 vccd1 _18734_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_235_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17673_ _15543_/X _19462_/Q _17683_/S vssd1 vssd1 vccd1 vccd1 _18579_/D sky130_fd_sc_hd__mux2_1
X_14885_ _14885_/A vssd1 vssd1 vccd1 vccd1 _14885_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_47_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17304__S _17518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19412_ _19984_/CLK _19412_/D repeater244/X vssd1 vssd1 vccd1 vccd1 _19412_/Q sky130_fd_sc_hd__dfrtp_4
X_16624_ _19045_/Q _16673_/B vssd1 vssd1 vccd1 vccd1 _16624_/Y sky130_fd_sc_hd__nand2_1
XFILLER_90_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12418__B1 hold256/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13836_ _19212_/Q _18723_/Q _13835_/Y _13910_/C vssd1 vssd1 vccd1 vccd1 _13850_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_223_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19343_ _19952_/CLK _19343_/D repeater244/X vssd1 vssd1 vccd1 vccd1 _19343_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17357__A0 _15963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16555_ _16555_/A vssd1 vssd1 vccd1 vccd1 _16555_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_31_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10979_ _10979_/A vssd1 vssd1 vccd1 vccd1 _10980_/B sky130_fd_sc_hd__inv_2
XFILLER_90_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13767_ _13775_/S vssd1 vssd1 vccd1 vccd1 _13772_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_15_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15506_ _18570_/Q _15498_/A _18571_/Q vssd1 vssd1 vccd1 vccd1 _15506_/X sky130_fd_sc_hd__o21a_1
XFILLER_231_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12718_ _14808_/A _12709_/X _12717_/X _12711_/X vssd1 vssd1 vccd1 vccd1 _18957_/D
+ sky130_fd_sc_hd__a22o_1
X_19274_ _19282_/CLK _19274_/D repeater216/X vssd1 vssd1 vccd1 vccd1 _19274_/Q sky130_fd_sc_hd__dfrtp_1
X_16486_ _19034_/Q vssd1 vssd1 vccd1 vccd1 _16486_/Y sky130_fd_sc_hd__inv_2
XFILLER_188_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13698_ _13700_/A _13506_/A _14668_/B vssd1 vssd1 vccd1 vccd1 _13698_/X sky130_fd_sc_hd__o21a_1
XFILLER_30_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17109__A0 _17486_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18225_ _20077_/CLK _18225_/D vssd1 vssd1 vccd1 vccd1 _18225_/Q sky130_fd_sc_hd__dfxtp_1
X_15437_ _19773_/Q _15437_/B vssd1 vssd1 vccd1 vccd1 _15437_/X sky130_fd_sc_hd__or2_1
XFILLER_248_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19087__RESET_B hold351/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12649_ _18999_/Q _12643_/X _12596_/X _12644_/X vssd1 vssd1 vccd1 vccd1 _18999_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_248_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18156_ _20123_/CLK _18156_/D vssd1 vssd1 vccd1 vccd1 _18156_/Q sky130_fd_sc_hd__dfxtp_1
X_15368_ _19784_/Q _10644_/B _10645_/B vssd1 vssd1 vccd1 vccd1 _15368_/X sky130_fd_sc_hd__a21bo_1
XFILLER_156_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17107_ _16546_/Y _20105_/Q _17535_/S vssd1 vssd1 vccd1 vccd1 _17107_/X sky130_fd_sc_hd__mux2_1
X_14319_ _14319_/A vssd1 vssd1 vccd1 vccd1 _14320_/A sky130_fd_sc_hd__inv_2
Xhold305 hold305/A vssd1 vssd1 vccd1 vccd1 hold305/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold316 HWDATA[21] vssd1 vssd1 vccd1 vccd1 input51/A sky130_fd_sc_hd__dlygate4sd3_1
X_18087_ _20077_/CLK _18087_/D vssd1 vssd1 vccd1 vccd1 _18087_/Q sky130_fd_sc_hd__dfxtp_1
X_15299_ _15334_/B _18513_/Q vssd1 vssd1 vccd1 vccd1 _15735_/B sky130_fd_sc_hd__or2_2
Xhold327 HWDATA[4] vssd1 vssd1 vccd1 vccd1 input64/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13146__A1 _19170_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold338 input78/X vssd1 vssd1 vccd1 vccd1 hold338/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14343__B1 _14326_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17038_ _16624_/Y _15660_/Y _17318_/S vssd1 vssd1 vccd1 vccd1 _17038_/X sky130_fd_sc_hd__mux2_2
Xhold349 hold366/X vssd1 vssd1 vccd1 vccd1 hold365/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09058__A hold233/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09860_ _09860_/A _09981_/A vssd1 vssd1 vccd1 vccd1 _09861_/B sky130_fd_sc_hd__or2_2
XANTENNA__19750__CLK _19900_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09791_ _09791_/A _09800_/A vssd1 vssd1 vccd1 vccd1 _09792_/B sky130_fd_sc_hd__or2_2
X_18989_ _19608_/CLK _18989_/D hold273/X vssd1 vssd1 vccd1 vccd1 _18989_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_97_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12657__B1 _12541_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_227_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12212__A _12228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater155 _17517_/S vssd1 vssd1 vccd1 vccd1 _17413_/S sky130_fd_sc_hd__buf_8
Xrepeater166 _17543_/S vssd1 vssd1 vccd1 vccd1 _17534_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_238_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrepeater177 _17518_/S vssd1 vssd1 vccd1 vccd1 _17524_/S sky130_fd_sc_hd__buf_8
XPHY_4309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater188 hold373/A vssd1 vssd1 vccd1 vccd1 repeater188/X sky130_fd_sc_hd__buf_8
XFILLER_27_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrepeater199 repeater200/X vssd1 vssd1 vccd1 vccd1 repeater199/X sky130_fd_sc_hd__buf_6
XFILLER_226_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17214__S _17524_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10683__A2 _10676_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12409__B1 _12408_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_92_HCLK_A clkbuf_4_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_179_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09225_ _18644_/Q vssd1 vssd1 vccd1 vccd1 _15709_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_210_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09156_ _09156_/A _09156_/B vssd1 vssd1 vccd1 vccd1 _09156_/Y sky130_fd_sc_hd__nor2_1
XFILLER_181_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09087_ _09087_/A vssd1 vssd1 vccd1 vccd1 _09087_/X sky130_fd_sc_hd__buf_1
XFILLER_174_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16323__B2 _15999_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18848__CLK _18866_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10000_ _09850_/A _10000_/A2 _09998_/Y _09990_/X vssd1 vssd1 vccd1 vccd1 _19941_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_67_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09989_ _09857_/B _09989_/A2 _19948_/Q _09988_/Y _09950_/X vssd1 vssd1 vccd1 vccd1
+ _19948_/D sky130_fd_sc_hd__o221a_1
XFILLER_237_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12648__B1 hold259/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_217_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10659__C1 _10658_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11951_ _19391_/Q _11948_/X _09033_/X _11949_/X vssd1 vssd1 vccd1 vccd1 _19391_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_29_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17124__S _17566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10902_ _19686_/Q _10894_/A _10868_/X _10895_/A vssd1 vssd1 vccd1 vccd1 _19686_/D
+ sky130_fd_sc_hd__a22o_1
X_11882_ _19429_/Q _11875_/X _09025_/X _11878_/X vssd1 vssd1 vccd1 vccd1 _19429_/D
+ sky130_fd_sc_hd__a22o_1
X_14670_ _14670_/A vssd1 vssd1 vccd1 vccd1 _14671_/A sky130_fd_sc_hd__inv_2
XFILLER_233_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10833_ _10833_/A vssd1 vssd1 vccd1 vccd1 _19720_/D sky130_fd_sc_hd__inv_2
X_13621_ _13613_/Y _17762_/S _13617_/A _13620_/Y vssd1 vssd1 vccd1 vccd1 _13621_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_32_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16963__S _17529_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_241_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16340_ _18344_/Q vssd1 vssd1 vccd1 vccd1 _16340_/Y sky130_fd_sc_hd__inv_2
X_13552_ _13552_/A _13569_/A vssd1 vssd1 vccd1 vccd1 _13553_/B sky130_fd_sc_hd__or2_2
X_10764_ _19752_/Q vssd1 vssd1 vccd1 vccd1 _10764_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12503_ _19084_/Q _12498_/X _12396_/X _12499_/X vssd1 vssd1 vccd1 vccd1 _19084_/D
+ sky130_fd_sc_hd__a22o_1
X_13483_ _13483_/A _13483_/B _13483_/C vssd1 vssd1 vccd1 vccd1 _13486_/A sky130_fd_sc_hd__or3_4
X_16271_ _19638_/Q _16095_/Y _16269_/X _16270_/X _16172_/Y vssd1 vssd1 vccd1 vccd1
+ _16271_/Y sky130_fd_sc_hd__o221ai_4
XANTENNA__19623__CLK _19920_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10695_ _10446_/A _17749_/X _17749_/S _19780_/Q _10694_/Y vssd1 vssd1 vccd1 vccd1
+ _19780_/D sky130_fd_sc_hd__a32o_1
XFILLER_185_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16562__B2 _16506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18010_ _18954_/CLK _18010_/D vssd1 vssd1 vccd1 vccd1 _18010_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_201_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12434_ _19127_/Q _12400_/A _12238_/X _12402_/A vssd1 vssd1 vccd1 vccd1 _19127_/D
+ sky130_fd_sc_hd__a22o_1
X_15222_ _15222_/A _15232_/B vssd1 vssd1 vccd1 vccd1 _15222_/Y sky130_fd_sc_hd__nor2_1
XFILLER_138_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20085__RESET_B repeater204/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12365_ _19162_/Q _12361_/X _12232_/X _12362_/X vssd1 vssd1 vccd1 vccd1 _19162_/D
+ sky130_fd_sc_hd__a22o_1
X_15153_ _17956_/Q _15146_/X _14709_/A _15148_/X vssd1 vssd1 vccd1 vccd1 _17956_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_181_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14104_ _14104_/A vssd1 vssd1 vccd1 vccd1 _14104_/Y sky130_fd_sc_hd__clkinv_1
XANTENNA__14325__B1 hold324/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11316_ _18962_/Q vssd1 vssd1 vccd1 vccd1 _11316_/Y sky130_fd_sc_hd__inv_2
XFILLER_153_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15084_ _15084_/A vssd1 vssd1 vccd1 vccd1 _15085_/A sky130_fd_sc_hd__inv_2
X_19961_ _19964_/CLK _19961_/D hold371/X vssd1 vssd1 vccd1 vccd1 _19961_/Q sky130_fd_sc_hd__dfrtp_1
X_12296_ _14273_/A vssd1 vssd1 vccd1 vccd1 _12296_/X sky130_fd_sc_hd__buf_2
X_14035_ _19070_/Q vssd1 vssd1 vccd1 vccd1 _14035_/Y sky130_fd_sc_hd__inv_2
X_18912_ _19222_/CLK _18912_/D repeater188/X vssd1 vssd1 vccd1 vccd1 _18912_/Q sky130_fd_sc_hd__dfrtp_1
X_11247_ _11468_/A _19002_/Q _11475_/A _19009_/Q _11246_/X vssd1 vssd1 vccd1 vccd1
+ _11248_/D sky130_fd_sc_hd__o221a_1
X_19892_ _20055_/CLK _19892_/D repeater205/X vssd1 vssd1 vccd1 vccd1 _19892_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_68_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18843_ _18866_/CLK _18843_/D repeater233/X vssd1 vssd1 vccd1 vccd1 _18843_/Q sky130_fd_sc_hd__dfrtp_1
X_11178_ _11192_/A vssd1 vssd1 vccd1 vccd1 _11178_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_79_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10129_ _15447_/B vssd1 vssd1 vccd1 vccd1 _10130_/B sky130_fd_sc_hd__inv_2
XFILLER_94_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13128__A _19173_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12639__B1 hold233/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18774_ _19855_/CLK _18774_/D repeater265/X vssd1 vssd1 vccd1 vccd1 _18774_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12032__A _12032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15986_ _19816_/Q vssd1 vssd1 vccd1 vccd1 _15986_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17725_ _19675_/Q _19688_/Q _18510_/Q vssd1 vssd1 vccd1 vccd1 _17725_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14937_ _18090_/Q _14922_/A _14868_/X _14923_/A vssd1 vssd1 vccd1 vccd1 _18090_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_75_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17034__S _17487_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17656_ _15610_/Y _19033_/Q _17664_/S vssd1 vssd1 vccd1 vccd1 _18596_/D sky130_fd_sc_hd__mux2_1
XANTENNA__19950__RESET_B hold371/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14868_ _20074_/Q vssd1 vssd1 vccd1 vccd1 _14868_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_235_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16250__B1 _16237_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16607_ _16572_/X _16607_/B _16607_/C vssd1 vssd1 vccd1 vccd1 _16607_/Y sky130_fd_sc_hd__nand3b_4
X_13819_ _13910_/D _13819_/B vssd1 vssd1 vccd1 vccd1 _13935_/A sky130_fd_sc_hd__or2_1
X_17587_ _15363_/X _19716_/Q _17600_/S vssd1 vssd1 vccd1 vccd1 _17587_/X sky130_fd_sc_hd__mux2_1
XANTENNA__16873__S _17543_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19268__RESET_B repeater212/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14799_ _19850_/Q vssd1 vssd1 vccd1 vccd1 _15034_/B sky130_fd_sc_hd__buf_1
X_19326_ _19971_/CLK _19326_/D repeater241/X vssd1 vssd1 vccd1 vccd1 _19326_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_177_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16538_ _17120_/X _16508_/X _17113_/X _15908_/X _16537_/X vssd1 vssd1 vccd1 vccd1
+ _16538_/X sky130_fd_sc_hd__o221a_1
XFILLER_188_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19257_ _19324_/CLK _19257_/D repeater237/X vssd1 vssd1 vccd1 vccd1 _19257_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_31_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17750__A0 _15735_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16469_ _16469_/A _16469_/B vssd1 vssd1 vccd1 vccd1 _16469_/Y sky130_fd_sc_hd__nor2_1
X_09010_ _19508_/Q _19507_/Q _09010_/C _09010_/D vssd1 vssd1 vccd1 vccd1 _11832_/C
+ sky130_fd_sc_hd__or4_4
X_18208_ _18333_/CLK _18208_/D vssd1 vssd1 vccd1 vccd1 _18208_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14564__B1 _14509_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19188_ _19293_/CLK _19188_/D repeater187/X vssd1 vssd1 vccd1 vccd1 _19188_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_163_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18139_ _18142_/CLK _18139_/D vssd1 vssd1 vccd1 vccd1 _18139_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold135 hold135/A vssd1 vssd1 vccd1 vccd1 hold135/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold146 HADDR[15] vssd1 vssd1 vccd1 vccd1 input7/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold157 HADDR[14] vssd1 vssd1 vccd1 vccd1 input6/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16621__B _16621_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20101_ _20122_/CLK _20101_/D repeater234/X vssd1 vssd1 vccd1 vccd1 _20101_/Q sky130_fd_sc_hd__dfrtp_2
Xhold168 input2/X vssd1 vssd1 vccd1 vccd1 hold168/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold179 hold179/A vssd1 vssd1 vccd1 vccd1 hold179/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17209__S _17546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09912_ _19352_/Q vssd1 vssd1 vccd1 vccd1 _09912_/Y sky130_fd_sc_hd__inv_2
XFILLER_160_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20032_ _20032_/CLK _20032_/D repeater240/X vssd1 vssd1 vccd1 vccd1 _20032_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_101_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09843_ _19943_/Q vssd1 vssd1 vccd1 vccd1 _09852_/A sky130_fd_sc_hd__inv_2
XFILLER_98_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17900__S1 _19632_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09774_ _09748_/A _09748_/B _09767_/X _09772_/Y vssd1 vssd1 vccd1 vccd1 _19992_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_37_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_61_HCLK clkbuf_opt_3_HCLK/A vssd1 vssd1 vccd1 vccd1 _19937_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_39_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19620__RESET_B repeater230/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16783__S _17512_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold134_A HADDR[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14555__B1 hold334/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09208_ _09205_/A _09198_/X _09205_/Y vssd1 vssd1 vccd1 vccd1 _20067_/D sky130_fd_sc_hd__a21oi_1
X_10480_ _17704_/X _10471_/A _19815_/Q _10472_/A vssd1 vssd1 vccd1 vccd1 _19815_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_183_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09139_ _09139_/A _09139_/B vssd1 vssd1 vccd1 vccd1 _09139_/Y sky130_fd_sc_hd__nor2_1
XFILLER_185_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14307__B1 _14277_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09982__B1 _09968_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12150_ _12150_/A vssd1 vssd1 vccd1 vccd1 _12150_/X sky130_fd_sc_hd__clkbuf_2
X_11101_ _15094_/A _10400_/B _19851_/Q _10400_/B vssd1 vssd1 vccd1 vccd1 _11101_/X
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__17119__S _17512_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12081_ _19321_/Q _12068_/X _12080_/X _12072_/X vssd1 vssd1 vccd1 vccd1 _19321_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_151_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18502__RESET_B repeater219/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11032_ _11022_/X _11026_/Y _17753_/S _11030_/X _11031_/X vssd1 vssd1 vccd1 vccd1
+ _11032_/X sky130_fd_sc_hd__o221a_1
XANTENNA__16958__S _17541_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15840_ _15840_/A vssd1 vssd1 vccd1 vccd1 _15840_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__18050__CLK _19851_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16480__B1 _16990_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15771_ _16721_/B vssd1 vssd1 vccd1 vccd1 _17522_/S sky130_fd_sc_hd__clkinv_8
XFILLER_94_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12983_ _12983_/A vssd1 vssd1 vccd1 vccd1 _12983_/Y sky130_fd_sc_hd__inv_2
XFILLER_91_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17510_ _17509_/X _10293_/Y _17548_/S vssd1 vssd1 vccd1 vccd1 _17510_/X sky130_fd_sc_hd__mux2_1
X_14722_ _18215_/Q _14717_/X _14606_/X _14719_/X vssd1 vssd1 vccd1 vccd1 _18215_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_94_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18490_ _19720_/CLK _18490_/D repeater201/X vssd1 vssd1 vccd1 vccd1 _18490_/Q sky130_fd_sc_hd__dfrtp_1
X_11934_ _11841_/X _19398_/Q _11934_/S vssd1 vssd1 vccd1 vccd1 _19398_/D sky130_fd_sc_hd__mux2_1
XFILLER_245_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17441_ _17486_/A0 _16047_/Y _17517_/S vssd1 vssd1 vccd1 vccd1 _17441_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14653_ _18250_/Q _14644_/A _14626_/X _14645_/A vssd1 vssd1 vccd1 vccd1 _18250_/D
+ sky130_fd_sc_hd__a22o_1
X_11865_ _13641_/A _11853_/A _11856_/A _11869_/B vssd1 vssd1 vccd1 vccd1 _11865_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__19361__RESET_B hold370/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output106_A _16327_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13604_ _13604_/A vssd1 vssd1 vccd1 vccd1 _13604_/Y sky130_fd_sc_hd__inv_2
XFILLER_159_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10816_ _17620_/X _10809_/A _19727_/Q _10810_/A vssd1 vssd1 vccd1 vccd1 _19727_/D
+ sky130_fd_sc_hd__a22o_1
X_17372_ _17371_/X _16294_/Y _17567_/S vssd1 vssd1 vccd1 vccd1 _17372_/X sky130_fd_sc_hd__mux2_1
XANTENNA__14794__B1 _14793_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14584_ _18291_/Q _14573_/A _14567_/X _14574_/A vssd1 vssd1 vccd1 vccd1 _18291_/D
+ sky130_fd_sc_hd__a22o_1
X_11796_ _19464_/Q _11793_/X _09033_/X _11794_/X vssd1 vssd1 vccd1 vccd1 _19464_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19111_ _19115_/CLK _19111_/D hold353/X vssd1 vssd1 vccd1 vccd1 _19111_/Q sky130_fd_sc_hd__dfrtp_2
X_16323_ _17368_/X _15904_/A _17373_/X _15999_/X vssd1 vssd1 vccd1 vccd1 _16323_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_185_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13535_ _13535_/A _13601_/A vssd1 vssd1 vccd1 vccd1 _13536_/B sky130_fd_sc_hd__or2_1
X_10747_ _19760_/Q _10741_/X _10418_/X _10743_/X vssd1 vssd1 vccd1 vccd1 _19760_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_13_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_repeater256_A repeater260/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19042_ _19566_/CLK _19042_/D repeater255/X vssd1 vssd1 vccd1 vccd1 _19042_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__10280__B1 _19646_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16254_ _18031_/Q vssd1 vssd1 vccd1 vccd1 _16254_/Y sky130_fd_sc_hd__inv_2
X_13466_ _13466_/A _13466_/B vssd1 vssd1 vccd1 vccd1 _13476_/A sky130_fd_sc_hd__or2_1
X_10678_ _17739_/X _10676_/X _19786_/Q _10677_/X vssd1 vssd1 vccd1 vccd1 _19786_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_185_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15205_ _19724_/Q vssd1 vssd1 vccd1 vccd1 _15205_/Y sky130_fd_sc_hd__inv_2
X_12417_ _19140_/Q _12412_/X hold281/X _12414_/X vssd1 vssd1 vccd1 vccd1 _19140_/D
+ sky130_fd_sc_hd__a22o_1
X_16185_ _18134_/Q vssd1 vssd1 vccd1 vccd1 _16185_/Y sky130_fd_sc_hd__inv_2
X_13397_ _20094_/Q vssd1 vssd1 vccd1 vccd1 _13397_/Y sky130_fd_sc_hd__clkinv_1
XFILLER_154_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15136_ _15136_/A vssd1 vssd1 vccd1 vccd1 _15136_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__09973__B1 _09968_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12348_ hold257/X vssd1 vssd1 vccd1 vccd1 hold256/A sky130_fd_sc_hd__buf_4
XFILLER_245_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15338__A _15364_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17029__S _17490_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15067_ _18012_/Q _15060_/A _14814_/A _15061_/A vssd1 vssd1 vccd1 vccd1 _18012_/D
+ sky130_fd_sc_hd__a22o_1
X_12279_ _19213_/Q _12276_/X _12098_/X _12277_/X vssd1 vssd1 vccd1 vccd1 _19213_/D
+ sky130_fd_sc_hd__a22o_1
X_19944_ _19976_/CLK _19944_/D repeater244/X vssd1 vssd1 vccd1 vccd1 _19944_/Q sky130_fd_sc_hd__dfrtp_1
X_14018_ _14018_/A _14018_/B vssd1 vssd1 vccd1 vccd1 _14123_/A sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_84_HCLK clkbuf_4_13_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19320_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__16868__S _17547_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19875_ _20059_/CLK _19875_/D repeater198/X vssd1 vssd1 vccd1 vccd1 _19875_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_67_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18826_ _19255_/CLK _18826_/D repeater217/X vssd1 vssd1 vccd1 vccd1 _18826_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__17894__S0 _19633_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_244_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18757_ _19900_/CLK _18757_/D repeater196/X vssd1 vssd1 vccd1 vccd1 _18757_/Q sky130_fd_sc_hd__dfstp_2
X_15969_ _10834_/Y _15854_/X _15968_/Y _15867_/B vssd1 vssd1 vccd1 vccd1 _15969_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_48_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19449__RESET_B repeater271/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_224_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17708_ _15432_/X _19769_/Q _18546_/D vssd1 vssd1 vccd1 vccd1 _17708_/X sky130_fd_sc_hd__mux2_1
X_09490_ _09490_/A _09490_/B vssd1 vssd1 vccd1 vccd1 _09574_/A sky130_fd_sc_hd__or2_1
XFILLER_236_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18688_ _18701_/CLK _18688_/D hold359/X vssd1 vssd1 vccd1 vccd1 _18688_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_64_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09071__A hold239/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17639_ _15684_/X _19050_/Q _17655_/S vssd1 vssd1 vccd1 vccd1 _18613_/D sky130_fd_sc_hd__mux2_1
XFILLER_91_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19309_ _20120_/CLK _19309_/D repeater238/X vssd1 vssd1 vccd1 vccd1 _19309_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_32_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14417__A hold331/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18073__CLK _18169_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_235_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16778__S _17474_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20015_ _20032_/CLK _20015_/D repeater240/X vssd1 vssd1 vccd1 vccd1 _20015_/Q sky130_fd_sc_hd__dfrtp_1
X_09826_ _19960_/Q vssd1 vssd1 vccd1 vccd1 _09868_/A sky130_fd_sc_hd__inv_2
XFILLER_246_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17885__S0 _17908_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16462__B1 _17086_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09757_ _09757_/A _09757_/B vssd1 vssd1 vccd1 vccd1 _09758_/C sky130_fd_sc_hd__nor2_1
XANTENNA__19801__RESET_B repeater222/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12400__A _12400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09688_ _19998_/Q _09684_/Y _19982_/Q _09685_/Y _09687_/X vssd1 vssd1 vccd1 vccd1
+ _09689_/D sky130_fd_sc_hd__o221a_1
XPHY_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17402__S _17566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11650_ _15270_/B _11650_/B _15271_/C vssd1 vssd1 vccd1 vccd1 _11672_/B sky130_fd_sc_hd__or3_4
XFILLER_187_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14776__B1 _14751_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10601_ _15334_/C _10938_/B _10584_/X _10598_/Y _10600_/Y vssd1 vssd1 vccd1 vccd1
+ _10601_/X sky130_fd_sc_hd__a41o_1
XPHY_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11581_ _11581_/A _11581_/B vssd1 vssd1 vccd1 vccd1 _11600_/A sky130_fd_sc_hd__or2_1
XANTENNA__12251__A1 _10954_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10532_ _10736_/B _10537_/A _10532_/C _10531_/X vssd1 vssd1 vccd1 vccd1 _11672_/C
+ sky130_fd_sc_hd__or4b_4
X_13320_ _18839_/Q vssd1 vssd1 vccd1 vccd1 _13322_/B sky130_fd_sc_hd__inv_4
XFILLER_155_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14528__B1 _14474_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18754__RESET_B repeater195/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10463_ _19825_/Q _10462_/A _10461_/Y _10462_/Y _18548_/Q vssd1 vssd1 vccd1 vccd1
+ _19825_/D sky130_fd_sc_hd__a221o_1
X_13251_ _18872_/Q _13242_/A _12543_/X _13243_/A vssd1 vssd1 vccd1 vccd1 _18872_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_182_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12202_ _19251_/Q _12198_/X _12088_/X _12199_/X vssd1 vssd1 vccd1 vccd1 _19251_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_170_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13182_ _13202_/A vssd1 vssd1 vccd1 vccd1 _13182_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_135_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10394_ _14256_/A _10403_/A vssd1 vssd1 vccd1 vccd1 _14476_/A sky130_fd_sc_hd__or2_2
XFILLER_124_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12133_ _12171_/A vssd1 vssd1 vccd1 vccd1 _12150_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_135_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17990_ _18169_/CLK _17990_/D vssd1 vssd1 vccd1 vccd1 _17990_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16150__C1 _16147_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16941_ _19485_/Q hold156/X _16946_/S vssd1 vssd1 vccd1 vccd1 _16941_/X sky130_fd_sc_hd__mux2_1
XFILLER_78_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12064_ _15774_/A _12066_/A vssd1 vssd1 vccd1 vccd1 _12065_/S sky130_fd_sc_hd__or2_1
XFILLER_238_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11015_ _11015_/A vssd1 vssd1 vccd1 vccd1 _19656_/D sky130_fd_sc_hd__inv_2
X_19660_ _19846_/CLK _19660_/D repeater270/X vssd1 vssd1 vccd1 vccd1 _19660_/Q sky130_fd_sc_hd__dfrtp_1
X_16872_ _16871_/X _13548_/A _17536_/S vssd1 vssd1 vccd1 vccd1 _16872_/X sky130_fd_sc_hd__mux2_1
XANTENNA__17876__S0 _17908_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08995__A _19516_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14059__A2 _14003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18611_ _19041_/CLK _18611_/D repeater266/X vssd1 vssd1 vccd1 vccd1 _18611_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_93_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15823_ _15823_/A vssd1 vssd1 vccd1 vccd1 _16303_/A sky130_fd_sc_hd__clkbuf_2
X_19591_ _19591_/CLK _19591_/D hold346/A vssd1 vssd1 vccd1 vccd1 _19591_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__19542__RESET_B repeater221/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18542_ _18886_/CLK hold328/X repeater221/X vssd1 vssd1 vccd1 vccd1 _18543_/D sky130_fd_sc_hd__dfrtp_1
XFILLER_161_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15754_ _11173_/A _17926_/Q _11175_/A vssd1 vssd1 vccd1 vccd1 _15755_/B sky130_fd_sc_hd__o21a_1
XFILLER_234_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12966_ _12965_/X _18935_/Q _18934_/Q _18936_/Q vssd1 vssd1 vccd1 vccd1 _12966_/X
+ sky130_fd_sc_hd__and4b_1
X_14705_ _14705_/A vssd1 vssd1 vccd1 vccd1 _14705_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_206_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18473_ _18473_/CLK _18473_/D vssd1 vssd1 vccd1 vccd1 _18473_/Q sky130_fd_sc_hd__dfxtp_1
X_11917_ _19406_/Q _11914_/X _10885_/X _11915_/X vssd1 vssd1 vccd1 vccd1 _19406_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_233_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15685_ _18614_/Q vssd1 vssd1 vccd1 vccd1 _15688_/A sky130_fd_sc_hd__inv_2
XPHY_4470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12897_ _19273_/Q vssd1 vssd1 vccd1 vccd1 _12897_/Y sky130_fd_sc_hd__inv_2
XPHY_4481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17424_ _15768_/Y _11224_/Y _17546_/S vssd1 vssd1 vccd1 vccd1 _17424_/X sky130_fd_sc_hd__mux2_1
XANTENNA__17312__S _17566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14636_ _18262_/Q _14630_/X _09177_/X _14632_/X vssd1 vssd1 vccd1 vccd1 _18262_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_33_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11848_ _19435_/Q vssd1 vssd1 vccd1 vccd1 _11848_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17355_ _17354_/X _09449_/Y _17413_/S vssd1 vssd1 vccd1 vccd1 _17355_/X sky130_fd_sc_hd__mux2_1
XFILLER_220_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14567_ _14780_/A vssd1 vssd1 vccd1 vccd1 _14567_/X sky130_fd_sc_hd__buf_2
X_11779_ _11936_/A vssd1 vssd1 vccd1 vccd1 _12371_/A sky130_fd_sc_hd__clkbuf_2
X_16306_ _19698_/Q vssd1 vssd1 vccd1 vccd1 _16306_/Y sky130_fd_sc_hd__inv_2
X_13518_ _13500_/Y _13509_/X _13721_/A vssd1 vssd1 vccd1 vccd1 _13518_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_174_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17286_ _17285_/X _14074_/Y _17544_/S vssd1 vssd1 vccd1 vccd1 _17286_/X sky130_fd_sc_hd__mux2_1
XANTENNA__17800__S0 _17918_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14498_ _18341_/Q _14491_/X _12726_/X _14493_/X vssd1 vssd1 vccd1 vccd1 _18341_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18495__RESET_B repeater203/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19025_ _19157_/CLK _19025_/D repeater266/X vssd1 vssd1 vccd1 vccd1 _19025_/Q sky130_fd_sc_hd__dfrtp_4
X_16237_ _17386_/X _16598_/A vssd1 vssd1 vccd1 vccd1 _16237_/Y sky130_fd_sc_hd__nand2_2
X_13449_ _13428_/B _13344_/B _13447_/Y _13445_/X vssd1 vssd1 vccd1 vccd1 _18857_/D
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__16452__A _19772_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16168_ _19649_/Q _15799_/Y _11023_/Y _18227_/Q vssd1 vssd1 vccd1 vccd1 _16168_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_142_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15119_ _17978_/Q _15111_/A _14935_/X _15112_/A vssd1 vssd1 vccd1 vccd1 _17978_/D
+ sky130_fd_sc_hd__a22o_1
X_08990_ _11830_/A vssd1 vssd1 vccd1 vccd1 _12130_/A sky130_fd_sc_hd__buf_1
X_16099_ _17948_/Q vssd1 vssd1 vccd1 vccd1 _16099_/Y sky130_fd_sc_hd__inv_2
X_19927_ _19927_/CLK _19927_/D repeater235/X vssd1 vssd1 vccd1 vccd1 _19927_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_130_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17867__S0 _17908_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19858_ _19859_/CLK _19858_/D repeater261/X vssd1 vssd1 vccd1 vccd1 _19858_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_96_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09611_ _09471_/A _09471_/B _09609_/Y _09607_/X vssd1 vssd1 vccd1 vccd1 _20010_/D
+ sky130_fd_sc_hd__a211oi_2
X_18809_ _20115_/CLK _18809_/D repeater217/X vssd1 vssd1 vccd1 vccd1 _18809_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__19283__RESET_B repeater212/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19789_ _20089_/CLK _19789_/D repeater203/X vssd1 vssd1 vccd1 vccd1 _19789_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_83_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09542_ _19316_/Q vssd1 vssd1 vccd1 vccd1 _16647_/A sky130_fd_sc_hd__inv_2
X_09473_ _09473_/A _09473_/B vssd1 vssd1 vccd1 vccd1 _09605_/A sky130_fd_sc_hd__or2_2
XFILLER_36_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20117__RESET_B repeater217/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17222__S _17566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_212_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12233__A1 _19231_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15183__B1 _17936_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_147_HCLK_A clkbuf_4_1_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11744__B1 _16928_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold299_A HWDATA[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17858__S0 _17908_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19984__CLK _19984_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09809_ _09809_/A _09809_/B _09813_/C vssd1 vssd1 vccd1 vccd1 _19975_/D sky130_fd_sc_hd__nor3_1
XANTENNA__13249__B1 _12538_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12820_ _12815_/Y _18825_/Q _12816_/Y _18813_/Q _12819_/X vssd1 vssd1 vccd1 vccd1
+ _12833_/B sky130_fd_sc_hd__o221a_1
XANTENNA__14997__B1 _14996_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_216_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_234_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12751_ _12746_/Y _18831_/Q _19241_/Q _13541_/A _12750_/X vssd1 vssd1 vccd1 vccd1
+ _12758_/C sky130_fd_sc_hd__o221a_1
XPHY_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17132__S _17318_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11702_ _18622_/Q vssd1 vssd1 vccd1 vccd1 _11703_/A sky130_fd_sc_hd__inv_2
XFILLER_242_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15470_ _15470_/A vssd1 vssd1 vccd1 vccd1 _15475_/B sky130_fd_sc_hd__inv_2
XPHY_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12682_ _18978_/Q _12677_/X hold310/X _12678_/X vssd1 vssd1 vccd1 vccd1 _18978_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14421_ _18387_/Q _14410_/A _14403_/X _14411_/A vssd1 vssd1 vccd1 vccd1 _18387_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11633_ _19553_/Q _11632_/Y _11624_/B _11563_/X vssd1 vssd1 vccd1 vccd1 _19553_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16971__S _17524_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17140_ _17139_/X _19140_/Q _17548_/S vssd1 vssd1 vccd1 vccd1 _17140_/X sky130_fd_sc_hd__mux2_1
XPHY_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19364__CLK _19984_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14352_ _14352_/A vssd1 vssd1 vccd1 vccd1 _14353_/A sky130_fd_sc_hd__inv_2
XPHY_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11564_ _19577_/Q _11569_/B _11453_/Y _11562_/A _11563_/X vssd1 vssd1 vccd1 vccd1
+ _19577_/D sky130_fd_sc_hd__o221a_1
XPHY_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11983__B1 _11918_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13303_ _18862_/Q vssd1 vssd1 vccd1 vccd1 _13433_/A sky130_fd_sc_hd__inv_2
XFILLER_6_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10515_ _10734_/A _19536_/Q _10525_/D _19535_/Q vssd1 vssd1 vccd1 vccd1 _10516_/B
+ sky130_fd_sc_hd__or4b_4
X_17071_ _16665_/Y _18984_/Q _17493_/S vssd1 vssd1 vccd1 vccd1 _17071_/X sky130_fd_sc_hd__mux2_1
XANTENNA__15174__B1 hold236/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11495_ _19607_/Q _11494_/Y _11490_/X _11488_/B vssd1 vssd1 vccd1 vccd1 _19607_/D
+ sky130_fd_sc_hd__o211a_1
X_14283_ _18460_/Q _14274_/A _13678_/X _14275_/A vssd1 vssd1 vccd1 vccd1 _18460_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_155_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16022_ _18044_/Q vssd1 vssd1 vccd1 vccd1 _16022_/Y sky130_fd_sc_hd__inv_2
X_13234_ _18884_/Q _13231_/X _18545_/Q _17584_/S vssd1 vssd1 vccd1 vccd1 _18884_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_171_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10446_ _10446_/A vssd1 vssd1 vccd1 vccd1 _10446_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__10538__A1 _19814_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10377_ _10372_/B _10376_/Y _10368_/X _10354_/A _10322_/A vssd1 vssd1 vccd1 vccd1
+ _10378_/A sky130_fd_sc_hd__o32a_1
X_13165_ _13089_/A _13165_/A2 _13090_/Y _13199_/B vssd1 vssd1 vccd1 vccd1 _18917_/D
+ sky130_fd_sc_hd__a211oi_4
XANTENNA__19794__RESET_B repeater219/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_69_HCLK_A clkbuf_opt_3_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16674__B1 _16996_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12116_ _19305_/Q _12114_/X _12035_/X _12115_/X vssd1 vssd1 vccd1 vccd1 _19305_/D
+ sky130_fd_sc_hd__a22o_1
X_17973_ _20124_/CLK _17973_/D vssd1 vssd1 vccd1 vccd1 _17973_/Q sky130_fd_sc_hd__dfxtp_1
X_13096_ _13092_/Y _18918_/Q _19167_/Q _13069_/B _13095_/X vssd1 vssd1 vccd1 vccd1
+ _13109_/A sky130_fd_sc_hd__o221a_1
XFILLER_111_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19712_ _19794_/CLK _19712_/D repeater219/X vssd1 vssd1 vccd1 vccd1 _19712_/Q sky130_fd_sc_hd__dfstp_1
X_16924_ _16923_/X _09489_/A _17414_/S vssd1 vssd1 vccd1 vccd1 _16924_/X sky130_fd_sc_hd__mux2_1
XANTENNA__17307__S _17545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12047_ _19335_/Q _12043_/X _11918_/X _12044_/X vssd1 vssd1 vccd1 vccd1 _19335_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17849__S0 _18760_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12160__B1 _12026_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_238_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19643_ _19647_/CLK _19643_/D repeater261/X vssd1 vssd1 vccd1 vccd1 _19643_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_37_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16855_ _16854_/X _09690_/Y _17523_/S vssd1 vssd1 vccd1 vccd1 _16855_/X sky130_fd_sc_hd__mux2_1
XANTENNA__16977__A1 _18980_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15806_ _18266_/Q vssd1 vssd1 vccd1 vccd1 _15806_/Y sky130_fd_sc_hd__inv_2
X_19574_ _19595_/CLK _19574_/D repeater282/X vssd1 vssd1 vccd1 vccd1 _19574_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__14988__B1 _14780_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16786_ _16785_/X _15569_/Y _17513_/S vssd1 vssd1 vccd1 vccd1 _16786_/X sky130_fd_sc_hd__mux2_1
X_13998_ _18676_/Q vssd1 vssd1 vccd1 vccd1 _14007_/A sky130_fd_sc_hd__inv_2
XFILLER_241_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_114_HCLK clkbuf_opt_0_HCLK/A vssd1 vssd1 vccd1 vccd1 _19119_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_234_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18525_ _18886_/CLK _18525_/D repeater220/X vssd1 vssd1 vccd1 vccd1 _18527_/D sky130_fd_sc_hd__dfstp_1
XFILLER_80_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15737_ _18488_/D _15737_/B vssd1 vssd1 vccd1 vccd1 _18509_/D sky130_fd_sc_hd__nor2_1
XFILLER_65_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12463__A1 _19110_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12949_ _19283_/Q _12964_/A _19279_/Q _12878_/A vssd1 vssd1 vccd1 vccd1 _12949_/Y
+ sky130_fd_sc_hd__a22oi_2
XANTENNA__13660__B1 _12028_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_221_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18456_ _18465_/CLK _18456_/D vssd1 vssd1 vccd1 vccd1 _18456_/Q sky130_fd_sc_hd__dfxtp_1
X_15668_ _15668_/A _15668_/B vssd1 vssd1 vccd1 vccd1 _15669_/A sky130_fd_sc_hd__or2_1
XFILLER_178_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18676__RESET_B repeater252/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17407_ _17486_/A0 _16121_/Y _17517_/S vssd1 vssd1 vccd1 vccd1 _17407_/X sky130_fd_sc_hd__mux2_1
X_14619_ _18273_/Q _14616_/X _09168_/X _14618_/X vssd1 vssd1 vccd1 vccd1 _18273_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16881__S _17414_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18387_ _19515_/CLK _18387_/D vssd1 vssd1 vccd1 vccd1 _18387_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15599_ _15602_/B _15598_/Y _15590_/X vssd1 vssd1 vccd1 vccd1 _15599_/X sky130_fd_sc_hd__o21a_1
XFILLER_159_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17338_ _17337_/X _16368_/Y _17548_/S vssd1 vssd1 vccd1 vccd1 _17338_/X sky130_fd_sc_hd__mux2_1
XFILLER_202_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11974__B1 _11911_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17269_ _17268_/X _13070_/A _17542_/S vssd1 vssd1 vccd1 vccd1 _17269_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19008_ _19595_/CLK _19008_/D hold346/A vssd1 vssd1 vccd1 vccd1 _19008_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_134_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08973_ _20070_/Q vssd1 vssd1 vccd1 vccd1 _08978_/A sky130_fd_sc_hd__inv_2
XFILLER_29_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17217__S _17487_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17090__A0 _17486_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_216_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_2_0_HCLK clkbuf_4_3_0_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_2_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_09525_ _19300_/Q vssd1 vssd1 vccd1 vccd1 _09525_/Y sky130_fd_sc_hd__inv_2
XFILLER_231_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09456_ _10043_/A _19387_/Q _10039_/A _19383_/Q _09455_/X vssd1 vssd1 vccd1 vccd1
+ _09463_/C sky130_fd_sc_hd__o221a_1
XPHY_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_196_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09387_ _10009_/A _19394_/Q _10082_/A _19370_/Q vssd1 vssd1 vccd1 vccd1 _09387_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__16791__S _17546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09083__B1 _09082_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09622__A2 _10079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11965__B1 _09058_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10300_ _18595_/Q _15601_/A vssd1 vssd1 vccd1 vccd1 _15605_/A sky130_fd_sc_hd__or2_2
XANTENNA__17979__CLK _20123_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11280_ _18997_/Q vssd1 vssd1 vccd1 vccd1 _11280_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10231_ _19659_/Q vssd1 vssd1 vccd1 vccd1 _10959_/A sky130_fd_sc_hd__inv_2
XFILLER_193_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10162_ _19890_/Q _10155_/A _09101_/X _10156_/A vssd1 vssd1 vccd1 vccd1 _19890_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_160_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17127__S _17543_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10093_ _10086_/A _10086_/B _10091_/Y _10107_/C vssd1 vssd1 vccd1 vccd1 _19914_/D
+ sky130_fd_sc_hd__a211oi_2
X_14970_ _18070_/Q _14964_/X _14810_/X _14966_/X vssd1 vssd1 vccd1 vccd1 _18070_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_48_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12142__B1 _12080_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_137_HCLK clkbuf_4_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19992_/CLK sky130_fd_sc_hd__clkbuf_16
X_13921_ _13921_/A vssd1 vssd1 vccd1 vccd1 _13921_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16966__S _17474_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16640_ _17041_/X _16577_/X _16921_/X _16578_/X _16639_/X vssd1 vssd1 vccd1 vccd1
+ _16641_/C sky130_fd_sc_hd__o221a_1
X_13852_ _19202_/Q vssd1 vssd1 vccd1 vccd1 _13852_/Y sky130_fd_sc_hd__inv_2
XFILLER_223_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12803_ _19231_/Q vssd1 vssd1 vccd1 vccd1 _16211_/A sky130_fd_sc_hd__inv_2
XFILLER_28_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16571_ _15901_/A _15999_/X _17566_/S _16504_/A _16484_/X vssd1 vssd1 vccd1 vccd1
+ _16682_/A sky130_fd_sc_hd__a2111oi_2
X_13783_ _18729_/Q vssd1 vssd1 vccd1 vccd1 _13914_/A sky130_fd_sc_hd__inv_2
XFILLER_216_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10995_ _10995_/A vssd1 vssd1 vccd1 vccd1 _19662_/D sky130_fd_sc_hd__inv_2
X_18310_ _18431_/CLK _18310_/D vssd1 vssd1 vccd1 vccd1 _18310_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15522_ _18575_/Q vssd1 vssd1 vccd1 vccd1 _15526_/A sky130_fd_sc_hd__inv_2
XANTENNA__10456__B1 _10423_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12734_ _19258_/Q vssd1 vssd1 vccd1 vccd1 _12734_/Y sky130_fd_sc_hd__inv_2
X_19290_ _19290_/CLK _19290_/D repeater211/X vssd1 vssd1 vccd1 vccd1 _19290_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_231_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18241_ _20077_/CLK _18241_/D vssd1 vssd1 vccd1 vccd1 _18241_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15453_ _15453_/A vssd1 vssd1 vccd1 vccd1 _15453_/Y sky130_fd_sc_hd__inv_2
XPHY_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12665_ _18991_/Q _12661_/X hold284/X _12664_/X vssd1 vssd1 vccd1 vccd1 _18991_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_repeater169_A _16950_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14404_ _18395_/Q _14395_/A _14403_/X _14396_/A vssd1 vssd1 vccd1 vccd1 _18395_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11616_ _19559_/Q _11615_/Y _11588_/A _11573_/B vssd1 vssd1 vccd1 vccd1 _19559_/D
+ sky130_fd_sc_hd__o211a_1
X_18172_ _18198_/CLK _18172_/D vssd1 vssd1 vccd1 vccd1 _18172_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15384_ _15384_/A _17585_/X vssd1 vssd1 vccd1 vccd1 _18512_/D sky130_fd_sc_hd__and2_1
XPHY_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12596_ _14273_/A vssd1 vssd1 vccd1 vccd1 _12596_/X sky130_fd_sc_hd__buf_4
XPHY_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17123_ _17122_/X _13844_/Y _17545_/S vssd1 vssd1 vccd1 vccd1 _17123_/X sky130_fd_sc_hd__mux2_1
X_14335_ _14335_/A _14545_/B _14598_/C vssd1 vssd1 vccd1 vccd1 _14337_/A sky130_fd_sc_hd__or3_4
XPHY_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11547_ _11547_/A _11547_/B vssd1 vssd1 vccd1 vccd1 _11585_/A sky130_fd_sc_hd__or2_1
XFILLER_7_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16895__A0 _17473_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19975__RESET_B repeater244/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17054_ _17053_/X _09872_/A _17524_/S vssd1 vssd1 vccd1 vccd1 _17054_/X sky130_fd_sc_hd__mux2_1
XANTENNA_output98_A _16705_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14266_ _18468_/Q _14259_/A _12729_/X _14260_/A vssd1 vssd1 vccd1 vccd1 _18468_/D
+ sky130_fd_sc_hd__a22o_1
X_11478_ _11478_/A _11478_/B vssd1 vssd1 vccd1 vccd1 _11508_/A sky130_fd_sc_hd__or2_1
XFILLER_109_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19904__RESET_B repeater195/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_130_HCLK_A clkbuf_4_4_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16005_ _17558_/S _15992_/X _15996_/X _16001_/X _16004_/X vssd1 vssd1 vccd1 vccd1
+ _16005_/X sky130_fd_sc_hd__o2111a_1
X_13217_ _18530_/Q _13217_/B vssd1 vssd1 vccd1 vccd1 _13218_/B sky130_fd_sc_hd__or2_1
X_10429_ _10429_/A _11842_/B vssd1 vssd1 vccd1 vccd1 _16492_/A sky130_fd_sc_hd__or2_4
X_14197_ _19114_/Q _14023_/A _14196_/Y _18691_/Q vssd1 vssd1 vccd1 vccd1 _14197_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12035__A hold239/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12381__B1 _12380_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13148_ _19179_/Q vssd1 vssd1 vccd1 vccd1 _13148_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17037__S _17474_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13079_ _13079_/A _13079_/B vssd1 vssd1 vccd1 vccd1 _13179_/A sky130_fd_sc_hd__or2_1
X_17956_ _20076_/CLK _17956_/D vssd1 vssd1 vccd1 vccd1 _17956_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16907_ _16906_/X _19215_/Q _17545_/S vssd1 vssd1 vccd1 vccd1 _16907_/X sky130_fd_sc_hd__mux2_1
X_17887_ _16034_/Y _16035_/Y _16036_/Y _16037_/Y _17908_/S0 _18759_/Q vssd1 vssd1
+ vccd1 vccd1 _17887_/X sky130_fd_sc_hd__mux4_1
XFILLER_226_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16876__S _17534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19626_ _19825_/CLK _19626_/D repeater220/X vssd1 vssd1 vccd1 vccd1 _19626_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_26_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16838_ _17473_/A0 _16700_/Y _17547_/S vssd1 vssd1 vccd1 vccd1 _16838_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18857__RESET_B repeater231/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16769_ _15768_/Y _11205_/Y _17546_/S vssd1 vssd1 vccd1 vccd1 _16769_/X sky130_fd_sc_hd__mux2_1
X_19557_ _19582_/CLK _19557_/D hold348/A vssd1 vssd1 vccd1 vccd1 _19557_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_202_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09310_ _09308_/Y _15726_/A _09308_/Y _15726_/A vssd1 vssd1 vccd1 vccd1 _09333_/B
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__10447__B1 _10446_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_234_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18508_ _19780_/CLK _18508_/D repeater226/X vssd1 vssd1 vccd1 vccd1 _18508_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_202_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19488_ _19513_/CLK hold155/X repeater260/X vssd1 vssd1 vccd1 vccd1 _19488_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_179_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09241_ _09222_/Y _09224_/Y _19885_/Q _15713_/A _09240_/X vssd1 vssd1 vccd1 vccd1
+ _09241_/X sky130_fd_sc_hd__o221a_1
XFILLER_167_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18439_ _18441_/CLK _18439_/D vssd1 vssd1 vccd1 vccd1 _18439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17500__S _17565_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09172_ _14705_/A _09163_/X _09171_/X _09165_/X vssd1 vssd1 vccd1 vccd1 _20079_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09065__B1 _09064_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_18_HCLK clkbuf_4_3_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _18869_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__11947__B1 _09027_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16624__B _16673_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_10_0_HCLK clkbuf_3_5_0_HCLK/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_1_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__15138__B1 hold236/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18542__D hold328/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_52_HCLK_A clkbuf_opt_1_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11784__A _11800_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08956_ _18784_/Q vssd1 vssd1 vccd1 vccd1 _08956_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12124__B1 _11981_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09254__A hold322/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16786__S _17513_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18598__RESET_B repeater267/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16810__A0 _15768_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18777__CLK _19847_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09508_ _19299_/Q vssd1 vssd1 vccd1 vccd1 _09508_/Y sky130_fd_sc_hd__inv_2
XANTENNA__10438__B1 _09064_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10780_ _17629_/X _10773_/A _19744_/Q _10774_/A vssd1 vssd1 vccd1 vccd1 _19744_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09439_ _19932_/Q _09374_/Y _19916_/Q _09435_/Y _09438_/X vssd1 vssd1 vccd1 vccd1
+ _09440_/D sky130_fd_sc_hd__o221a_1
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15916__A2 _16683_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17410__S _17517_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09056__B1 hold276/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12450_ _12457_/A vssd1 vssd1 vccd1 vccd1 _12450_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_200_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11401_ _19573_/Q vssd1 vssd1 vccd1 vccd1 _11547_/B sky130_fd_sc_hd__inv_2
X_12381_ _19156_/Q _12374_/X _12380_/X _12378_/X vssd1 vssd1 vccd1 vccd1 _19156_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16326__C1 _16324_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14120_ _14120_/A vssd1 vssd1 vccd1 vccd1 _14120_/Y sky130_fd_sc_hd__clkinv_1
X_11332_ _18981_/Q vssd1 vssd1 vccd1 vccd1 _11332_/Y sky130_fd_sc_hd__inv_2
XFILLER_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14051_ _19071_/Q _14012_/A _19081_/Q _14022_/A vssd1 vssd1 vccd1 vccd1 _14051_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19402__CLK _19984_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11263_ _19605_/Q vssd1 vssd1 vccd1 vccd1 _11485_/A sky130_fd_sc_hd__inv_2
XFILLER_106_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12363__B1 _12299_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13002_ _13002_/A _13019_/A vssd1 vssd1 vccd1 vccd1 _13017_/A sky130_fd_sc_hd__or2_2
X_10214_ _19664_/Q vssd1 vssd1 vccd1 vccd1 _10964_/A sky130_fd_sc_hd__inv_2
XFILLER_122_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11194_ _17716_/X _11191_/X _19615_/Q _11192_/X vssd1 vssd1 vccd1 vccd1 _19615_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_106_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17810_ _18332_/Q _18212_/Q _18204_/Q _18196_/Q _17918_/S0 _18750_/Q vssd1 vssd1
+ vccd1 vccd1 _17810_/X sky130_fd_sc_hd__mux4_2
X_10145_ _19897_/Q _10136_/A _16980_/X _10138_/A vssd1 vssd1 vccd1 vccd1 _19897_/D
+ sky130_fd_sc_hd__a22o_1
X_18790_ _19647_/CLK _18790_/D repeater261/X vssd1 vssd1 vccd1 vccd1 _18790_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_95_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17741_ _15368_/X _19704_/Q _18508_/D vssd1 vssd1 vccd1 vccd1 _17741_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09164__A _09164_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10076_ _10036_/A _10036_/B _10079_/A _10074_/Y vssd1 vssd1 vccd1 vccd1 _19920_/D
+ sky130_fd_sc_hd__a211oi_2
X_14953_ _14953_/A vssd1 vssd1 vccd1 vccd1 _14954_/A sky130_fd_sc_hd__inv_2
XANTENNA_output136_A _19610_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13904_ _13927_/A vssd1 vssd1 vccd1 vccd1 _13970_/C sky130_fd_sc_hd__clkbuf_2
X_17672_ _15548_/X _19463_/Q _17683_/S vssd1 vssd1 vccd1 vccd1 _18580_/D sky130_fd_sc_hd__mux2_1
X_14884_ _14884_/A vssd1 vssd1 vccd1 vccd1 _14885_/A sky130_fd_sc_hd__inv_2
XFILLER_63_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16801__A0 _15963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16623_ _16723_/B vssd1 vssd1 vccd1 vccd1 _16673_/B sky130_fd_sc_hd__buf_2
X_19411_ _19984_/CLK _19411_/D repeater243/X vssd1 vssd1 vccd1 vccd1 _19411_/Q sky130_fd_sc_hd__dfrtp_4
X_13835_ _19212_/Q vssd1 vssd1 vccd1 vccd1 _13835_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15080__A2 _15072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16554_ _17138_/X _16508_/X _17132_/X _15908_/X _16553_/Y vssd1 vssd1 vccd1 vccd1
+ _16554_/X sky130_fd_sc_hd__o221a_1
X_19342_ _19964_/CLK _19342_/D hold372/X vssd1 vssd1 vccd1 vccd1 _19342_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__09295__B1 _09094_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13766_ _20039_/Q _19738_/Q _19733_/Q _13766_/D vssd1 vssd1 vccd1 vccd1 _13775_/S
+ sky130_fd_sc_hd__or4_4
X_10978_ _10978_/A vssd1 vssd1 vccd1 vccd1 _10978_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_15_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15505_ _15509_/B vssd1 vssd1 vccd1 vccd1 _15511_/B sky130_fd_sc_hd__inv_2
X_12717_ _14806_/A vssd1 vssd1 vccd1 vccd1 _12717_/X sky130_fd_sc_hd__clkbuf_2
X_19273_ _19283_/CLK _19273_/D repeater216/X vssd1 vssd1 vccd1 vccd1 _19273_/Q sky130_fd_sc_hd__dfrtp_1
X_16485_ _19448_/Q vssd1 vssd1 vccd1 vccd1 _16485_/Y sky130_fd_sc_hd__inv_2
XFILLER_231_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13697_ _14857_/A _14629_/B _13506_/Y _17760_/X _13696_/X vssd1 vssd1 vccd1 vccd1
+ _18765_/D sky130_fd_sc_hd__a41o_1
XANTENNA__17320__S _17524_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18224_ _20077_/CLK _18224_/D vssd1 vssd1 vccd1 vccd1 _18224_/Q sky130_fd_sc_hd__dfxtp_1
X_15436_ _15436_/A _18633_/Q vssd1 vssd1 vccd1 vccd1 _17569_/S sky130_fd_sc_hd__nor2_1
XFILLER_175_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12648_ _19000_/Q _12643_/X hold259/X _12644_/X vssd1 vssd1 vccd1 vccd1 _19000_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_129_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18155_ _18869_/CLK _18155_/D vssd1 vssd1 vccd1 vccd1 _18155_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15367_ _19783_/Q _10643_/B _10644_/B vssd1 vssd1 vccd1 vccd1 _15367_/X sky130_fd_sc_hd__a21bo_1
X_12579_ _19045_/Q _12576_/X _12404_/X _12577_/X vssd1 vssd1 vccd1 vccd1 _19045_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17106_ _16484_/X _08956_/Y _17566_/S vssd1 vssd1 vccd1 vccd1 _17106_/X sky130_fd_sc_hd__mux2_1
X_14318_ _14319_/A vssd1 vssd1 vccd1 vccd1 _14318_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__09339__A _14780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18086_ _20077_/CLK _18086_/D vssd1 vssd1 vccd1 vccd1 _18086_/Q sky130_fd_sc_hd__dfxtp_1
X_15298_ _15298_/A _15298_/B _15298_/C _15298_/D vssd1 vssd1 vccd1 vccd1 _15298_/X
+ sky130_fd_sc_hd__or4_1
Xhold306 input54/X vssd1 vssd1 vccd1 vccd1 hold306/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold317 hold317/A vssd1 vssd1 vccd1 vccd1 hold317/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold328 input76/X vssd1 vssd1 vccd1 vccd1 hold328/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold339 sda_i_S5 vssd1 vssd1 vccd1 vccd1 input78/A sky130_fd_sc_hd__dlygate4sd3_1
X_17037_ _17036_/X _15552_/A _17474_/S vssd1 vssd1 vccd1 vccd1 _17037_/X sky130_fd_sc_hd__mux2_1
X_14249_ _14366_/A _14758_/B _14758_/C vssd1 vssd1 vccd1 vccd1 _14251_/A sky130_fd_sc_hd__or3_4
XFILLER_113_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09790_ _09790_/A _09790_/B vssd1 vssd1 vccd1 vccd1 _09800_/A sky130_fd_sc_hd__or2_1
X_18988_ _19115_/CLK _18988_/D hold273/X vssd1 vssd1 vccd1 vccd1 _18988_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_39_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09074__A hold251/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17939_ _20036_/CLK _17939_/D vssd1 vssd1 vccd1 vccd1 _17939_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_227_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater156 _17523_/S vssd1 vssd1 vccd1 vccd1 _17517_/S sky130_fd_sc_hd__buf_8
Xrepeater167 _17522_/S vssd1 vssd1 vccd1 vccd1 _17543_/S sky130_fd_sc_hd__clkbuf_16
XFILLER_227_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater178 _17414_/S vssd1 vssd1 vccd1 vccd1 _17518_/S sky130_fd_sc_hd__buf_8
Xrepeater189 repeater190/X vssd1 vssd1 vccd1 vccd1 repeater189/X sky130_fd_sc_hd__buf_8
XANTENNA__18691__RESET_B hold359/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16619__B _16621_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19609_ _19609_/CLK _19609_/D hold359/X vssd1 vssd1 vccd1 vccd1 _19609_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10948__A _11771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18620__RESET_B hold351/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_195_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19897__RESET_B repeater195/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10840__A0 _10715_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17230__S _17566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09224_ _15713_/A vssd1 vssd1 vccd1 vccd1 _09224_/Y sky130_fd_sc_hd__inv_2
XANTENNA__09038__B1 _09037_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16571__A2 _15999_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19826__RESET_B repeater271/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11779__A _11936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09155_ _09144_/C _09154_/X _09151_/Y vssd1 vssd1 vccd1 vccd1 _20084_/D sky130_fd_sc_hd__a21oi_1
XFILLER_147_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12593__B1 _12356_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09086_ _10448_/A vssd1 vssd1 vccd1 vccd1 _09086_/X sky130_fd_sc_hd__buf_4
XFILLER_174_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12345__B1 _12344_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09988_ _09988_/A vssd1 vssd1 vccd1 vccd1 _09988_/Y sky130_fd_sc_hd__inv_2
X_08939_ _19859_/Q _18779_/Q _19859_/Q _18779_/Q vssd1 vssd1 vccd1 vccd1 _08943_/C
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__17036__A0 _17473_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17405__S _17512_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11950_ _19392_/Q _11948_/X _09030_/X _11949_/X vssd1 vssd1 vccd1 vccd1 _19392_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_245_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10901_ _19687_/Q _10894_/A _10866_/X _10895_/A vssd1 vssd1 vccd1 vccd1 _19687_/D
+ sky130_fd_sc_hd__a22o_1
X_11881_ _19430_/Q _11875_/X hold288/X _11878_/X vssd1 vssd1 vccd1 vccd1 _19430_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_245_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13620_ _13620_/A _13620_/B vssd1 vssd1 vccd1 vccd1 _13620_/Y sky130_fd_sc_hd__nand2_1
XFILLER_232_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10832_ _15349_/A _10831_/B _10829_/Y _10702_/Y _10840_/S vssd1 vssd1 vccd1 vccd1
+ _10833_/A sky130_fd_sc_hd__o32a_1
XFILLER_32_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09277__B1 _09101_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_213_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13551_ _13551_/A _13551_/B vssd1 vssd1 vccd1 vccd1 _13569_/A sky130_fd_sc_hd__or2_1
XFILLER_25_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10763_ _19753_/Q _10762_/X _10758_/B vssd1 vssd1 vccd1 vccd1 _19753_/D sky130_fd_sc_hd__o21a_1
XFILLER_241_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17140__S _17548_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12502_ _19085_/Q _12498_/X _12394_/X _12499_/X vssd1 vssd1 vccd1 vccd1 _19085_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_157_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16270_ _19637_/Q _16024_/Y _19638_/Q _16095_/Y vssd1 vssd1 vccd1 vccd1 _16270_/X
+ sky130_fd_sc_hd__a22o_1
X_13482_ _18841_/Q _13485_/A _13479_/A _13421_/X vssd1 vssd1 vccd1 vccd1 _18841_/D
+ sky130_fd_sc_hd__o211a_1
X_10694_ _17749_/X vssd1 vssd1 vccd1 vccd1 _10694_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16562__A2 _16505_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15221_ _15388_/A _15217_/Y _15218_/Y _15204_/X _15220_/Y vssd1 vssd1 vccd1 vccd1
+ _18638_/D sky130_fd_sc_hd__o221ai_1
XFILLER_185_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11689__A _15823_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12433_ _19128_/Q _12427_/X _12236_/X _12428_/X vssd1 vssd1 vccd1 vccd1 _19128_/D
+ sky130_fd_sc_hd__a22o_1
X_15152_ _17957_/Q _15146_/X _14707_/A _15148_/X vssd1 vssd1 vccd1 vccd1 _17957_/D
+ sky130_fd_sc_hd__a22o_1
X_12364_ _19163_/Q _12361_/X _12302_/X _12362_/X vssd1 vssd1 vccd1 vccd1 _19163_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_153_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14103_ _14030_/A _14030_/B _14101_/Y _14135_/B vssd1 vssd1 vccd1 vccd1 _18700_/D
+ sky130_fd_sc_hd__a211oi_2
X_11315_ _11303_/X _11315_/B _11315_/C _11315_/D vssd1 vssd1 vccd1 vccd1 _11362_/A
+ sky130_fd_sc_hd__and4b_1
X_15083_ _15084_/A vssd1 vssd1 vccd1 vccd1 _15083_/X sky130_fd_sc_hd__clkbuf_2
X_19960_ _19964_/CLK _19960_/D hold372/X vssd1 vssd1 vccd1 vccd1 _19960_/Q sky130_fd_sc_hd__dfrtp_1
X_12295_ _19201_/Q _12290_/X _12225_/X _12291_/X vssd1 vssd1 vccd1 vccd1 _19201_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08998__A _13280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12336__B1 _12095_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14034_ _18703_/Q vssd1 vssd1 vccd1 vccd1 _14034_/Y sky130_fd_sc_hd__inv_2
X_18911_ _19222_/CLK _18911_/D repeater188/X vssd1 vssd1 vccd1 vccd1 _18911_/Q sky130_fd_sc_hd__dfrtp_1
X_11246_ _19588_/Q _11244_/Y _19582_/Q _16208_/A vssd1 vssd1 vccd1 vccd1 _11246_/X
+ sky130_fd_sc_hd__o22a_1
X_19891_ _20055_/CLK _19891_/D repeater207/X vssd1 vssd1 vccd1 vccd1 _19891_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__20054__RESET_B repeater205/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18842_ _20107_/CLK _18842_/D repeater233/X vssd1 vssd1 vccd1 vccd1 _18842_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__10898__B1 _10885_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17814__A2 _17812_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11177_ _11191_/A vssd1 vssd1 vccd1 vccd1 _11192_/A sky130_fd_sc_hd__inv_2
XANTENNA__12313__A _12313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10128_ _18587_/Q _18586_/Q _15566_/A vssd1 vssd1 vccd1 vccd1 _15447_/B sky130_fd_sc_hd__or3_4
X_15985_ _18517_/Q vssd1 vssd1 vccd1 vccd1 _15985_/Y sky130_fd_sc_hd__inv_2
X_18773_ _19855_/CLK _18773_/D repeater264/X vssd1 vssd1 vccd1 vccd1 _18773_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_94_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17315__S _17566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17724_ _19676_/Q _19689_/Q _18510_/Q vssd1 vssd1 vccd1 vccd1 _17724_/X sky130_fd_sc_hd__mux2_1
X_10059_ _10059_/A vssd1 vssd1 vccd1 vccd1 _10059_/Y sky130_fd_sc_hd__inv_2
X_14936_ _18091_/Q _14922_/A _14935_/X _14923_/A vssd1 vssd1 vccd1 vccd1 _18091_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_36_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17655_ _15615_/X _19034_/Q _17655_/S vssd1 vssd1 vccd1 vccd1 _18597_/D sky130_fd_sc_hd__mux2_1
X_14867_ _18131_/Q _14859_/A _14713_/X _14860_/A vssd1 vssd1 vccd1 vccd1 _18131_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_24_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16250__A1 _17379_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16606_ _17240_/X _16577_/X _16863_/X _16578_/X _16605_/X vssd1 vssd1 vccd1 vccd1
+ _16607_/C sky130_fd_sc_hd__o221a_1
X_13818_ _13911_/A _13938_/A vssd1 vssd1 vccd1 vccd1 _13819_/B sky130_fd_sc_hd__or2_2
X_17586_ _19680_/Q _19717_/Q _18481_/Q vssd1 vssd1 vccd1 vccd1 _17586_/X sky130_fd_sc_hd__mux2_1
X_14798_ _18170_/Q _14786_/A _14782_/X _14787_/A vssd1 vssd1 vccd1 vccd1 _18170_/D
+ sky130_fd_sc_hd__a22o_1
X_19325_ _19325_/CLK _19325_/D repeater213/X vssd1 vssd1 vccd1 vccd1 _19325_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_32_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11075__B1 _19632_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16537_ _17196_/X _16687_/A _17187_/X _16509_/X vssd1 vssd1 vccd1 vccd1 _16537_/X
+ sky130_fd_sc_hd__o22a_1
X_13749_ _18746_/Q vssd1 vssd1 vccd1 vccd1 _13749_/Y sky130_fd_sc_hd__inv_2
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19990__RESET_B repeater192/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17050__S _17459_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19256_ _19324_/CLK _19256_/D repeater237/X vssd1 vssd1 vccd1 vccd1 _19256_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_31_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16468_ _16468_/A _16469_/B vssd1 vssd1 vccd1 vccd1 _16468_/Y sky130_fd_sc_hd__nor2_1
XFILLER_31_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15419_ _15419_/A _17571_/X vssd1 vssd1 vccd1 vccd1 _18541_/D sky130_fd_sc_hd__and2_1
XFILLER_164_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18207_ _19849_/CLK _18207_/D vssd1 vssd1 vccd1 vccd1 _18207_/Q sky130_fd_sc_hd__dfxtp_1
X_19187_ _19293_/CLK _19187_/D repeater187/X vssd1 vssd1 vccd1 vccd1 _19187_/Q sky130_fd_sc_hd__dfrtp_1
X_16399_ _18025_/Q vssd1 vssd1 vccd1 vccd1 _16399_/Y sky130_fd_sc_hd__inv_2
XFILLER_145_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_3_6_0_HCLK clkbuf_3_7_0_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_6_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12575__B1 _12398_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09069__A _09084_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18138_ _18142_/CLK _18138_/D vssd1 vssd1 vccd1 vccd1 _18138_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18069_ _18142_/CLK _18069_/D vssd1 vssd1 vccd1 vccd1 _18069_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold136 input15/X vssd1 vssd1 vccd1 vccd1 hold136/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold147 hold147/A vssd1 vssd1 vccd1 vccd1 hold147/X sky130_fd_sc_hd__dlygate4sd3_1
X_20100_ _20107_/CLK _20100_/D repeater234/X vssd1 vssd1 vccd1 vccd1 _20100_/Q sky130_fd_sc_hd__dfrtp_1
Xhold158 hold158/A vssd1 vssd1 vccd1 vccd1 hold158/X sky130_fd_sc_hd__dlygate4sd3_1
X_09911_ _09899_/X _09911_/B _09911_/C _09911_/D vssd1 vssd1 vccd1 vccd1 _09948_/B
+ sky130_fd_sc_hd__and4b_1
XFILLER_171_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold169 HADDR[10] vssd1 vssd1 vccd1 vccd1 input2/A sky130_fd_sc_hd__dlygate4sd3_1
X_20031_ _20115_/CLK _20031_/D repeater240/X vssd1 vssd1 vccd1 vccd1 _20031_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__10889__B1 _10866_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09842_ _19944_/Q vssd1 vssd1 vccd1 vccd1 _09853_/A sky130_fd_sc_hd__inv_2
XFILLER_59_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12223__A hold268/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18872__RESET_B repeater208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09773_ _19993_/Q _09772_/Y _09763_/X _09750_/B vssd1 vssd1 vccd1 vccd1 _19993_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__17225__S _17545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11302__A1 _11487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_227_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18815__CLK _20115_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_195_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19660__RESET_B repeater270/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09207_ _20068_/Q _09205_/Y _09205_/B _09206_/Y vssd1 vssd1 vccd1 vccd1 _20068_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_182_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12566__B1 _12382_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09138_ _09138_/A vssd1 vssd1 vccd1 vccd1 _15322_/B sky130_fd_sc_hd__buf_1
XFILLER_147_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09069_ _09084_/A vssd1 vssd1 vccd1 vccd1 _09069_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_163_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11100_ _19851_/Q vssd1 vssd1 vccd1 vccd1 _15094_/A sky130_fd_sc_hd__buf_1
XFILLER_135_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12080_ hold286/X vssd1 vssd1 vccd1 vccd1 _12080_/X sky130_fd_sc_hd__buf_2
XFILLER_116_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11031_ _19651_/Q _11022_/X _19651_/Q _11022_/X vssd1 vssd1 vccd1 vccd1 _11031_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_150_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17009__A0 _15768_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18542__RESET_B repeater221/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17135__S _17414_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16480__B2 _16688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15770_ _16669_/A vssd1 vssd1 vccd1 vccd1 _16721_/B sky130_fd_sc_hd__buf_4
X_12982_ _12967_/B _12883_/B _12978_/Y _13027_/C vssd1 vssd1 vccd1 vccd1 _18941_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_91_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14721_ _18216_/Q _14717_/X _14604_/X _14719_/X vssd1 vssd1 vccd1 vccd1 _18216_/D
+ sky130_fd_sc_hd__a22o_1
X_11933_ _11933_/A _12372_/A vssd1 vssd1 vccd1 vccd1 _11934_/S sky130_fd_sc_hd__or2_1
XFILLER_217_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16974__S _17536_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_232_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17440_ _17439_/X _15583_/Y _17513_/S vssd1 vssd1 vccd1 vccd1 _17440_/X sky130_fd_sc_hd__mux2_1
XFILLER_73_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14652_ _18251_/Q _14644_/A _09185_/X _14645_/A vssd1 vssd1 vccd1 vccd1 _18251_/D
+ sky130_fd_sc_hd__a22o_1
X_11864_ _19435_/Q _15233_/A _11856_/Y _10954_/B _11862_/A vssd1 vssd1 vccd1 vccd1
+ _11869_/B sky130_fd_sc_hd__a41o_1
XFILLER_232_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19748__RESET_B repeater205/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13603_ _13534_/A _13534_/B _13588_/X _13601_/Y vssd1 vssd1 vccd1 vccd1 _18810_/D
+ sky130_fd_sc_hd__a211oi_2
XPHY_3951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10815_ _17619_/X _10808_/X _19728_/Q _10810_/A vssd1 vssd1 vccd1 vccd1 _19728_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_14_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17371_ _16296_/Y _08937_/Y _17566_/S vssd1 vssd1 vccd1 vccd1 _17371_/X sky130_fd_sc_hd__mux2_1
XPHY_3962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14583_ _18292_/Q _14573_/A _14582_/X _14574_/A vssd1 vssd1 vccd1 vccd1 _18292_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_220_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11795_ _19465_/Q _11793_/X _09030_/X _11794_/X vssd1 vssd1 vccd1 vccd1 _19465_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19110_ _19115_/CLK _19110_/D hold353/X vssd1 vssd1 vccd1 vccd1 _19110_/Q sky130_fd_sc_hd__dfrtp_2
X_16322_ _17356_/X _16069_/X _17353_/X _16070_/X _16321_/X vssd1 vssd1 vccd1 vccd1
+ _16322_/X sky130_fd_sc_hd__o221a_1
X_13534_ _13534_/A _13534_/B vssd1 vssd1 vccd1 vccd1 _13601_/A sky130_fd_sc_hd__or2_1
X_10746_ _19761_/Q _10741_/X _10451_/X _10743_/X vssd1 vssd1 vccd1 vccd1 _19761_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19740__CLK _20051_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19041_ _19041_/CLK _19041_/D repeater266/X vssd1 vssd1 vccd1 vccd1 _19041_/Q sky130_fd_sc_hd__dfrtp_1
X_16253_ _18023_/Q vssd1 vssd1 vccd1 vccd1 _16253_/Y sky130_fd_sc_hd__inv_2
X_13465_ _13465_/A _13479_/A vssd1 vssd1 vccd1 vccd1 _13466_/B sky130_fd_sc_hd__or2_2
XFILLER_185_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_repeater151_A _17459_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10677_ _10677_/A vssd1 vssd1 vccd1 vccd1 _10677_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_repeater249_A hold370/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15204_ _15213_/A _18481_/Q vssd1 vssd1 vccd1 vccd1 _15204_/X sky130_fd_sc_hd__or2_2
X_12416_ _19141_/Q _12412_/X _12344_/X _12414_/X vssd1 vssd1 vccd1 vccd1 _19141_/D
+ sky130_fd_sc_hd__a22o_1
X_16184_ _18222_/Q vssd1 vssd1 vccd1 vccd1 _16184_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13396_ _13394_/Y _18843_/Q _20094_/Q _13322_/A _13395_/X vssd1 vssd1 vccd1 vccd1
+ _13402_/C sky130_fd_sc_hd__o221a_1
XFILLER_182_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15135_ _15135_/A vssd1 vssd1 vccd1 vccd1 _15136_/A sky130_fd_sc_hd__inv_2
XFILLER_142_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12347_ _19172_/Q _12341_/X hold281/X _12342_/X vssd1 vssd1 vccd1 vccd1 _19172_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19890__CLK _20070_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output80_A _16516_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15066_ _18013_/Q _15059_/X _14812_/A _15061_/X vssd1 vssd1 vccd1 vccd1 _18013_/D
+ sky130_fd_sc_hd__a22o_1
X_19943_ _19984_/CLK _19943_/D repeater244/X vssd1 vssd1 vccd1 vccd1 _19943_/Q sky130_fd_sc_hd__dfrtp_1
X_12278_ _19214_/Q _12276_/X _12095_/X _12277_/X vssd1 vssd1 vccd1 vccd1 _19214_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_4_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14017_ _14017_/A _14126_/A vssd1 vssd1 vccd1 vccd1 _14018_/B sky130_fd_sc_hd__or2_2
X_11229_ _19581_/Q _11224_/Y _19591_/Q _11225_/Y _11228_/X vssd1 vssd1 vccd1 vccd1
+ _11248_/A sky130_fd_sc_hd__o221a_1
X_19874_ _20064_/CLK _19874_/D repeater198/X vssd1 vssd1 vccd1 vccd1 _19874_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_122_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18825_ _19255_/CLK _18825_/D repeater217/X vssd1 vssd1 vccd1 vccd1 _18825_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_56_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17894__S1 _19634_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17045__S _17318_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18756_ _18869_/CLK _18756_/D repeater195/X vssd1 vssd1 vccd1 vccd1 _18756_/Q sky130_fd_sc_hd__dfrtp_4
X_15968_ _19686_/Q vssd1 vssd1 vccd1 vccd1 _15968_/Y sky130_fd_sc_hd__inv_2
X_17707_ _15433_/X _19770_/Q _18546_/D vssd1 vssd1 vccd1 vccd1 _17707_/X sky130_fd_sc_hd__mux2_1
XFILLER_224_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14919_ _15121_/A _15109_/B _14951_/C vssd1 vssd1 vccd1 vccd1 _14922_/A sky130_fd_sc_hd__or3_4
X_18687_ _18701_/CLK _18687_/D hold359/X vssd1 vssd1 vccd1 vccd1 _18687_/Q sky130_fd_sc_hd__dfrtp_4
X_15899_ _15899_/A vssd1 vssd1 vccd1 vccd1 _15900_/A sky130_fd_sc_hd__buf_1
XANTENNA__16884__S _17524_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16223__B2 _16055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17638_ _15689_/X _19051_/Q _17655_/S vssd1 vssd1 vccd1 vccd1 _18614_/D sky130_fd_sc_hd__mux2_1
XFILLER_64_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15801__B _16096_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17569_ _15438_/X _19822_/Q _17569_/S vssd1 vssd1 vccd1 vccd1 _17569_/X sky130_fd_sc_hd__mux2_1
XFILLER_210_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19418__RESET_B repeater271/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19308_ _20120_/CLK _19308_/D repeater238/X vssd1 vssd1 vccd1 vccd1 _19308_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_210_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19239_ _19314_/CLK _19239_/D repeater239/X vssd1 vssd1 vccd1 vccd1 _19239_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_192_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18667__SET_B repeater222/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20014_ _20032_/CLK _20014_/D repeater240/X vssd1 vssd1 vccd1 vccd1 _20014_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_58_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09825_ _19961_/Q vssd1 vssd1 vccd1 vccd1 _09869_/A sky130_fd_sc_hd__inv_2
XFILLER_101_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17885__S1 _18759_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09756_ _20001_/Q _09755_/Y _09667_/C _09755_/A _09731_/X vssd1 vssd1 vccd1 vccd1
+ _20001_/D sky130_fd_sc_hd__o221a_1
XFILLER_246_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14473__B1 hold334/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_107_HCLK_A clkbuf_4_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16794__S _17544_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09687_ _09744_/A _19417_/Q _19988_/Q _09686_/Y vssd1 vssd1 vccd1 vccd1 _09687_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_242_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13028__A1 _13021_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_199_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_214_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19841__RESET_B repeater270/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_202_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19159__RESET_B repeater188/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10600_ _18508_/Q _15224_/A vssd1 vssd1 vccd1 vccd1 _10600_/Y sky130_fd_sc_hd__nor2_2
XPHY_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11580_ _11580_/A _11603_/A vssd1 vssd1 vccd1 vccd1 _11581_/B sky130_fd_sc_hd__or2_1
XPHY_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10531_ _11655_/A _10531_/B vssd1 vssd1 vccd1 vccd1 _10531_/X sky130_fd_sc_hd__or2_2
XPHY_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12539__B1 _12538_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13250_ _18873_/Q _13242_/A _12541_/X _13243_/A vssd1 vssd1 vccd1 vccd1 _18873_/D
+ sky130_fd_sc_hd__a22o_1
X_10462_ _10462_/A vssd1 vssd1 vccd1 vccd1 _10462_/Y sky130_fd_sc_hd__inv_2
XFILLER_155_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16542__B _16544_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12201_ _19252_/Q _12198_/X _12086_/X _12199_/X vssd1 vssd1 vccd1 vccd1 _19252_/D
+ sky130_fd_sc_hd__a22o_1
X_13181_ _18908_/Q _13179_/Y _13180_/X _13181_/C1 vssd1 vssd1 vccd1 vccd1 _18908_/D
+ sky130_fd_sc_hd__o211a_1
X_10393_ _19848_/Q vssd1 vssd1 vccd1 vccd1 _10403_/A sky130_fd_sc_hd__inv_2
XFILLER_108_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18794__RESET_B repeater261/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12132_ _15772_/A _12316_/B vssd1 vssd1 vccd1 vccd1 _12171_/A sky130_fd_sc_hd__or2_2
XFILLER_124_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16969__S _17522_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18723__RESET_B repeater253/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16940_ _19484_/Q hold165/X _16946_/S vssd1 vssd1 vccd1 vccd1 _16940_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09707__B2 _19423_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12063_ _11991_/X _19327_/Q _12063_/S vssd1 vssd1 vccd1 vccd1 _19327_/D sky130_fd_sc_hd__mux2_1
XFILLER_49_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11014_ _11010_/B _11013_/X _10978_/X _10989_/A _10956_/D vssd1 vssd1 vccd1 vccd1
+ _11015_/A sky130_fd_sc_hd__o32a_1
XFILLER_238_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16871_ _16870_/X _13410_/Y _17535_/S vssd1 vssd1 vccd1 vccd1 _16871_/X sky130_fd_sc_hd__mux2_1
XANTENNA__17876__S1 _18759_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18610_ _19566_/CLK _18610_/D repeater266/X vssd1 vssd1 vccd1 vccd1 _18610_/Q sky130_fd_sc_hd__dfrtp_1
X_15822_ _19701_/Q vssd1 vssd1 vccd1 vccd1 _15822_/Y sky130_fd_sc_hd__inv_2
X_19590_ _19591_/CLK _19590_/D hold346/X vssd1 vssd1 vccd1 vccd1 _19590_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_93_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18541_ _19825_/CLK _18541_/D repeater223/X vssd1 vssd1 vccd1 vccd1 _18541_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_206_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15753_ _15753_/A _15753_/B vssd1 vssd1 vccd1 vccd1 _18518_/D sky130_fd_sc_hd__and2_1
X_12965_ _12965_/A _12965_/B _12965_/C _12965_/D vssd1 vssd1 vccd1 vccd1 _12965_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_161_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11916_ _19407_/Q _11914_/X _10882_/X _11915_/X vssd1 vssd1 vccd1 vccd1 _19407_/D
+ sky130_fd_sc_hd__a22o_1
X_14704_ _18224_/Q _14698_/X _14703_/X _14701_/X vssd1 vssd1 vccd1 vccd1 _18224_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_233_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15684_ _15688_/B _15683_/Y _15673_/X vssd1 vssd1 vccd1 vccd1 _15684_/X sky130_fd_sc_hd__o21a_1
X_18472_ _18473_/CLK _18472_/D vssd1 vssd1 vccd1 vccd1 _18472_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19582__RESET_B hold348/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12896_ _19268_/Q _13004_/A _19289_/Q _12888_/B _12895_/X vssd1 vssd1 vccd1 vccd1
+ _12908_/A sky130_fd_sc_hd__o221a_1
XPHY_4460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16717__B _16718_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_29_HCLK_A clkbuf_4_9_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17423_ _17422_/X _13887_/Y _17545_/S vssd1 vssd1 vccd1 vccd1 _17423_/X sky130_fd_sc_hd__mux2_1
X_14635_ _18263_/Q _14630_/X _09174_/X _14632_/X vssd1 vssd1 vccd1 vccd1 _18263_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11847_ _11841_/X _19436_/Q _11847_/S vssd1 vssd1 vccd1 vccd1 _19436_/D sky130_fd_sc_hd__mux2_1
XFILLER_199_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14518__A _14519_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17354_ _15963_/X _09508_/Y _17534_/S vssd1 vssd1 vccd1 vccd1 _17354_/X sky130_fd_sc_hd__mux2_1
X_14566_ _18300_/Q _14559_/A _14513_/X _14560_/A vssd1 vssd1 vccd1 vccd1 _18300_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_20_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17705__A1 _19772_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11778_ _12659_/A vssd1 vssd1 vccd1 vccd1 _15772_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_186_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16305_ _19714_/Q vssd1 vssd1 vccd1 vccd1 _16305_/Y sky130_fd_sc_hd__inv_2
X_13517_ _18759_/Q _13516_/A _13704_/A _13516_/Y vssd1 vssd1 vccd1 vccd1 _13721_/A
+ sky130_fd_sc_hd__o22a_1
X_10729_ _19766_/Q _10721_/A _10425_/X _10722_/A vssd1 vssd1 vccd1 vccd1 _19766_/D
+ sky130_fd_sc_hd__a22o_1
X_17285_ _15768_/Y _14194_/Y _17546_/S vssd1 vssd1 vccd1 vccd1 _17285_/X sky130_fd_sc_hd__mux2_1
XANTENNA__17800__S1 _18750_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12038__A hold250/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14497_ _18342_/Q _14491_/X _12723_/X _14493_/X vssd1 vssd1 vccd1 vccd1 _18342_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_118_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19024_ _19970_/CLK _19024_/D repeater249/X vssd1 vssd1 vccd1 vccd1 _19024_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_118_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16236_ _16633_/A vssd1 vssd1 vccd1 vccd1 _16598_/A sky130_fd_sc_hd__inv_2
X_13448_ _18858_/Q _13447_/Y _13426_/X _13346_/B vssd1 vssd1 vccd1 vccd1 _18858_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_162_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_51_HCLK clkbuf_opt_1_HCLK/A vssd1 vssd1 vccd1 vccd1 _19795_/CLK sky130_fd_sc_hd__clkbuf_16
X_16167_ _18046_/Q vssd1 vssd1 vccd1 vccd1 _16167_/Y sky130_fd_sc_hd__inv_2
X_13379_ _13377_/Y _18846_/Q _20100_/Q _13469_/A _13378_/X vssd1 vssd1 vccd1 vccd1
+ _13386_/B sky130_fd_sc_hd__o221a_1
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12950__B1 _12948_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15118_ _17979_/Q _15111_/A _14933_/X _15112_/A vssd1 vssd1 vccd1 vccd1 _17979_/D
+ sky130_fd_sc_hd__a22o_1
X_16098_ _18093_/Q vssd1 vssd1 vccd1 vccd1 _16098_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16879__S _17534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18510__CLK _19780_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19636__CLK _19851_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19926_ _19927_/CLK _19926_/D repeater235/X vssd1 vssd1 vccd1 vccd1 _19926_/Q sky130_fd_sc_hd__dfrtp_1
X_15049_ _15049_/A vssd1 vssd1 vccd1 vccd1 _15049_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_123_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12702__B1 _12533_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19857_ _19859_/CLK _19857_/D repeater265/X vssd1 vssd1 vccd1 vccd1 _19857_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17867__S1 _18759_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09610_ _20011_/Q _09609_/Y _09585_/A _09473_/B vssd1 vssd1 vccd1 vccd1 _20011_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_95_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18808_ _20122_/CLK _18808_/D repeater217/X vssd1 vssd1 vccd1 vccd1 _18808_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_28_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_228_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19788_ _20089_/CLK _19788_/D repeater203/X vssd1 vssd1 vccd1 vccd1 _19788_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__14455__B1 _14441_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09082__A _10446_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09541_ _19304_/Q vssd1 vssd1 vccd1 vccd1 _09541_/Y sky130_fd_sc_hd__inv_2
X_18739_ _20051_/CLK _18739_/D repeater209/X vssd1 vssd1 vccd1 vccd1 _18739_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17503__S _17568_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09472_ _09472_/A _09609_/A vssd1 vssd1 vccd1 vccd1 _09473_/B sky130_fd_sc_hd__or2_2
XPHY_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18040__CLK _19851_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11787__A _11801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10691__A _12257_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11744__B2 _11738_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16789__S _17459_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18190__CLK _18198_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14143__C1 _14112_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold194_A HADDR[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14694__B1 _14693_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17858__S1 _18759_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09808_ _09635_/B _09810_/A _09635_/A vssd1 vssd1 vccd1 vccd1 _09809_/B sky130_fd_sc_hd__o21a_1
XFILLER_75_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10180__B1 _09108_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14446__B1 _14417_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_216_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09739_ _09787_/B _09739_/B vssd1 vssd1 vccd1 vccd1 _09740_/B sky130_fd_sc_hd__or2_2
XFILLER_28_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12130__B _12130_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17413__S _17413_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11027__A _15296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12750_ _19256_/Q _13556_/A _16668_/A _18828_/Q vssd1 vssd1 vccd1 vccd1 _12750_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_28_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11701_ _19520_/Q _11671_/X _11661_/Y vssd1 vssd1 vccd1 vccd1 _19520_/D sky130_fd_sc_hd__o21a_1
XFILLER_203_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12681_ _18979_/Q _12677_/X hold318/X _12678_/X vssd1 vssd1 vccd1 vccd1 _18979_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_230_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10866__A _13678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_242_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14420_ _18388_/Q _14410_/A _14419_/X _14411_/A vssd1 vssd1 vccd1 vccd1 _18388_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11632_ _11632_/A vssd1 vssd1 vccd1 vccd1 _11632_/Y sky130_fd_sc_hd__inv_2
XPHY_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19509__CLK _19510_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_74_HCLK clkbuf_opt_4_HCLK/A vssd1 vssd1 vccd1 vccd1 _18852_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14351_ _14745_/A vssd1 vssd1 vccd1 vccd1 _14351_/X sky130_fd_sc_hd__clkbuf_2
XPHY_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11563_ _11592_/A vssd1 vssd1 vccd1 vccd1 _11563_/X sky130_fd_sc_hd__clkbuf_2
XPHY_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13302_ _18863_/Q vssd1 vssd1 vccd1 vccd1 _13350_/A sky130_fd_sc_hd__inv_2
XANTENNA__17794__S0 _19647_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10514_ _19534_/Q _19533_/Q _10514_/C _10514_/D vssd1 vssd1 vccd1 vccd1 _10525_/D
+ sky130_fd_sc_hd__or4_4
XPHY_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17070_ _17069_/X _20028_/Q _17414_/S vssd1 vssd1 vccd1 vccd1 _17070_/X sky130_fd_sc_hd__mux2_2
XPHY_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14282_ _18461_/Q _14272_/X _13676_/X _14275_/X vssd1 vssd1 vccd1 vccd1 _18461_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_144_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11494_ _11494_/A vssd1 vssd1 vccd1 vccd1 _11494_/Y sky130_fd_sc_hd__inv_2
X_16021_ _18468_/Q vssd1 vssd1 vccd1 vccd1 _16021_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18904__RESET_B repeater212/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13233_ _18885_/Q _13231_/X _18884_/Q _17584_/S vssd1 vssd1 vccd1 vccd1 _18885_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__15169__A _15169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10445_ _19834_/Q _10441_/X _09079_/X _10442_/X vssd1 vssd1 vccd1 vccd1 _19834_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_108_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13164_ _13202_/A vssd1 vssd1 vccd1 vccd1 _13199_/B sky130_fd_sc_hd__clkbuf_4
X_10376_ _19856_/Q _10376_/B vssd1 vssd1 vccd1 vccd1 _10376_/Y sky130_fd_sc_hd__nor2_1
XFILLER_124_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12115_ _12122_/A vssd1 vssd1 vccd1 vccd1 _12115_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__13488__A1 _13483_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13095_ _16468_/A _18895_/Q _16585_/A _18904_/Q vssd1 vssd1 vccd1 vccd1 _13095_/X
+ sky130_fd_sc_hd__o22a_1
X_17972_ _18765_/CLK _17972_/D vssd1 vssd1 vccd1 vccd1 _17972_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14685__B1 _14600_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19711_ _19720_/CLK _19711_/D repeater201/X vssd1 vssd1 vccd1 vccd1 _19711_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_111_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16923_ _16922_/X _09420_/Y _17413_/S vssd1 vssd1 vccd1 vccd1 _16923_/X sky130_fd_sc_hd__mux2_1
X_12046_ _19336_/Q _12043_/X _11981_/X _12044_/X vssd1 vssd1 vccd1 vccd1 _19336_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_120_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17849__S1 _18761_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19642_ _19647_/CLK _19642_/D repeater261/X vssd1 vssd1 vccd1 vccd1 _19642_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_238_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16854_ _17473_/A0 _09883_/Y _17522_/S vssd1 vssd1 vccd1 vccd1 _16854_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12321__A _12335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10171__B1 _09082_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15805_ _17969_/Q vssd1 vssd1 vccd1 vccd1 _15805_/Y sky130_fd_sc_hd__inv_2
X_19573_ _19576_/CLK _19573_/D repeater282/X vssd1 vssd1 vccd1 vccd1 _19573_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_92_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13997_ _18677_/Q vssd1 vssd1 vccd1 vccd1 _14008_/A sky130_fd_sc_hd__inv_2
X_16785_ _17473_/A0 _16729_/Y _17512_/S vssd1 vssd1 vccd1 vccd1 _16785_/X sky130_fd_sc_hd__mux2_1
XFILLER_92_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17323__S _17518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18524_ _18886_/CLK _18524_/D repeater220/X vssd1 vssd1 vccd1 vccd1 _18526_/D sky130_fd_sc_hd__dfstp_2
XFILLER_52_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15736_ _10658_/A _17925_/Q _10660_/A vssd1 vssd1 vccd1 vccd1 _15737_/B sky130_fd_sc_hd__o21a_1
X_12948_ _19277_/Q vssd1 vssd1 vccd1 vccd1 _12948_/Y sky130_fd_sc_hd__inv_2
XFILLER_234_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20016__CLK _20091_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_153_HCLK_A clkbuf_4_1_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18455_ _18465_/CLK _18455_/D vssd1 vssd1 vccd1 vccd1 _18455_/Q sky130_fd_sc_hd__dfxtp_1
X_12879_ _12965_/B _12879_/B vssd1 vssd1 vccd1 vccd1 _12988_/A sky130_fd_sc_hd__or2_1
X_15667_ _18610_/Q vssd1 vssd1 vccd1 vccd1 _15667_/Y sky130_fd_sc_hd__inv_2
XPHY_4290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17406_ _17405_/X _15587_/Y _17513_/S vssd1 vssd1 vccd1 vccd1 _17406_/X sky130_fd_sc_hd__mux2_1
X_14618_ _14618_/A vssd1 vssd1 vccd1 vccd1 _14618_/X sky130_fd_sc_hd__clkbuf_2
X_18386_ _19515_/CLK _18386_/D vssd1 vssd1 vccd1 vccd1 _18386_/Q sky130_fd_sc_hd__dfxtp_1
X_15598_ _15598_/A _15598_/B vssd1 vssd1 vccd1 vccd1 _15598_/Y sky130_fd_sc_hd__nor2_1
XFILLER_60_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14549_ _18313_/Q _14546_/X _14531_/X _14548_/X vssd1 vssd1 vccd1 vccd1 _18313_/D
+ sky130_fd_sc_hd__a22o_1
X_17337_ _17336_/X _11328_/Y _17459_/S vssd1 vssd1 vccd1 vccd1 _17337_/X sky130_fd_sc_hd__mux2_1
XANTENNA__17785__S0 _17923_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15165__B2 _15160_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17268_ _17267_/X _12897_/Y _17541_/S vssd1 vssd1 vccd1 vccd1 _17268_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19007_ _19595_/CLK _19007_/D hold346/A vssd1 vssd1 vccd1 vccd1 _19007_/Q sky130_fd_sc_hd__dfrtp_4
X_16219_ _19697_/Q vssd1 vssd1 vccd1 vccd1 _16219_/Y sky130_fd_sc_hd__inv_2
X_17199_ _17198_/X _11380_/Y _17548_/S vssd1 vssd1 vccd1 vccd1 _17199_/X sky130_fd_sc_hd__mux2_1
XFILLER_155_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09077__A hold268/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_216_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08972_ _13496_/C vssd1 vssd1 vccd1 vccd1 _17605_/S sky130_fd_sc_hd__clkbuf_4
X_19909_ _20006_/CLK _19909_/D repeater191/X vssd1 vssd1 vccd1 vccd1 _19909_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_69_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10162__B1 _09101_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_232_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16638__A _16638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09524_ _20004_/Q _09521_/Y _09483_/A _19313_/Q _09523_/X vssd1 vssd1 vccd1 vccd1
+ _09528_/C sky130_fd_sc_hd__o221a_1
XANTENNA__17233__S _17545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_97_HCLK clkbuf_4_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19968_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_25_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09455_ _19921_/Q _09453_/Y _10037_/A _19381_/Q vssd1 vssd1 vccd1 vccd1 _09455_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09386_ _19916_/Q vssd1 vssd1 vccd1 vccd1 _10088_/A sky130_fd_sc_hd__inv_2
XFILLER_12_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_12_HCLK_A clkbuf_4_2_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_0_HCLK_A clkbuf_4_0_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17776__S0 _17923_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold207_A HADDR[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_3_HCLK clkbuf_4_0_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19851_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__12406__A hold318/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12914__B1 _12913_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10230_ _19832_/Q vssd1 vssd1 vccd1 vccd1 _10230_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17408__S _17518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15717__A _19876_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10161_ _19891_/Q _10154_/X _09098_/X _10156_/X vssd1 vssd1 vccd1 vccd1 _19891_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_160_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10092_ _19915_/Q _10091_/Y _10088_/B _10026_/X vssd1 vssd1 vccd1 vccd1 _19915_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_48_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_248_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13920_ _13829_/A _13829_/B _13919_/X _13917_/Y vssd1 vssd1 vccd1 vccd1 _18730_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20039__CLK _20051_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13851_ _19206_/Q vssd1 vssd1 vccd1 vccd1 _13851_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15092__B1 _09339_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12802_ _18814_/Q vssd1 vssd1 vccd1 vccd1 _13537_/A sky130_fd_sc_hd__inv_2
XANTENNA__17143__S _17548_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16570_ _19041_/Q vssd1 vssd1 vccd1 vccd1 _16570_/Y sky130_fd_sc_hd__inv_2
X_13782_ _13782_/A vssd1 vssd1 vccd1 vccd1 _13829_/A sky130_fd_sc_hd__inv_2
X_10994_ _10988_/B _10978_/A _10993_/Y _10989_/X _10962_/A vssd1 vssd1 vccd1 vccd1
+ _10995_/A sky130_fd_sc_hd__o32a_1
XFILLER_231_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20079__RESET_B repeater205/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15521_ _15526_/B _15520_/X _15512_/X vssd1 vssd1 vccd1 vccd1 _15521_/X sky130_fd_sc_hd__o21a_1
X_12733_ _19259_/Q vssd1 vssd1 vccd1 vccd1 _12733_/Y sky130_fd_sc_hd__inv_2
XFILLER_231_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20008__RESET_B repeater241/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15452_ _18558_/Q vssd1 vssd1 vccd1 vccd1 _15452_/Y sky130_fd_sc_hd__inv_2
X_18240_ _20079_/CLK _18240_/D vssd1 vssd1 vccd1 vccd1 _18240_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12664_ _12678_/A vssd1 vssd1 vccd1 vccd1 _12664_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_70_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16592__B1 _17237_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14403_ hold335/X vssd1 vssd1 vccd1 vccd1 _14403_/X sky130_fd_sc_hd__buf_2
XPHY_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11615_ _11615_/A vssd1 vssd1 vccd1 vccd1 _11615_/Y sky130_fd_sc_hd__inv_2
XPHY_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15383_ _18639_/Q _17586_/X _18637_/Q _15382_/X vssd1 vssd1 vccd1 vccd1 _15383_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18171_ _18460_/CLK _18171_/D vssd1 vssd1 vccd1 vccd1 _18171_/Q sky130_fd_sc_hd__dfxtp_1
X_12595_ _19033_/Q _12590_/X hold259/X _12591_/X vssd1 vssd1 vccd1 vccd1 _19033_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17767__S0 _17923_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14334_ _14334_/A _19641_/Q _15296_/B vssd1 vssd1 vccd1 vccd1 _14598_/C sky130_fd_sc_hd__or3_4
XPHY_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17122_ _17121_/X _14087_/Y _17544_/S vssd1 vssd1 vccd1 vccd1 _17122_/X sky130_fd_sc_hd__mux2_1
X_11546_ _11570_/A vssd1 vssd1 vccd1 vccd1 _11639_/B sky130_fd_sc_hd__clkbuf_2
XPHY_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17053_ _17052_/X _09673_/Y _17523_/S vssd1 vssd1 vccd1 vccd1 _17053_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14265_ _18469_/Q _14258_/X _12726_/X _14260_/X vssd1 vssd1 vccd1 vccd1 _18469_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_repeater231_A repeater232/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11477_ _11477_/A _11511_/A vssd1 vssd1 vccd1 vccd1 _11478_/B sky130_fd_sc_hd__or2_1
XFILLER_143_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12316__A _15769_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16004_ _17476_/X _16002_/X _17485_/X _16003_/X vssd1 vssd1 vccd1 vccd1 _16004_/X
+ sky130_fd_sc_hd__o22a_1
X_13216_ _18529_/Q _18528_/Q vssd1 vssd1 vccd1 vccd1 _13217_/B sky130_fd_sc_hd__or2_1
X_10428_ _19842_/Q _10417_/X _10427_/X _10419_/Y vssd1 vssd1 vccd1 vccd1 _19842_/D
+ sky130_fd_sc_hd__a22o_1
X_14196_ _19112_/Q vssd1 vssd1 vccd1 vccd1 _14196_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17844__A0 _17840_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17318__S _17318_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13147_ _19162_/Q _13064_/A _13145_/Y _18890_/Q _13146_/X vssd1 vssd1 vccd1 vccd1
+ _13159_/A sky130_fd_sc_hd__o221a_1
X_10359_ _10353_/B _10368_/A _10358_/Y _10354_/X _10327_/A vssd1 vssd1 vccd1 vccd1
+ _10360_/A sky130_fd_sc_hd__o32a_1
XFILLER_98_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19944__RESET_B repeater244/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17955_ _20076_/CLK _17955_/D vssd1 vssd1 vccd1 vccd1 _17955_/Q sky130_fd_sc_hd__dfxtp_1
X_13078_ _13078_/A _13184_/A vssd1 vssd1 vccd1 vccd1 _13079_/B sky130_fd_sc_hd__or2_2
X_16906_ _16644_/Y _19083_/Q _17490_/S vssd1 vssd1 vccd1 vccd1 _16906_/X sky130_fd_sc_hd__mux2_2
XFILLER_39_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12029_ _19345_/Q _12023_/X _12028_/X _12024_/X vssd1 vssd1 vccd1 vccd1 _19345_/D
+ sky130_fd_sc_hd__a22o_1
X_17886_ _16030_/Y _16031_/Y _16032_/Y _16033_/Y _17908_/S0 _18759_/Q vssd1 vssd1
+ vccd1 vccd1 _17886_/X sky130_fd_sc_hd__mux4_2
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19625_ _19920_/CLK _19625_/D repeater229/X vssd1 vssd1 vccd1 vccd1 _19625_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__10695__A1 _10446_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16837_ _16836_/X _13091_/Y _17488_/S vssd1 vssd1 vccd1 vccd1 _16837_/X sky130_fd_sc_hd__mux2_2
XANTENNA__17053__S _17523_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15362__A _15364_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19556_ _19582_/CLK _19556_/D hold346/A vssd1 vssd1 vccd1 vccd1 _19556_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_81_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16768_ _16767_/X _13535_/A _17386_/S vssd1 vssd1 vccd1 vccd1 _16768_/X sky130_fd_sc_hd__mux2_2
XFILLER_19_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14830__B1 _14782_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18507_ _19812_/CLK _18507_/D repeater222/X vssd1 vssd1 vccd1 vccd1 _18507_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_202_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15719_ _19879_/Q _10286_/A _15718_/Y _19872_/Q _10759_/C vssd1 vssd1 vccd1 vccd1
+ _17631_/S sky130_fd_sc_hd__a221oi_2
X_19487_ _19510_/CLK hold161/X repeater260/X vssd1 vssd1 vccd1 vccd1 _19487_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__16892__S _17543_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_221_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16699_ _19466_/Q vssd1 vssd1 vccd1 vccd1 _16699_/Y sky130_fd_sc_hd__inv_2
X_09240_ _19883_/Q _15711_/A _09232_/X _09236_/X _09239_/X vssd1 vssd1 vccd1 vccd1
+ _09240_/X sky130_fd_sc_hd__o2111a_1
XFILLER_178_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18438_ _18441_/CLK _18438_/D vssd1 vssd1 vccd1 vccd1 _18438_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18826__RESET_B repeater217/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09171_ _14703_/A vssd1 vssd1 vccd1 vccd1 _09171_/X sky130_fd_sc_hd__clkbuf_2
X_18369_ _18441_/CLK _18369_/D vssd1 vssd1 vccd1 vccd1 _18369_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19974__CLK _19984_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10080__C1 _10107_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17228__S _17517_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09535__A _19317_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08955_ _10321_/D _18775_/Q _10331_/A _18785_/Q _08954_/X vssd1 vssd1 vccd1 vccd1
+ _08969_/B sky130_fd_sc_hd__o221a_1
XFILLER_130_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11883__B1 _09027_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15074__B1 hold247/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16368__A _19132_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_hold157_A HADDR[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09507_ _09491_/A _19321_/Q _20018_/Q _16547_/A _09506_/X vssd1 vssd1 vccd1 vccd1
+ _09512_/C sky130_fd_sc_hd__o221a_1
XFILLER_25_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09270__A _09270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09438_ _19922_/Q _09436_/Y _10038_/A _19382_/Q vssd1 vssd1 vccd1 vccd1 _09438_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_13_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18567__RESET_B repeater271/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09369_ _20008_/Q vssd1 vssd1 vccd1 vccd1 _09469_/A sky130_fd_sc_hd__inv_1
XFILLER_178_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11399__C1 _11398_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11400_ _19548_/Q vssd1 vssd1 vccd1 vccd1 _11548_/B sky130_fd_sc_hd__inv_2
X_12380_ hold291/X vssd1 vssd1 vccd1 vccd1 _12380_/X sky130_fd_sc_hd__buf_2
XFILLER_193_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16877__A1 _09414_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11331_ _11319_/X _11331_/B _11331_/C _11331_/D vssd1 vssd1 vccd1 vccd1 _11362_/B
+ sky130_fd_sc_hd__and4b_1
XFILLER_193_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14888__B1 _14808_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14050_ _19067_/Q vssd1 vssd1 vccd1 vccd1 _14050_/Y sky130_fd_sc_hd__inv_2
XFILLER_180_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11262_ _19598_/Q vssd1 vssd1 vccd1 vccd1 _11478_/A sky130_fd_sc_hd__inv_2
XFILLER_4_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_104_HCLK clkbuf_4_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19290_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_134_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16550__B _16622_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13001_ _13021_/A _13021_/B _13001_/C vssd1 vssd1 vccd1 vccd1 _13019_/A sky130_fd_sc_hd__or3_1
X_10213_ _19837_/Q vssd1 vssd1 vccd1 vccd1 _10213_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17138__S _17513_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11975__A _14273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15447__A _15479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11193_ _17715_/X _11191_/X _19616_/Q _11192_/X vssd1 vssd1 vccd1 vccd1 _19616_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_239_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17921__S0 _17923_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10144_ _16981_/X _10136_/A _19898_/Q _10138_/A vssd1 vssd1 vccd1 vccd1 _19898_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_239_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16977__S _17493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19355__RESET_B hold370/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17740_ _15369_/X _19705_/Q _18508_/D vssd1 vssd1 vccd1 vccd1 _17740_/X sky130_fd_sc_hd__mux2_1
X_10075_ _19921_/Q _10074_/Y _10026_/A _10038_/B vssd1 vssd1 vccd1 vccd1 _19921_/D
+ sky130_fd_sc_hd__o211a_1
X_14952_ _14953_/A vssd1 vssd1 vccd1 vccd1 _14952_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_75_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13903_ _13903_/A vssd1 vssd1 vccd1 vccd1 _13927_/A sky130_fd_sc_hd__clkbuf_2
X_17671_ _15553_/X _19464_/Q _17683_/S vssd1 vssd1 vccd1 vccd1 _18581_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14883_ _14884_/A vssd1 vssd1 vccd1 vccd1 _14883_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_75_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output129_A _19732_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19847__CLK _19847_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19410_ _19984_/CLK _19410_/D repeater193/X vssd1 vssd1 vccd1 vccd1 _19410_/Q sky130_fd_sc_hd__dfrtp_4
X_16622_ _19459_/Q _16622_/B vssd1 vssd1 vccd1 vccd1 _16622_/Y sky130_fd_sc_hd__nand2_1
XFILLER_75_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13834_ _18735_/Q vssd1 vssd1 vccd1 vccd1 _13834_/Y sky130_fd_sc_hd__inv_2
XFILLER_235_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19341_ _19352_/CLK _19341_/D repeater245/X vssd1 vssd1 vccd1 vccd1 _19341_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16553_ _17140_/X _16594_/A _17131_/X _16595_/A vssd1 vssd1 vccd1 vccd1 _16553_/Y
+ sky130_fd_sc_hd__a22oi_4
X_13765_ _18745_/Q _13760_/X _18745_/Q _13760_/X vssd1 vssd1 vccd1 vccd1 _18745_/D
+ sky130_fd_sc_hd__o2bb2a_1
X_10977_ _10973_/A _10955_/Y _10976_/X _10954_/A _19666_/Q vssd1 vssd1 vccd1 vccd1
+ _19666_/D sky130_fd_sc_hd__a32o_1
XFILLER_203_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15504_ _18571_/Q vssd1 vssd1 vccd1 vccd1 _15504_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15910__A _15999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17601__S _17605_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12716_ _18957_/Q vssd1 vssd1 vccd1 vccd1 _14808_/A sky130_fd_sc_hd__clkbuf_2
X_19272_ _19282_/CLK _19272_/D repeater216/X vssd1 vssd1 vccd1 vccd1 _19272_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_231_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16565__B1 _17169_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16484_ _16484_/A vssd1 vssd1 vccd1 vccd1 _16484_/X sky130_fd_sc_hd__buf_2
X_13696_ _13700_/A _13523_/A _14642_/A vssd1 vssd1 vccd1 vccd1 _13696_/X sky130_fd_sc_hd__o21a_1
XFILLER_231_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18223_ _20077_/CLK _18223_/D vssd1 vssd1 vccd1 vccd1 _18223_/Q sky130_fd_sc_hd__dfxtp_1
X_15435_ _19626_/Q _11170_/X _19626_/Q _11170_/X vssd1 vssd1 vccd1 vccd1 _15435_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_30_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12647_ _19001_/Q _12643_/X hold267/X _12644_/X vssd1 vssd1 vccd1 vccd1 _19001_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_129_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14040__A1 _14039_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15366_ _19782_/Q _19781_/Q _10643_/B vssd1 vssd1 vccd1 vccd1 _15366_/X sky130_fd_sc_hd__a21bo_1
X_18154_ _19900_/CLK _18154_/D vssd1 vssd1 vccd1 vccd1 _18154_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12051__B1 _11926_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12578_ _19046_/Q _12576_/X _12401_/X _12577_/X vssd1 vssd1 vccd1 vccd1 _19046_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_8_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17105_ _17104_/X _19201_/Q _17545_/S vssd1 vssd1 vccd1 vccd1 _17105_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14317_ _14335_/A _14317_/B _15070_/C vssd1 vssd1 vccd1 vccd1 _14319_/A sky130_fd_sc_hd__or3_4
XFILLER_8_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11529_ _11529_/A vssd1 vssd1 vccd1 vccd1 _11529_/Y sky130_fd_sc_hd__inv_2
XFILLER_117_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15297_ _15297_/A _15297_/B vssd1 vssd1 vccd1 vccd1 _15298_/B sky130_fd_sc_hd__or2_1
X_18085_ _20076_/CLK _18085_/D vssd1 vssd1 vccd1 vccd1 _18085_/Q sky130_fd_sc_hd__dfxtp_1
Xhold307 HWDATA[24] vssd1 vssd1 vccd1 vccd1 input54/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold318 input48/X vssd1 vssd1 vccd1 vccd1 hold318/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold329 scl_i_S5 vssd1 vssd1 vccd1 vccd1 input76/A sky130_fd_sc_hd__dlygate4sd3_1
X_17036_ _17473_/A0 _16680_/Y _17042_/S vssd1 vssd1 vccd1 vccd1 _17036_/X sky130_fd_sc_hd__mux2_1
X_14248_ _18754_/Q _14270_/B _15192_/A vssd1 vssd1 vccd1 vccd1 _14758_/C sky130_fd_sc_hd__or3_4
XANTENNA__17048__S _17545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11885__A _11892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14179_ _19109_/Q _14018_/A _16617_/A _18692_/Q _14178_/X vssd1 vssd1 vccd1 vccd1
+ _14184_/C sky130_fd_sc_hd__o221a_1
XFILLER_152_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17912__S0 _17913_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18987_ _19115_/CLK _18987_/D hold273/X vssd1 vssd1 vccd1 vccd1 _18987_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__16887__S _17473_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_239_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17938_ _19842_/CLK _17938_/D vssd1 vssd1 vccd1 vccd1 _17938_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater146 _17664_/S vssd1 vssd1 vccd1 vccd1 _17655_/S sky130_fd_sc_hd__buf_8
XFILLER_227_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater157 _17459_/S vssd1 vssd1 vccd1 vccd1 _17523_/S sky130_fd_sc_hd__buf_8
XFILLER_226_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrepeater168 _17548_/S vssd1 vssd1 vccd1 vccd1 _17545_/S sky130_fd_sc_hd__clkbuf_16
X_17869_ _17865_/X _17866_/X _17867_/X _17868_/X _18760_/Q _18761_/Q vssd1 vssd1 vccd1
+ vccd1 _17869_/X sky130_fd_sc_hd__mux4_2
Xrepeater179 _17414_/S vssd1 vssd1 vccd1 vccd1 _17482_/S sky130_fd_sc_hd__buf_6
XANTENNA__15056__B1 _15006_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19608_ _19608_/CLK _19608_/D hold355/X vssd1 vssd1 vccd1 vccd1 _19608_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_38_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17969__CLK _20123_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09090__A _10451_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19539_ _19540_/CLK _19539_/D repeater221/X vssd1 vssd1 vccd1 vccd1 _19539_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16005__C1 _16001_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17511__S _17539_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18660__RESET_B repeater210/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09223_ _18648_/Q _09238_/A _09211_/A vssd1 vssd1 vccd1 vccd1 _15713_/A sky130_fd_sc_hd__o21ai_2
XFILLER_195_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10840__A1 _19717_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09154_ _09154_/A _09156_/A _09156_/B vssd1 vssd1 vccd1 vccd1 _09154_/X sky130_fd_sc_hd__or3_2
XANTENNA__12042__B1 _11975_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_127_HCLK clkbuf_4_4_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19577_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_175_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09085_ hold237/X vssd1 vssd1 vccd1 vccd1 _10448_/A sky130_fd_sc_hd__buf_4
XFILLER_163_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12345__A1 _19173_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17903__S0 _17913_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09987_ _09987_/A _09987_/B _09987_/C vssd1 vssd1 vccd1 vccd1 _19949_/D sky130_fd_sc_hd__nor3_1
XANTENNA__16797__S _17535_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08938_ _10323_/A _08937_/Y _19857_/Q _18777_/Q vssd1 vssd1 vccd1 vccd1 _08943_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_85_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10900_ _19688_/Q _10893_/X _10863_/X _10895_/X vssd1 vssd1 vccd1 vccd1 _19688_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_84_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13515__A _18759_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11880_ _19431_/Q _11875_/X _09021_/X _11878_/X vssd1 vssd1 vccd1 vccd1 _19431_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_189_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10831_ _15336_/A _10831_/B vssd1 vssd1 vccd1 vccd1 _10840_/S sky130_fd_sc_hd__or2_2
XFILLER_16_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17421__S _17546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13550_ _13550_/A _13573_/A vssd1 vssd1 vccd1 vccd1 _13551_/B sky130_fd_sc_hd__or2_2
XFILLER_213_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12281__B1 _12102_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10762_ _19752_/Q _19751_/Q _10771_/B vssd1 vssd1 vccd1 vccd1 _10762_/X sky130_fd_sc_hd__and3_1
XFILLER_197_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12501_ _19086_/Q _12498_/X _12392_/X _12499_/X vssd1 vssd1 vccd1 vccd1 _19086_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19640__SET_B repeater258/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_213_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13481_ _13481_/A vssd1 vssd1 vccd1 vccd1 _13485_/A sky130_fd_sc_hd__inv_2
X_10693_ _10704_/B vssd1 vssd1 vccd1 vccd1 _17749_/S sky130_fd_sc_hd__inv_2
XFILLER_157_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15220_ _19721_/Q _15208_/Y _15219_/Y _10909_/A _15209_/X vssd1 vssd1 vccd1 vccd1
+ _15220_/Y sky130_fd_sc_hd__o2111ai_4
X_12432_ _19129_/Q _12427_/X _12234_/X _12428_/X vssd1 vssd1 vccd1 vccd1 _19129_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11689__B _13252_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12033__B1 _12032_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15151_ _17958_/Q _15146_/X _14705_/A _15148_/X vssd1 vssd1 vccd1 vccd1 _17958_/D
+ sky130_fd_sc_hd__a22o_1
X_12363_ _19164_/Q _12361_/X _12299_/X _12362_/X vssd1 vssd1 vccd1 vccd1 _19164_/D
+ sky130_fd_sc_hd__a22o_1
X_14102_ _18701_/Q _14101_/Y _14096_/X _14102_/C1 vssd1 vssd1 vccd1 vccd1 _18701_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_4_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11314_ _11466_/A _18967_/Q _19583_/Q _11311_/Y _11313_/X vssd1 vssd1 vccd1 vccd1
+ _11315_/D sky130_fd_sc_hd__o221a_1
X_15082_ _15082_/A _18755_/Q _15082_/C vssd1 vssd1 vccd1 vccd1 _15084_/A sky130_fd_sc_hd__or3_4
X_12294_ _19202_/Q _12290_/X _12223_/X _12291_/X vssd1 vssd1 vccd1 vccd1 _19202_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19536__RESET_B repeater221/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14033_ _14033_/A vssd1 vssd1 vccd1 vccd1 _14033_/Y sky130_fd_sc_hd__inv_2
X_18910_ _19288_/CLK _18910_/D repeater188/X vssd1 vssd1 vccd1 vccd1 _18910_/Q sky130_fd_sc_hd__dfrtp_1
X_11245_ _18996_/Q vssd1 vssd1 vccd1 vccd1 _16208_/A sky130_fd_sc_hd__inv_2
X_19890_ _20070_/CLK _19890_/D repeater206/X vssd1 vssd1 vccd1 vccd1 _19890_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_106_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18841_ _20107_/CLK _18841_/D repeater233/X vssd1 vssd1 vccd1 vccd1 _18841_/Q sky130_fd_sc_hd__dfrtp_1
X_11176_ _11191_/A vssd1 vssd1 vccd1 vccd1 _11176_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_122_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10127_ _18585_/Q _18584_/Q _15562_/A vssd1 vssd1 vccd1 vccd1 _15566_/A sky130_fd_sc_hd__or3_4
X_18772_ _19855_/CLK _18772_/D repeater265/X vssd1 vssd1 vccd1 vccd1 _18772_/Q sky130_fd_sc_hd__dfrtp_1
X_15984_ _18873_/Q vssd1 vssd1 vccd1 vccd1 _15984_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17027__A1 _19409_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17723_ _19677_/Q _19690_/Q _18510_/Q vssd1 vssd1 vccd1 vccd1 _17723_/X sky130_fd_sc_hd__mux2_1
X_10058_ _19932_/Q _10052_/C _10057_/X _10055_/A vssd1 vssd1 vccd1 vccd1 _19932_/D
+ sky130_fd_sc_hd__o211a_1
X_14935_ _20075_/Q vssd1 vssd1 vccd1 vccd1 _14935_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_209_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15038__B1 _14992_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17654_ _15619_/X _19035_/Q _17655_/S vssd1 vssd1 vccd1 vccd1 _18598_/D sky130_fd_sc_hd__mux2_1
X_14866_ _18132_/Q _14859_/A _14711_/X _14860_/A vssd1 vssd1 vccd1 vccd1 _18132_/D
+ sky130_fd_sc_hd__a22o_1
X_16605_ _16856_/X _15889_/X _16861_/X _15887_/X vssd1 vssd1 vccd1 vccd1 _16605_/X
+ sky130_fd_sc_hd__o22a_2
XANTENNA__16250__A2 _16235_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13817_ _13911_/B _13817_/B vssd1 vssd1 vccd1 vccd1 _13938_/A sky130_fd_sc_hd__or2_1
X_17585_ _15383_/X _19680_/Q _17585_/S vssd1 vssd1 vccd1 vccd1 _17585_/X sky130_fd_sc_hd__mux2_1
XFILLER_23_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14797_ _18171_/Q _14786_/A _14780_/X _14787_/A vssd1 vssd1 vccd1 vccd1 _18171_/D
+ sky130_fd_sc_hd__a22o_1
X_19324_ _19324_/CLK _19324_/D repeater213/X vssd1 vssd1 vccd1 vccd1 _19324_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_90_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17331__S _17487_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16536_ _08922_/Y _16505_/X _10234_/Y _16506_/X vssd1 vssd1 vccd1 vccd1 _16536_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12272__B1 _12086_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16538__B1 _17113_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13748_ _13748_/A vssd1 vssd1 vccd1 vccd1 _13760_/B sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_opt_3_HCLK_A clkbuf_opt_3_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19255_ _19255_/CLK _19255_/D repeater237/X vssd1 vssd1 vccd1 vccd1 _19255_/Q sky130_fd_sc_hd__dfrtp_1
X_16467_ _16467_/A _16469_/B vssd1 vssd1 vccd1 vccd1 _16467_/Y sky130_fd_sc_hd__nor2_1
X_13679_ _18774_/Q _13671_/X _13678_/X _13672_/X vssd1 vssd1 vccd1 vccd1 _18774_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18206_ _18216_/CLK _18206_/D vssd1 vssd1 vccd1 vccd1 _18206_/Q sky130_fd_sc_hd__dfxtp_1
X_15418_ _18541_/Q _13228_/B _17584_/S vssd1 vssd1 vccd1 vccd1 _15418_/X sky130_fd_sc_hd__a21o_1
XFILLER_157_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19186_ _19293_/CLK _19186_/D repeater186/X vssd1 vssd1 vccd1 vccd1 _19186_/Q sky130_fd_sc_hd__dfrtp_1
X_16398_ _18145_/Q vssd1 vssd1 vccd1 vccd1 _16398_/Y sky130_fd_sc_hd__inv_2
XANTENNA__09976__C1 _09964_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18137_ _18137_/CLK _18137_/D vssd1 vssd1 vccd1 vccd1 _18137_/Q sky130_fd_sc_hd__dfxtp_1
X_15349_ _15349_/A vssd1 vssd1 vccd1 vccd1 _15358_/A sky130_fd_sc_hd__buf_1
XFILLER_145_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18068_ _19851_/CLK _18068_/D vssd1 vssd1 vccd1 vccd1 _18068_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold137 HADDR[22] vssd1 vssd1 vccd1 vccd1 input15/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold148 input70/X vssd1 vssd1 vccd1 vccd1 hold148/X sky130_fd_sc_hd__dlygate4sd3_1
X_17019_ _15963_/X _09538_/Y _17534_/S vssd1 vssd1 vccd1 vccd1 _17019_/X sky130_fd_sc_hd__mux2_1
Xhold159 input8/X vssd1 vssd1 vccd1 vccd1 hold159/X sky130_fd_sc_hd__dlygate4sd3_1
X_09910_ _09865_/A _19349_/Q _19945_/Q _09908_/Y _09909_/X vssd1 vssd1 vccd1 vccd1
+ _09911_/D sky130_fd_sc_hd__o221a_1
XFILLER_208_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20030_ _20032_/CLK _20030_/D repeater240/X vssd1 vssd1 vccd1 vccd1 _20030_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__09085__A hold237/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09841_ _19945_/Q vssd1 vssd1 vccd1 vccd1 _09854_/A sky130_fd_sc_hd__inv_2
XANTENNA__17506__S _17566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09772_ _09772_/A vssd1 vssd1 vccd1 vccd1 _09772_/Y sky130_fd_sc_hd__inv_2
XFILLER_246_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15029__B1 _15000_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11302__A2 _18989_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18841__RESET_B repeater233/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17241__S _17546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16529__B1 _17126_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19713__SET_B repeater219/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09206_ _20068_/Q _20067_/Q _09198_/A vssd1 vssd1 vccd1 vccd1 _09206_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__12015__B1 _09039_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14555__A2 _14547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13212__C1 _13202_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09137_ _20088_/Q _09136_/Y _09131_/X vssd1 vssd1 vccd1 vccd1 _20088_/D sky130_fd_sc_hd__o21a_1
XFILLER_163_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09068_ _20103_/Q _09053_/X _09067_/X _09055_/X vssd1 vssd1 vccd1 vccd1 _20103_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_163_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11030_ _11023_/Y _17753_/S _11026_/A _11029_/Y vssd1 vssd1 vccd1 vccd1 _11030_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__17257__A1 _19078_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17416__S _17529_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16480__A2 _16638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11829__B1 _10870_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12981_ _18942_/Q _12978_/Y _12885_/B _12980_/X vssd1 vssd1 vccd1 vccd1 _18942_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_45_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14720_ _18217_/Q _14717_/X _14600_/X _14719_/X vssd1 vssd1 vccd1 vccd1 _18217_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11932_ _11841_/X _15512_/A _11932_/S vssd1 vssd1 vccd1 vccd1 _19399_/D sky130_fd_sc_hd__mux2_2
XFILLER_150_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_232_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11863_ _11863_/A vssd1 vssd1 vccd1 vccd1 _15233_/A sky130_fd_sc_hd__inv_2
X_14651_ _18252_/Q _14644_/A _09183_/X _14645_/A vssd1 vssd1 vccd1 vccd1 _18252_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17151__S _17529_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13602_ _18811_/Q _13601_/Y _13591_/X _13602_/C1 vssd1 vssd1 vccd1 vccd1 _18811_/D
+ sky130_fd_sc_hd__o211a_1
X_10814_ _17618_/X _10808_/X _19729_/Q _10810_/X vssd1 vssd1 vccd1 vccd1 _19729_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_32_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17370_ _16297_/Y _09233_/Y _19498_/Q vssd1 vssd1 vccd1 vccd1 _17370_/X sky130_fd_sc_hd__mux2_1
XPHY_3963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14582_ _14727_/A vssd1 vssd1 vccd1 vccd1 _14582_/X sky130_fd_sc_hd__clkbuf_2
X_11794_ _11801_/A vssd1 vssd1 vccd1 vccd1 _11794_/X sky130_fd_sc_hd__buf_1
XFILLER_186_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16321_ _17377_/X _15900_/A _17348_/X _15908_/A vssd1 vssd1 vccd1 vccd1 _16321_/X
+ sky130_fd_sc_hd__o22a_2
XPHY_3996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10745_ _19762_/Q _10741_/X _10448_/X _10743_/X vssd1 vssd1 vccd1 vccd1 _19762_/D
+ sky130_fd_sc_hd__a22o_1
X_13533_ _13533_/A _13604_/A vssd1 vssd1 vccd1 vccd1 _13534_/B sky130_fd_sc_hd__or2_1
XANTENNA__16990__S _17474_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19788__RESET_B repeater203/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19040_ _19041_/CLK _19040_/D repeater263/X vssd1 vssd1 vccd1 vccd1 _19040_/Q sky130_fd_sc_hd__dfrtp_1
X_13464_ _13464_/A _13481_/A vssd1 vssd1 vccd1 vccd1 _13479_/A sky130_fd_sc_hd__or2_1
XFILLER_146_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16252_ _18143_/Q vssd1 vssd1 vccd1 vccd1 _16252_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12006__B1 hold288/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10676_ _10676_/A vssd1 vssd1 vccd1 vccd1 _10676_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_9_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13203__C1 _13202_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15203_ _18639_/Q vssd1 vssd1 vccd1 vccd1 _15211_/A sky130_fd_sc_hd__inv_2
X_12415_ _19142_/Q _12412_/X _12413_/X _12414_/X vssd1 vssd1 vccd1 vccd1 _19142_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_139_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13395_ _20095_/Q _13464_/A _20119_/Q _13387_/Y vssd1 vssd1 vccd1 vccd1 _13395_/X
+ sky130_fd_sc_hd__o22a_1
X_16183_ _18238_/Q vssd1 vssd1 vccd1 vccd1 _16183_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12346_ hold282/X vssd1 vssd1 vccd1 vccd1 hold281/A sky130_fd_sc_hd__buf_4
X_15134_ _15135_/A vssd1 vssd1 vccd1 vccd1 _15134_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_154_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19370__RESET_B repeater241/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15065_ _18014_/Q _15059_/X _14810_/A _15061_/X vssd1 vssd1 vccd1 vccd1 _18014_/D
+ sky130_fd_sc_hd__a22o_1
X_19942_ _20013_/CLK _19942_/D repeater244/X vssd1 vssd1 vccd1 vccd1 _19942_/Q sky130_fd_sc_hd__dfrtp_1
X_12277_ _12277_/A vssd1 vssd1 vccd1 vccd1 _12277_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_99_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14016_ _14016_/A _14016_/B vssd1 vssd1 vccd1 vccd1 _14126_/A sky130_fd_sc_hd__or2_1
X_11228_ _11465_/A _18998_/Q _11227_/Y _19023_/Q vssd1 vssd1 vccd1 vccd1 _11228_/X
+ sky130_fd_sc_hd__o22a_1
X_19873_ _19873_/CLK _19873_/D repeater261/X vssd1 vssd1 vccd1 vccd1 _19873_/Q sky130_fd_sc_hd__dfstp_1
X_18824_ _19255_/CLK _18824_/D repeater217/X vssd1 vssd1 vccd1 vccd1 _18824_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__17326__S _17530_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11159_ _19614_/Q _11159_/B vssd1 vssd1 vccd1 vccd1 _11160_/B sky130_fd_sc_hd__or2_1
XFILLER_68_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18755_ _18869_/CLK _18755_/D repeater195/X vssd1 vssd1 vccd1 vccd1 _18755_/Q sky130_fd_sc_hd__dfrtp_2
X_15967_ _19702_/Q vssd1 vssd1 vccd1 vccd1 _15967_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19415__CLK _19984_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17706_ _15434_/X _19771_/Q _18546_/D vssd1 vssd1 vccd1 vccd1 _17706_/X sky130_fd_sc_hd__mux2_1
X_14918_ _18098_/Q _14909_/A _14868_/X _14910_/A vssd1 vssd1 vccd1 vccd1 _18098_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12493__B1 _12375_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18686_ _18686_/CLK _18686_/D hold359/X vssd1 vssd1 vccd1 vccd1 _18686_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_91_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15898_ _16634_/A vssd1 vssd1 vccd1 vccd1 _15898_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_224_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17637_ _15691_/X _19052_/Q _17655_/S vssd1 vssd1 vccd1 vccd1 _18615_/D sky130_fd_sc_hd__mux2_1
XFILLER_224_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14849_ _18144_/Q _14845_/X _14806_/X _14847_/X vssd1 vssd1 vccd1 vccd1 _18144_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_212_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17061__S _17546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17568_ _17567_/X _17914_/X _17568_/S vssd1 vssd1 vccd1 vccd1 _17568_/X sky130_fd_sc_hd__mux2_1
XANTENNA__15982__B2 _15867_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19307_ _20120_/CLK _19307_/D repeater238/X vssd1 vssd1 vccd1 vccd1 _19307_/Q sky130_fd_sc_hd__dfrtp_1
X_16519_ _17293_/X _16505_/X _17277_/X _16506_/X vssd1 vssd1 vccd1 vccd1 _16519_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_220_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17499_ _15958_/Y _15957_/Y _17564_/S vssd1 vssd1 vccd1 vccd1 _17499_/X sky130_fd_sc_hd__mux2_1
XFILLER_210_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_220_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19238_ _19282_/CLK _19238_/D repeater215/X vssd1 vssd1 vccd1 vccd1 _19238_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_192_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19458__RESET_B repeater272/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19169_ _19208_/CLK _19169_/D hold363/X vssd1 vssd1 vccd1 vccd1 _19169_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_129_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17487__A1 _12936_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16695__C1 _16694_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20013_ _20013_/CLK _20013_/D repeater242/X vssd1 vssd1 vccd1 vccd1 _20013_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17236__S _17542_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09824_ _19962_/Q vssd1 vssd1 vccd1 vccd1 _09870_/A sky130_fd_sc_hd__inv_2
XFILLER_98_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09755_ _09755_/A vssd1 vssd1 vccd1 vccd1 _09755_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12484__B1 _12236_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09686_ _19417_/Q vssd1 vssd1 vccd1 vccd1 _09686_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10530_ _10530_/A _19543_/Q _10530_/C vssd1 vssd1 vccd1 vccd1 _10531_/B sky130_fd_sc_hd__or3_1
XPHY_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16922__A0 _15963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14528__A2 _14519_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10461_ _19825_/Q vssd1 vssd1 vccd1 vccd1 _10461_/Y sky130_fd_sc_hd__inv_2
XFILLER_182_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12200_ _19253_/Q _12198_/X _12083_/X _12199_/X vssd1 vssd1 vccd1 vccd1 _19253_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_6_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13180_ _13180_/A vssd1 vssd1 vccd1 vccd1 _13180_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_202_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10392_ _19849_/Q vssd1 vssd1 vccd1 vccd1 _14256_/A sky130_fd_sc_hd__inv_2
XFILLER_124_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12131_ _12371_/A _15895_/A vssd1 vssd1 vccd1 vccd1 _12316_/B sky130_fd_sc_hd__or2_4
XANTENNA__16686__C1 _16685_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16150__A1 _15749_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12062_ _15776_/A _12066_/A vssd1 vssd1 vccd1 vccd1 _12063_/S sky130_fd_sc_hd__or2_1
XANTENNA__18312__CLK _19847_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17146__S _17536_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11013_ _10224_/X _10211_/X _10956_/C _10956_/D vssd1 vssd1 vccd1 vccd1 _11013_/X
+ sky130_fd_sc_hd__o31a_1
XANTENNA__15455__A _15479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16870_ _15963_/X _12815_/Y _17534_/S vssd1 vssd1 vccd1 vccd1 _16870_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_238_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18763__RESET_B repeater195/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15821_ _15961_/A _15821_/B vssd1 vssd1 vccd1 vccd1 _17558_/S sky130_fd_sc_hd__nor2_4
XFILLER_38_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18540_ _19825_/CLK _18540_/D repeater229/X vssd1 vssd1 vccd1 vccd1 _18540_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_246_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15752_ _19780_/Q _15751_/Y _15439_/A vssd1 vssd1 vccd1 vccd1 _18515_/D sky130_fd_sc_hd__o21ai_1
XANTENNA__11278__B2 _18994_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12475__B1 _12223_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12964_ _12964_/A _12964_/B _12964_/C _12964_/D vssd1 vssd1 vccd1 vccd1 _12965_/D
+ sky130_fd_sc_hd__or4_1
XFILLER_234_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14703_ _14703_/A vssd1 vssd1 vccd1 vccd1 _14703_/X sky130_fd_sc_hd__clkbuf_2
X_18471_ _18954_/CLK _18471_/D vssd1 vssd1 vccd1 vccd1 _18471_/Q sky130_fd_sc_hd__dfxtp_1
X_11915_ _11915_/A vssd1 vssd1 vccd1 vccd1 _11915_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_206_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15683_ _15683_/A _15683_/B vssd1 vssd1 vccd1 vccd1 _15683_/Y sky130_fd_sc_hd__nor2_1
XPHY_4450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14216__B2 _14004_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12895_ _12894_/Y _18944_/Q _19287_/Q _12887_/A vssd1 vssd1 vccd1 vccd1 _12895_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_4461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19969__RESET_B repeater274/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17422_ _17421_/X _14081_/Y _17544_/S vssd1 vssd1 vccd1 vccd1 _17422_/X sky130_fd_sc_hd__mux2_1
XANTENNA__15190__A _15190_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12227__B1 _11975_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14634_ _18264_/Q _14630_/X _09171_/X _14632_/X vssd1 vssd1 vccd1 vccd1 _18264_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11846_ _12558_/B _15774_/A vssd1 vssd1 vccd1 vccd1 _11847_/S sky130_fd_sc_hd__or2_1
XPHY_4494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17353_ _17352_/X _09853_/A _17518_/S vssd1 vssd1 vccd1 vccd1 _17353_/X sky130_fd_sc_hd__mux2_1
XFILLER_202_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11777_ hold193/X _11771_/X _19471_/Q _11772_/X vssd1 vssd1 vccd1 vccd1 hold195/A
+ sky130_fd_sc_hd__o22a_1
X_14565_ _18301_/Q _14558_/X hold330/X _14560_/X vssd1 vssd1 vccd1 vccd1 _18301_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16304_ _16302_/Y _16303_/X _15733_/Y _15850_/B vssd1 vssd1 vccd1 vccd1 _16304_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_202_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10728_ _19767_/Q _10721_/A _10423_/X _10722_/A vssd1 vssd1 vccd1 vccd1 _19767_/D
+ sky130_fd_sc_hd__a22o_1
X_13516_ _13516_/A vssd1 vssd1 vccd1 vccd1 _13516_/Y sky130_fd_sc_hd__inv_2
X_17284_ _17283_/X _15618_/A _17318_/S vssd1 vssd1 vccd1 vccd1 _17284_/X sky130_fd_sc_hd__mux2_1
XFILLER_201_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_1_0_HCLK_A clkbuf_4_1_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14496_ _18343_/Q _14491_/X _12720_/X _14493_/X vssd1 vssd1 vccd1 vccd1 _18343_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19551__RESET_B repeater274/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19023_ _19609_/CLK _19023_/D hold357/X vssd1 vssd1 vccd1 vccd1 _19023_/Q sky130_fd_sc_hd__dfrtp_2
X_16235_ _16688_/A vssd1 vssd1 vccd1 vccd1 _16235_/X sky130_fd_sc_hd__buf_2
X_13447_ _13447_/A vssd1 vssd1 vccd1 vccd1 _13447_/Y sky130_fd_sc_hd__inv_2
X_10659_ _19796_/Q _10655_/X _19700_/Q _10658_/X vssd1 vssd1 vccd1 vccd1 _18508_/D
+ sky130_fd_sc_hd__o211ai_4
XFILLER_127_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13378_ _20120_/Q _18866_/Q _20120_/Q _18866_/Q vssd1 vssd1 vccd1 vccd1 _13378_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_16166_ _18470_/Q vssd1 vssd1 vccd1 vccd1 _16166_/Y sky130_fd_sc_hd__inv_2
XFILLER_170_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15117_ _17980_/Q _15110_/X _14931_/X _15112_/X vssd1 vssd1 vccd1 vccd1 _17980_/D
+ sky130_fd_sc_hd__a22o_1
X_12329_ _19184_/Q _12327_/X _12083_/X _12328_/X vssd1 vssd1 vccd1 vccd1 _19184_/D
+ sky130_fd_sc_hd__a22o_1
X_16097_ _18125_/Q vssd1 vssd1 vccd1 vccd1 _16097_/Y sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_113_HCLK_A clkbuf_opt_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19925_ _19927_/CLK _19925_/D repeater235/X vssd1 vssd1 vccd1 vccd1 _19925_/Q sky130_fd_sc_hd__dfrtp_1
X_15048_ _15048_/A vssd1 vssd1 vccd1 vccd1 _15049_/A sky130_fd_sc_hd__inv_2
XFILLER_69_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17056__S _17542_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19856_ _19865_/CLK _19856_/D repeater265/X vssd1 vssd1 vccd1 vccd1 _19856_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_84_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18807_ _18856_/CLK _18807_/D repeater231/X vssd1 vssd1 vccd1 vccd1 _18807_/Q sky130_fd_sc_hd__dfrtp_1
X_19787_ _20089_/CLK _19787_/D repeater203/X vssd1 vssd1 vccd1 vccd1 _19787_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__16895__S _17473_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16999_ _16998_/X _09487_/A _17386_/S vssd1 vssd1 vccd1 vccd1 _16999_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09540_ _20030_/Q _09538_/Y _09465_/A _19294_/Q _09539_/X vssd1 vssd1 vccd1 vccd1
+ _09545_/C sky130_fd_sc_hd__o221a_1
X_18738_ _20051_/CLK _18738_/D repeater200/X vssd1 vssd1 vccd1 vccd1 _18738_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12466__B1 _12413_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_243_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09471_ _09471_/A _09471_/B vssd1 vssd1 vccd1 vccd1 _09609_/A sky130_fd_sc_hd__or2_1
X_18669_ _19812_/CLK _18669_/D repeater222/X vssd1 vssd1 vccd1 vccd1 _18669_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__12218__B1 _12032_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_211_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19639__RESET_B repeater257/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_212_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16643__B _16647_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10691__B _15858_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11744__A2 _11737_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_35_HCLK_A _18641_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold187_A HADDR[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_98_HCLK_A clkbuf_4_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09807_ _09807_/A _09807_/B _09807_/C vssd1 vssd1 vccd1 vccd1 _09810_/A sky130_fd_sc_hd__or3_4
XANTENNA_clkbuf_4_12_0_HCLK_A clkbuf_3_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11308__A _18969_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09738_ _09738_/A _09813_/C _09738_/C vssd1 vssd1 vccd1 vccd1 _20002_/D sky130_fd_sc_hd__nor3_1
XFILLER_216_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09669_ _09669_/A vssd1 vssd1 vccd1 vccd1 _09738_/A sky130_fd_sc_hd__inv_2
XPHY_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11700_ _19521_/Q _11691_/A _10870_/X _11692_/A vssd1 vssd1 vccd1 vccd1 _19521_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12209__B1 _12100_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12680_ _18980_/Q _12677_/X hold301/X _12678_/X vssd1 vssd1 vccd1 vccd1 _18980_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_70_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11631_ _11624_/A _11624_/B _11629_/Y _11645_/C vssd1 vssd1 vccd1 vccd1 _19554_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_230_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11562_ _11562_/A vssd1 vssd1 vccd1 vccd1 _11569_/B sky130_fd_sc_hd__inv_2
X_14350_ hold248/X vssd1 vssd1 vccd1 vccd1 _14745_/A sky130_fd_sc_hd__clkbuf_2
XPHY_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10513_ _10526_/B _19531_/Q _19532_/Q vssd1 vssd1 vccd1 vccd1 _10516_/A sky130_fd_sc_hd__or3b_1
X_13301_ _18867_/Q vssd1 vssd1 vccd1 vccd1 _13354_/A sky130_fd_sc_hd__inv_2
XANTENNA__17794__S1 _19648_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14281_ _18462_/Q _14272_/X _13674_/X _14275_/X vssd1 vssd1 vccd1 vccd1 _18462_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11978__A _14277_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11493_ _11488_/A _11488_/B _11528_/A _11489_/Y vssd1 vssd1 vccd1 vccd1 _19608_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_10_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10882__A _14277_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13232_ _18886_/Q _13231_/X _18885_/Q _17584_/S vssd1 vssd1 vccd1 vccd1 _18886_/D
+ sky130_fd_sc_hd__a22o_1
X_16020_ _18404_/Q vssd1 vssd1 vccd1 vccd1 _16020_/Y sky130_fd_sc_hd__inv_2
XFILLER_171_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10444_ _19835_/Q _10441_/X _09077_/X _10442_/X vssd1 vssd1 vccd1 vccd1 _19835_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_152_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12932__A1 _12929_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19260__CLK _20013_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13163_ _18918_/Q _13090_/Y _13091_/Y _13090_/A _13162_/X vssd1 vssd1 vccd1 vccd1
+ _18918_/D sky130_fd_sc_hd__o221a_1
X_10375_ _10375_/A vssd1 vssd1 vccd1 vccd1 _10376_/B sky130_fd_sc_hd__inv_2
X_12114_ _12121_/A vssd1 vssd1 vccd1 vccd1 _12114_/X sky130_fd_sc_hd__clkbuf_2
X_17971_ _18765_/CLK _17971_/D vssd1 vssd1 vccd1 vccd1 _17971_/Q sky130_fd_sc_hd__dfxtp_1
X_13094_ _19175_/Q vssd1 vssd1 vccd1 vccd1 _16585_/A sky130_fd_sc_hd__inv_2
X_19710_ _19720_/CLK _19710_/D repeater201/X vssd1 vssd1 vccd1 vccd1 _19710_/Q sky130_fd_sc_hd__dfstp_1
X_16922_ _15963_/X _09556_/Y _17534_/S vssd1 vssd1 vccd1 vccd1 _16922_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12045_ _19337_/Q _12043_/X _11978_/X _12044_/X vssd1 vssd1 vccd1 vccd1 _19337_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12696__B1 hold259/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12602__A _14279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19641_ _19647_/CLK _19641_/D repeater261/X vssd1 vssd1 vccd1 vccd1 _19641_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_120_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16853_ _16852_/X _13546_/A _17536_/S vssd1 vssd1 vccd1 vccd1 _16853_/X sky130_fd_sc_hd__mux2_1
XFILLER_238_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17604__S _17605_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15804_ _17945_/Q vssd1 vssd1 vccd1 vccd1 _15804_/Y sky130_fd_sc_hd__inv_2
X_19572_ _19595_/CLK _19572_/D repeater282/X vssd1 vssd1 vccd1 vccd1 _19572_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__12448__B1 _12384_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16784_ _16783_/X _09877_/A _17513_/S vssd1 vssd1 vccd1 vccd1 _16784_/X sky130_fd_sc_hd__mux2_1
XFILLER_225_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13996_ _18678_/Q vssd1 vssd1 vccd1 vccd1 _14009_/A sky130_fd_sc_hd__inv_2
XFILLER_218_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18523_ _19825_/CLK _18523_/D repeater223/X vssd1 vssd1 vccd1 vccd1 _18523_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__16728__B _16728_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15735_ _15735_/A _15735_/B vssd1 vssd1 vccd1 vccd1 _18480_/D sky130_fd_sc_hd__and2_1
X_12947_ _19263_/Q _13021_/C _12945_/Y _18924_/Q _12946_/X vssd1 vssd1 vccd1 vccd1
+ _12955_/B sky130_fd_sc_hd__o221a_1
XFILLER_18_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18454_ _19842_/CLK _18454_/D vssd1 vssd1 vccd1 vccd1 _18454_/Q sky130_fd_sc_hd__dfxtp_1
X_15666_ _15666_/A _15666_/B vssd1 vssd1 vccd1 vccd1 _15666_/Y sky130_fd_sc_hd__nor2_1
XPHY_4280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12878_ _12878_/A _12991_/A vssd1 vssd1 vccd1 vccd1 _12879_/B sky130_fd_sc_hd__or2_1
XPHY_4291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17405_ _17473_/A0 _16122_/Y _17512_/S vssd1 vssd1 vccd1 vccd1 _17405_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14617_ _14617_/A vssd1 vssd1 vccd1 vccd1 _14618_/A sky130_fd_sc_hd__inv_2
X_18385_ _18441_/CLK _18385_/D vssd1 vssd1 vccd1 vccd1 _18385_/Q sky130_fd_sc_hd__dfxtp_1
X_11829_ _19439_/Q _11800_/A _10870_/X _11801_/A vssd1 vssd1 vccd1 vccd1 _19439_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_221_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15597_ _15597_/A vssd1 vssd1 vccd1 vccd1 _15602_/B sky130_fd_sc_hd__inv_2
XPHY_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17336_ _15768_/Y _11264_/Y _17546_/S vssd1 vssd1 vccd1 vccd1 _17336_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12620__B1 _12384_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14548_ _14548_/A vssd1 vssd1 vccd1 vccd1 _14548_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_186_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17785__S1 _19646_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15165__A2 _15158_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17267_ _17486_/A0 _13137_/Y _17543_/S vssd1 vssd1 vccd1 vccd1 _17267_/X sky130_fd_sc_hd__mux2_1
X_14479_ _14479_/A vssd1 vssd1 vccd1 vccd1 _14480_/A sky130_fd_sc_hd__inv_2
X_19006_ _19595_/CLK _19006_/D hold346/A vssd1 vssd1 vccd1 vccd1 _19006_/Q sky130_fd_sc_hd__dfrtp_4
X_16218_ _19713_/Q vssd1 vssd1 vccd1 vccd1 _16218_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14373__B1 hold324/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09919__A2 _09918_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_160_HCLK clkbuf_4_0_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19515_/CLK sky130_fd_sc_hd__clkbuf_16
X_17198_ _17197_/X _11354_/Y _17493_/S vssd1 vssd1 vccd1 vccd1 _17198_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12923__A1 _12922_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16149_ _17408_/X _16148_/X _17417_/X _16003_/X vssd1 vssd1 vccd1 vccd1 _16149_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__18685__RESET_B repeater252/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19753__CLK _19900_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08971_ _13285_/A vssd1 vssd1 vccd1 vccd1 _13496_/C sky130_fd_sc_hd__inv_2
XFILLER_216_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19908_ _20006_/CLK _19908_/D repeater241/X vssd1 vssd1 vccd1 vccd1 _19908_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__09147__A3 hold344/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12687__B1 hold233/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12512__A _12528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09093__A _14791_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19839_ _19846_/CLK _19839_/D repeater270/X vssd1 vssd1 vccd1 vccd1 _19839_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_57_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17514__S _17537_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_232_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15823__A _15823_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09523_ _20032_/Q _09522_/Y _09492_/A _19322_/Q vssd1 vssd1 vccd1 vccd1 _09523_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_43_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09454_ _19921_/Q vssd1 vssd1 vccd1 vccd1 _10037_/A sky130_fd_sc_hd__inv_2
XPHY_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19473__RESET_B repeater260/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09385_ _10011_/A _19369_/Q _19912_/Q _09381_/Y _09384_/X vssd1 vssd1 vccd1 vccd1
+ _09385_/X sky130_fd_sc_hd__a221o_1
XFILLER_178_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19402__RESET_B repeater244/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17776__S1 _19646_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17550__A0 _15847_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13167__A1 _18916_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14364__B1 _14312_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17302__A0 _17486_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10160_ _19892_/Q _10154_/X _09094_/X _10156_/X vssd1 vssd1 vccd1 vccd1 _19892_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_121_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10091_ _10091_/A vssd1 vssd1 vccd1 vccd1 _10091_/Y sky130_fd_sc_hd__inv_2
XFILLER_126_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_248_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17424__S _17546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13850_ _13850_/A _13850_/B _13850_/C _13849_/X vssd1 vssd1 vccd1 vccd1 _13850_/X
+ sky130_fd_sc_hd__or4b_4
XFILLER_235_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16548__B _16583_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12801_ _19253_/Q _13553_/A _12797_/Y _18804_/Q _12800_/X vssd1 vssd1 vccd1 vccd1
+ _12808_/C sky130_fd_sc_hd__o221a_1
Xclkbuf_leaf_41_HCLK clkbuf_opt_1_HCLK/A vssd1 vssd1 vccd1 vccd1 _19808_/CLK sky130_fd_sc_hd__clkbuf_16
X_10993_ _19662_/Q _10993_/B vssd1 vssd1 vccd1 vccd1 _10993_/Y sky130_fd_sc_hd__nor2_1
XFILLER_62_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13781_ _18731_/Q vssd1 vssd1 vccd1 vccd1 _13830_/B sky130_fd_sc_hd__inv_2
XANTENNA__10877__A _14273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11102__B1 _19634_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15520_ _18573_/Q _15518_/C _18574_/Q vssd1 vssd1 vccd1 vccd1 _15520_/X sky130_fd_sc_hd__o21a_1
XFILLER_243_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12732_ _18952_/Q _12710_/A _12731_/X _12711_/A vssd1 vssd1 vccd1 vccd1 _18952_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_231_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15451_ _15453_/A _15450_/X _15571_/A vssd1 vssd1 vccd1 vccd1 _15451_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_231_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12663_ _12699_/A vssd1 vssd1 vccd1 vccd1 _12678_/A sky130_fd_sc_hd__clkbuf_2
XPHY_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14402_ _18396_/Q _14395_/A _14329_/X _14396_/A vssd1 vssd1 vccd1 vccd1 _18396_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11614_ _11573_/A _11573_/B _11617_/A _11612_/Y vssd1 vssd1 vccd1 vccd1 _19560_/D
+ sky130_fd_sc_hd__a211oi_2
X_18170_ _18869_/CLK _18170_/D vssd1 vssd1 vccd1 vccd1 _18170_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15382_ _19717_/Q _18481_/Q vssd1 vssd1 vccd1 vccd1 _15382_/X sky130_fd_sc_hd__or2_1
XPHY_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12594_ _19034_/Q _12590_/X hold267/X _12591_/X vssd1 vssd1 vccd1 vccd1 _19034_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17767__S1 _19646_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17121_ _15768_/Y _14156_/Y _17546_/S vssd1 vssd1 vccd1 vccd1 _17121_/X sky130_fd_sc_hd__mux2_1
X_14333_ _19643_/Q vssd1 vssd1 vccd1 vccd1 _14545_/B sky130_fd_sc_hd__buf_1
XANTENNA__20048__RESET_B repeater208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11545_ _19024_/Q vssd1 vssd1 vccd1 vccd1 _11570_/A sky130_fd_sc_hd__inv_2
XPHY_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14084__A _19082_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17052_ _17473_/A0 _09939_/Y _17522_/S vssd1 vssd1 vccd1 vccd1 _17052_/X sky130_fd_sc_hd__mux2_1
X_11476_ _11476_/A _11476_/B vssd1 vssd1 vccd1 vccd1 _11511_/A sky130_fd_sc_hd__or2_1
X_14264_ _18470_/Q _14258_/X _12723_/X _14260_/X vssd1 vssd1 vccd1 vccd1 _18470_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_167_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12316__B _12316_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16003_ _16633_/A vssd1 vssd1 vccd1 vccd1 _16003_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_137_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10427_ _11926_/A vssd1 vssd1 vccd1 vccd1 _10427_/X sky130_fd_sc_hd__buf_4
X_13215_ _18887_/Q _12986_/A _13215_/B1 _13176_/X vssd1 vssd1 vccd1 vccd1 _18887_/D
+ sky130_fd_sc_hd__o211a_1
X_14195_ _19099_/Q vssd1 vssd1 vccd1 vccd1 _14195_/Y sky130_fd_sc_hd__inv_2
XFILLER_136_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14107__B1 _14106_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10358_ _19861_/Q _10358_/B vssd1 vssd1 vccd1 vccd1 _10358_/Y sky130_fd_sc_hd__nor2_1
X_13146_ _19170_/Q _13071_/A _19178_/Q _13079_/A vssd1 vssd1 vccd1 vccd1 _13146_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_97_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17954_ _20076_/CLK _17954_/D vssd1 vssd1 vccd1 vccd1 _17954_/Q sky130_fd_sc_hd__dfxtp_1
X_13077_ _13077_/A _13077_/B vssd1 vssd1 vccd1 vccd1 _13184_/A sky130_fd_sc_hd__or2_1
XANTENNA__12669__B1 hold286/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10289_ _17630_/S vssd1 vssd1 vccd1 vccd1 _10771_/A sky130_fd_sc_hd__inv_2
XFILLER_111_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12028_ _12028_/A vssd1 vssd1 vccd1 vccd1 _12028_/X sky130_fd_sc_hd__buf_4
X_16905_ _16904_/X _18895_/Q _17542_/S vssd1 vssd1 vccd1 vccd1 _16905_/X sky130_fd_sc_hd__mux2_1
X_17885_ _16026_/Y _16027_/Y _16028_/Y _16029_/Y _17908_/S0 _18759_/Q vssd1 vssd1
+ vccd1 vccd1 _17885_/X sky130_fd_sc_hd__mux4_2
XFILLER_39_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19984__RESET_B repeater193/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15643__A _15643_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17334__S _17544_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19624_ _19920_/CLK _19624_/D repeater229/X vssd1 vssd1 vccd1 vccd1 _19624_/Q sky130_fd_sc_hd__dfrtp_1
X_16836_ _16835_/X _12898_/Y _17487_/S vssd1 vssd1 vccd1 vccd1 _16836_/X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_81_HCLK_A clkbuf_4_13_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19555_ _19582_/CLK _19555_/D hold348/A vssd1 vssd1 vccd1 vccd1 _19555_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_81_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16767_ _16766_/X _13383_/Y _17385_/S vssd1 vssd1 vccd1 vccd1 _16767_/X sky130_fd_sc_hd__mux2_1
XFILLER_53_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13979_ _18695_/Q vssd1 vssd1 vccd1 vccd1 _14025_/A sky130_fd_sc_hd__inv_2
XANTENNA__14259__A _14259_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18506_ _18506_/CLK hold274/X repeater233/X vssd1 vssd1 vccd1 vccd1 _18507_/D sky130_fd_sc_hd__dfrtp_1
XFILLER_18_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15718_ _19879_/Q vssd1 vssd1 vccd1 vccd1 _15718_/Y sky130_fd_sc_hd__inv_2
X_19486_ _19510_/CLK hold147/X repeater260/X vssd1 vssd1 vccd1 vccd1 _19486_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_202_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16698_ _16682_/X _16698_/B _16698_/C vssd1 vssd1 vccd1 vccd1 _16698_/Y sky130_fd_sc_hd__nand3b_4
XFILLER_33_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18437_ _18441_/CLK _18437_/D vssd1 vssd1 vccd1 vccd1 _18437_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15649_ _18605_/Q _18606_/Q _15649_/C vssd1 vssd1 vccd1 vccd1 _15654_/B sky130_fd_sc_hd__or3_1
XFILLER_61_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09170_ _20079_/Q vssd1 vssd1 vccd1 vccd1 _14705_/A sky130_fd_sc_hd__clkbuf_2
X_18368_ _19637_/CLK _18368_/D vssd1 vssd1 vccd1 vccd1 _18368_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17319_ _17486_/A0 _16369_/Y _17517_/S vssd1 vssd1 vccd1 vccd1 _17319_/X sky130_fd_sc_hd__mux2_1
XFILLER_186_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18299_ _18435_/CLK _18299_/D vssd1 vssd1 vccd1 vccd1 _18299_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09718__A2_N _19415_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18866__RESET_B repeater232/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14346__B1 _14314_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17509__S _17537_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08954_ _19855_/Q _08952_/Y _10361_/A _18780_/Q vssd1 vssd1 vccd1 vccd1 _08954_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_69_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_64_HCLK clkbuf_opt_4_HCLK/A vssd1 vssd1 vccd1 vccd1 _20120_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_56_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17244__S _17385_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_245_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09506_ _20033_/Q _16720_/A _09488_/A _19318_/Q vssd1 vssd1 vccd1 vccd1 _09506_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09437_ _19922_/Q vssd1 vssd1 vccd1 vccd1 _10038_/A sky130_fd_sc_hd__inv_2
XFILLER_188_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16384__A _19771_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13388__A1 _20095_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14585__B1 hold320/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09368_ _20009_/Q vssd1 vssd1 vccd1 vccd1 _09470_/A sky130_fd_sc_hd__inv_2
XFILLER_40_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16326__A1 _15749_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09299_ _20040_/Q _09293_/X _09108_/X _09294_/X vssd1 vssd1 vccd1 vccd1 _20040_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_20_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11330_ _11476_/A _18978_/Q _19584_/Q _11328_/Y _11329_/X vssd1 vssd1 vccd1 vccd1
+ _11331_/D sky130_fd_sc_hd__o221a_1
XFILLER_138_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15728__A _20038_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11261_ _11261_/A _11261_/B _11261_/C _11260_/X vssd1 vssd1 vccd1 vccd1 _11261_/X
+ sky130_fd_sc_hd__or4b_1
XANTENNA__17419__S _17459_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10212_ _19826_/Q vssd1 vssd1 vccd1 vccd1 _10212_/Y sky130_fd_sc_hd__inv_2
X_13000_ _13000_/A vssd1 vssd1 vccd1 vccd1 _13021_/A sky130_fd_sc_hd__clkbuf_2
X_11192_ _11192_/A vssd1 vssd1 vccd1 vccd1 _11192_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_134_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17921__S1 _19646_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10143_ _16982_/X _10136_/A _19899_/Q _10138_/X vssd1 vssd1 vccd1 vccd1 _19899_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_121_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10074_ _10074_/A vssd1 vssd1 vccd1 vccd1 _10074_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14951_ _15109_/A _15109_/B _14951_/C vssd1 vssd1 vccd1 vccd1 _14953_/A sky130_fd_sc_hd__or3_4
XFILLER_102_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13902_ _18735_/Q _13833_/Y _13834_/Y _13833_/A _13901_/X vssd1 vssd1 vccd1 vccd1
+ _18735_/D sky130_fd_sc_hd__o221a_1
XANTENNA__17154__S _17518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11991__A _12313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17670_ _15558_/X _19465_/Q _17683_/S vssd1 vssd1 vccd1 vccd1 _18582_/D sky130_fd_sc_hd__mux2_1
X_14882_ _14990_/A _15034_/B _15009_/C vssd1 vssd1 vccd1 vccd1 _14884_/A sky130_fd_sc_hd__or3_4
XFILLER_247_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10103__C _10107_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16621_ _16621_/A _16621_/B vssd1 vssd1 vccd1 vccd1 _16621_/Y sky130_fd_sc_hd__nor2_1
X_13833_ _13833_/A vssd1 vssd1 vccd1 vccd1 _13833_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16993__S _17546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19340_ _19352_/CLK _19340_/D hold373/X vssd1 vssd1 vccd1 vccd1 _19340_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_189_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16552_ _17155_/X _16505_/X _17167_/X _16506_/X vssd1 vssd1 vccd1 vccd1 _16552_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_16_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13764_ _18746_/Q _13287_/X _13748_/A _13763_/X vssd1 vssd1 vccd1 vccd1 _18746_/D
+ sky130_fd_sc_hd__a31o_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10976_ _19666_/Q _10976_/B vssd1 vssd1 vccd1 vccd1 _10976_/X sky130_fd_sc_hd__or2_1
XFILLER_16_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15503_ _15535_/A _15503_/B vssd1 vssd1 vccd1 vccd1 _15503_/Y sky130_fd_sc_hd__nor2_1
XFILLER_16_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12715_ _14806_/A _12709_/X _12714_/X _12711_/X vssd1 vssd1 vccd1 vccd1 _18958_/D
+ sky130_fd_sc_hd__a22o_1
X_19271_ _19282_/CLK _19271_/D repeater216/X vssd1 vssd1 vccd1 vccd1 _19271_/Q sky130_fd_sc_hd__dfrtp_1
X_16483_ _17565_/S _16483_/B _17564_/S vssd1 vssd1 vccd1 vccd1 _16484_/A sky130_fd_sc_hd__or3_1
XANTENNA_repeater174_A _17474_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13695_ _17760_/X vssd1 vssd1 vccd1 vccd1 _13700_/A sky130_fd_sc_hd__inv_2
XFILLER_203_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16565__B2 _15908_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18222_ _20077_/CLK _18222_/D vssd1 vssd1 vccd1 vccd1 _18222_/Q sky130_fd_sc_hd__dfxtp_1
X_15434_ _19625_/Q _11170_/B _11170_/X vssd1 vssd1 vccd1 vccd1 _15434_/X sky130_fd_sc_hd__a21bo_1
XFILLER_188_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_175_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12646_ _19002_/Q _12643_/X hold250/X _12644_/X vssd1 vssd1 vccd1 vccd1 _19002_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_203_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18153_ _18165_/CLK _18153_/D vssd1 vssd1 vccd1 vccd1 _18153_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15365_ _19781_/Q vssd1 vssd1 vccd1 vccd1 _15365_/Y sky130_fd_sc_hd__inv_2
X_12577_ _12577_/A vssd1 vssd1 vccd1 vccd1 _12577_/X sky130_fd_sc_hd__clkbuf_2
XPHY_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12327__A _12334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12051__B2 _12017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17104_ _16467_/Y _19069_/Q _17544_/S vssd1 vssd1 vccd1 vccd1 _17104_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14316_ _19642_/Q _14316_/B _15296_/B vssd1 vssd1 vccd1 vccd1 _15070_/C sky130_fd_sc_hd__or3_4
XPHY_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11528_ _11528_/A _11528_/B _11528_/C vssd1 vssd1 vccd1 vccd1 _19588_/D sky130_fd_sc_hd__nor3_1
X_18084_ _18260_/CLK _18084_/D vssd1 vssd1 vccd1 vccd1 _18084_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15296_ _15296_/A _15296_/B vssd1 vssd1 vccd1 vccd1 _15296_/Y sky130_fd_sc_hd__nor2_1
XFILLER_183_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold308 input55/X vssd1 vssd1 vccd1 vccd1 hold308/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17329__S _17536_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold319 HWDATA[19] vssd1 vssd1 vccd1 vccd1 input48/A sky130_fd_sc_hd__dlygate4sd3_1
X_17035_ _17034_/X _13084_/A _17488_/S vssd1 vssd1 vccd1 vccd1 _17035_/X sky130_fd_sc_hd__mux2_1
X_14247_ _14247_/A vssd1 vssd1 vccd1 vccd1 _15192_/A sky130_fd_sc_hd__buf_1
XFILLER_171_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11459_ _11459_/A _11592_/A vssd1 vssd1 vccd1 vccd1 _11541_/A sky130_fd_sc_hd__or2_1
XFILLER_98_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_87_HCLK clkbuf_4_13_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20032_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_152_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14178_ _19106_/Q _14015_/A _14177_/Y _18674_/Q vssd1 vssd1 vccd1 vccd1 _14178_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_112_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17912__S1 _19632_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13129_ _13128_/Y _18902_/Q _19173_/Q _13074_/A vssd1 vssd1 vccd1 vccd1 _13129_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12062__A _15776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18986_ _19608_/CLK _18986_/D hold273/X vssd1 vssd1 vccd1 vccd1 _18986_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_239_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17937_ _18869_/CLK _17937_/D vssd1 vssd1 vccd1 vccd1 _17937_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18546__CLK _19920_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17064__S _17541_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_239_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater147 _17683_/S vssd1 vssd1 vccd1 vccd1 _17696_/S sky130_fd_sc_hd__buf_6
XFILLER_226_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater158 _17544_/S vssd1 vssd1 vccd1 vccd1 _17459_/S sky130_fd_sc_hd__buf_8
X_17868_ _16191_/Y _16192_/Y _16193_/Y _16194_/Y _17908_/S0 _18759_/Q vssd1 vssd1
+ vccd1 vccd1 _17868_/X sky130_fd_sc_hd__mux4_2
Xrepeater169 _16950_/S vssd1 vssd1 vccd1 vccd1 _16946_/S sky130_fd_sc_hd__buf_6
XFILLER_94_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19607_ _19609_/CLK _19607_/D hold359/X vssd1 vssd1 vccd1 vccd1 _19607_/Q sky130_fd_sc_hd__dfrtp_4
X_16819_ _17486_/A0 _13118_/Y _17543_/S vssd1 vssd1 vccd1 vccd1 _16819_/X sky130_fd_sc_hd__mux2_1
X_17799_ _17795_/X _17796_/X _17797_/X _17798_/X _19647_/Q _19648_/Q vssd1 vssd1 vccd1
+ vccd1 _17799_/X sky130_fd_sc_hd__mux4_2
XFILLER_242_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19538_ _19545_/CLK _19538_/D repeater221/X vssd1 vssd1 vccd1 vccd1 _19538_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_62_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19941__CLK _20013_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19469_ _19470_/CLK _19469_/D repeater274/X vssd1 vssd1 vccd1 vccd1 _19469_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__15820__B _16096_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09222_ _19885_/Q vssd1 vssd1 vccd1 vccd1 _09222_/Y sky130_fd_sc_hd__inv_2
XFILLER_139_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09153_ _09153_/A vssd1 vssd1 vccd1 vccd1 _20085_/D sky130_fd_sc_hd__inv_2
XFILLER_238_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09084_ _09084_/A vssd1 vssd1 vccd1 vccd1 _09084_/X sky130_fd_sc_hd__buf_1
XFILLER_108_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16651__B _16673_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17239__S _17493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18076__CLK _18198_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17903__S1 _19632_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09986_ _09857_/B _09986_/A2 _09857_/A vssd1 vssd1 vccd1 vccd1 _09987_/C sky130_fd_sc_hd__o21a_1
XFILLER_107_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08937_ _18777_/Q vssd1 vssd1 vccd1 vccd1 _08937_/Y sky130_fd_sc_hd__inv_2
XFILLER_229_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09281__A _19498_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16795__A1 _19222_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10830_ _19700_/Q vssd1 vssd1 vccd1 vccd1 _15336_/A sky130_fd_sc_hd__inv_2
XFILLER_16_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09277__A2 _09270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10761_ _10761_/A vssd1 vssd1 vccd1 vccd1 _10771_/B sky130_fd_sc_hd__inv_2
XFILLER_197_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12500_ _19087_/Q _12498_/X _12389_/X _12499_/X vssd1 vssd1 vccd1 vccd1 _19087_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_13_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18788__RESET_B repeater260/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13480_ _18842_/Q _13479_/Y _13466_/B _13421_/X vssd1 vssd1 vccd1 vccd1 _18842_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_200_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10692_ _15854_/A _10718_/A vssd1 vssd1 vccd1 vccd1 _10704_/B sky130_fd_sc_hd__or2_4
XFILLER_157_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10874__B _14245_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18717__RESET_B repeater253/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12431_ _19130_/Q _12427_/X _12232_/X _12428_/X vssd1 vssd1 vccd1 vccd1 _19130_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_148_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15150_ _17959_/Q _15146_/X _14703_/A _15148_/X vssd1 vssd1 vccd1 vccd1 _17959_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09985__B1 _09968_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12362_ _12362_/A vssd1 vssd1 vccd1 vccd1 _12362_/X sky130_fd_sc_hd__buf_1
XFILLER_138_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14101_ _14101_/A vssd1 vssd1 vccd1 vccd1 _14101_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11792__B1 _09027_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11313_ _11487_/A _18989_/Q _19585_/Q _11312_/Y vssd1 vssd1 vccd1 vccd1 _11313_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__17149__S _17414_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15081_ _18002_/Q _15072_/A _14782_/X _15073_/A vssd1 vssd1 vccd1 vccd1 _18002_/D
+ sky130_fd_sc_hd__a22o_1
X_12293_ _19203_/Q _12290_/X _12038_/X _12291_/X vssd1 vssd1 vccd1 vccd1 _19203_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_107_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14032_ _14032_/A _14032_/B vssd1 vssd1 vccd1 vccd1 _14033_/A sky130_fd_sc_hd__or2_1
X_11244_ _19002_/Q vssd1 vssd1 vccd1 vccd1 _11244_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14730__B1 _14693_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16988__S _17493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11175_ _11175_/A _18546_/D vssd1 vssd1 vccd1 vccd1 _11191_/A sky130_fd_sc_hd__or2_4
X_18840_ _20107_/CLK _18840_/D repeater233/X vssd1 vssd1 vccd1 vccd1 _18840_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_79_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10126_ _18583_/Q _18582_/Q _10126_/C _15547_/B vssd1 vssd1 vccd1 vccd1 _15562_/A
+ sky130_fd_sc_hd__or4_4
XANTENNA__08960__B2 _08959_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18771_ _19842_/CLK _18771_/D repeater271/X vssd1 vssd1 vccd1 vccd1 _18771_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_output141_A _19814_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15983_ _19766_/Q vssd1 vssd1 vccd1 vccd1 _15983_/Y sky130_fd_sc_hd__inv_2
XFILLER_121_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17722_ _19678_/Q _19691_/Q _18510_/Q vssd1 vssd1 vccd1 vccd1 _17722_/X sky130_fd_sc_hd__mux2_1
X_10057_ _10057_/A vssd1 vssd1 vccd1 vccd1 _10057_/X sky130_fd_sc_hd__clkbuf_2
X_14934_ _18092_/Q _14922_/A _14933_/X _14923_/A vssd1 vssd1 vccd1 vccd1 _18092_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_209_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17653_ _15623_/X _19036_/Q _17655_/S vssd1 vssd1 vccd1 vccd1 _18599_/D sky130_fd_sc_hd__mux2_1
X_14865_ _18133_/Q _14858_/X _14709_/X _14860_/X vssd1 vssd1 vccd1 vccd1 _18133_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_224_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17612__S _17614_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16604_ _17243_/X _16573_/X _17236_/X _16574_/X _16603_/X vssd1 vssd1 vccd1 vccd1
+ _16607_/B sky130_fd_sc_hd__o221a_4
XFILLER_217_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13816_ _13909_/C _13941_/A vssd1 vssd1 vccd1 vccd1 _13817_/B sky130_fd_sc_hd__or2_1
XANTENNA__14797__B1 _14780_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17584_ _18528_/Q _15390_/Y _17584_/S vssd1 vssd1 vccd1 vccd1 _17584_/X sky130_fd_sc_hd__mux2_1
X_14796_ _18172_/Q _14786_/A hold263/X _14787_/A vssd1 vssd1 vccd1 vccd1 _18172_/D
+ sky130_fd_sc_hd__a22o_1
X_19323_ _19324_/CLK _19323_/D repeater213/X vssd1 vssd1 vccd1 vccd1 _19323_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_44_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16535_ _19038_/Q vssd1 vssd1 vccd1 vccd1 _16535_/Y sky130_fd_sc_hd__inv_2
X_13747_ _18870_/Q _15191_/A vssd1 vssd1 vccd1 vccd1 _13748_/A sky130_fd_sc_hd__or2_2
XFILLER_44_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16538__B2 _15908_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10959_ _10959_/A _11001_/A vssd1 vssd1 vccd1 vccd1 _10999_/B sky130_fd_sc_hd__nor2_1
XFILLER_189_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19254_ _19324_/CLK _19254_/D repeater237/X vssd1 vssd1 vccd1 vccd1 _19254_/Q sky130_fd_sc_hd__dfrtp_4
X_16466_ _16466_/A _16469_/B vssd1 vssd1 vccd1 vccd1 _16466_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__17830__S0 _17918_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_231_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13678_ _13678_/A vssd1 vssd1 vccd1 vccd1 _13678_/X sky130_fd_sc_hd__clkbuf_4
X_18205_ _18460_/CLK _18205_/D vssd1 vssd1 vccd1 vccd1 _18205_/Q sky130_fd_sc_hd__dfxtp_1
X_15417_ _15419_/A _17572_/X vssd1 vssd1 vccd1 vccd1 _18540_/D sky130_fd_sc_hd__and2_1
XPHY_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12629_ _12629_/A vssd1 vssd1 vccd1 vccd1 _12629_/X sky130_fd_sc_hd__clkbuf_2
X_19185_ _19293_/CLK _19185_/D repeater187/X vssd1 vssd1 vccd1 vccd1 _19185_/Q sky130_fd_sc_hd__dfrtp_4
X_16397_ _15846_/A _16379_/X _15859_/A _16388_/X _16396_/X vssd1 vssd1 vccd1 vccd1
+ _16397_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_129_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18136_ _18137_/CLK _18136_/D vssd1 vssd1 vccd1 vccd1 _18136_/Q sky130_fd_sc_hd__dfxtp_1
X_15348_ _18496_/Q _14226_/B _14227_/B vssd1 vssd1 vccd1 vccd1 _15348_/X sky130_fd_sc_hd__a21bo_1
XFILLER_184_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16471__B _16544_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17059__S _17385_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18067_ _18142_/CLK _18067_/D vssd1 vssd1 vccd1 vccd1 _18067_/Q sky130_fd_sc_hd__dfxtp_1
X_15279_ _10908_/A _15278_/X _15227_/Y _15213_/A vssd1 vssd1 vccd1 vccd1 _15326_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_172_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold138 hold138/A vssd1 vssd1 vccd1 vccd1 hold138/X sky130_fd_sc_hd__dlygate4sd3_1
X_17018_ _16651_/Y _15667_/Y _17318_/S vssd1 vssd1 vccd1 vccd1 _17018_/X sky130_fd_sc_hd__mux2_2
Xhold149 HWRITE vssd1 vssd1 vccd1 vccd1 input70/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14721__B1 _14604_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16898__S _17512_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09840_ _19946_/Q vssd1 vssd1 vccd1 vccd1 _09855_/A sky130_fd_sc_hd__inv_2
XANTENNA__17897__S0 _17908_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09771_ _09750_/A _09750_/B _09767_/X _09769_/Y vssd1 vssd1 vccd1 vccd1 _19994_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_246_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18969_ _19137_/CLK _18969_/D hold348/X vssd1 vssd1 vccd1 vccd1 _18969_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_101_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17522__S _17522_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_242_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14788__B1 _14745_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_242_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16646__B _16647_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16529__B2 _16235_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17821__S0 _17918_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_210_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18810__RESET_B repeater217/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09205_ _09205_/A _09205_/B vssd1 vssd1 vccd1 vccd1 _09205_/Y sky130_fd_sc_hd__nor2_1
XFILLER_148_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09136_ _15322_/A _09136_/B vssd1 vssd1 vccd1 vccd1 _09136_/Y sky130_fd_sc_hd__nor2_1
XFILLER_182_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09067_ _12032_/A vssd1 vssd1 vccd1 vccd1 _09067_/X sky130_fd_sc_hd__buf_4
XFILLER_136_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_4_8_0_HCLK clkbuf_4_9_0_HCLK/A vssd1 vssd1 vccd1 vccd1 _18641_/CLK sky130_fd_sc_hd__clkbuf_1
XFILLER_150_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17888__S0 _17908_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_238_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18861__CLK _18866_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16465__B1 _15859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19987__CLK _19992_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08942__B2 _08941_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09969_ _19960_/Q _09967_/Y _09968_/X _09869_/B vssd1 vssd1 vccd1 vccd1 _19960_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_103_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20089_ _20089_/CLK _20089_/D repeater204/X vssd1 vssd1 vccd1 vccd1 _20089_/Q sky130_fd_sc_hd__dfrtp_1
X_12980_ _12980_/A vssd1 vssd1 vccd1 vccd1 _12980_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__11829__B2 _11801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_245_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11931_ _11933_/A _12183_/B vssd1 vssd1 vccd1 vccd1 _11932_/S sky130_fd_sc_hd__or2_1
XPHY_4610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17432__S _17567_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14650_ _18253_/Q _14643_/X _09180_/X _14645_/X vssd1 vssd1 vccd1 vccd1 _18253_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_205_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11862_ _11862_/A vssd1 vssd1 vccd1 vccd1 _11862_/Y sky130_fd_sc_hd__inv_2
XFILLER_232_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13601_ _13601_/A vssd1 vssd1 vccd1 vccd1 _13601_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10813_ _17617_/X _10808_/X _19730_/Q _10810_/X vssd1 vssd1 vccd1 vccd1 _19730_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12254__A1 _10954_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14581_ _18293_/Q _14572_/X _14580_/X _14574_/X vssd1 vssd1 vccd1 vccd1 _18293_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_14_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11793_ _11800_/A vssd1 vssd1 vccd1 vccd1 _11793_/X sky130_fd_sc_hd__buf_1
XANTENNA__10885__A _14279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16320_ _17370_/X _15884_/A _17369_/X _15915_/A vssd1 vssd1 vccd1 vccd1 _16320_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_3986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13532_ _13532_/A _13532_/B vssd1 vssd1 vccd1 vccd1 _13604_/A sky130_fd_sc_hd__or2_1
XANTENNA__19367__CLK _20091_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10744_ _19763_/Q _10741_/X _10446_/X _10743_/X vssd1 vssd1 vccd1 vccd1 _19763_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17812__S0 _17918_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16251_ _15846_/X _16225_/X _15859_/X _16233_/X _16250_/X vssd1 vssd1 vccd1 vccd1
+ _16251_/Y sky130_fd_sc_hd__o221ai_4
XANTENNA__12006__A1 _19360_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13463_ _13483_/A _13483_/B _13463_/C vssd1 vssd1 vccd1 vccd1 _13481_/A sky130_fd_sc_hd__or3_1
XFILLER_13_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10675_ _17738_/X _10669_/X _19787_/Q _10670_/X vssd1 vssd1 vccd1 vccd1 _19787_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16572__A _16682_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15202_ _15233_/B vssd1 vssd1 vccd1 vccd1 _15202_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12414_ _12428_/A vssd1 vssd1 vccd1 vccd1 _12414_/X sky130_fd_sc_hd__buf_1
XFILLER_139_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16182_ _18254_/Q vssd1 vssd1 vccd1 vccd1 _16182_/Y sky130_fd_sc_hd__inv_2
X_13394_ _20097_/Q vssd1 vssd1 vccd1 vccd1 _13394_/Y sky130_fd_sc_hd__clkinvlp_2
XFILLER_126_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15133_ _15169_/A _15196_/A vssd1 vssd1 vccd1 vccd1 _15135_/A sky130_fd_sc_hd__or2_2
XFILLER_126_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12345_ _19173_/Q _12341_/X _12344_/X _12342_/X vssd1 vssd1 vccd1 vccd1 _19173_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_127_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15064_ _18015_/Q _15059_/X _14808_/A _15061_/X vssd1 vssd1 vccd1 vccd1 _18015_/D
+ sky130_fd_sc_hd__a22o_1
X_19941_ _20013_/CLK _19941_/D repeater243/X vssd1 vssd1 vccd1 vccd1 _19941_/Q sky130_fd_sc_hd__dfrtp_1
X_12276_ _12276_/A vssd1 vssd1 vccd1 vccd1 _12276_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_175_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14015_ _14015_/A _14129_/A vssd1 vssd1 vccd1 vccd1 _14016_/B sky130_fd_sc_hd__or2_2
X_11227_ _19609_/Q vssd1 vssd1 vccd1 vccd1 _11227_/Y sky130_fd_sc_hd__inv_2
XFILLER_141_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19872_ _20059_/CLK _19872_/D repeater197/X vssd1 vssd1 vccd1 vccd1 _19872_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__17879__S0 _18760_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18823_ _18827_/CLK _18823_/D repeater217/X vssd1 vssd1 vccd1 vccd1 _18823_/Q sky130_fd_sc_hd__dfrtp_1
X_11158_ _19613_/Q _11158_/B vssd1 vssd1 vccd1 vccd1 _11159_/B sky130_fd_sc_hd__or2_1
XFILLER_1_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10109_ _19398_/Q vssd1 vssd1 vccd1 vccd1 _10109_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15966_ _19026_/Q vssd1 vssd1 vccd1 vccd1 _15966_/Y sky130_fd_sc_hd__inv_2
X_11089_ _14255_/A vssd1 vssd1 vccd1 vccd1 _15295_/B sky130_fd_sc_hd__inv_2
X_18754_ _18869_/CLK _18754_/D repeater195/X vssd1 vssd1 vccd1 vccd1 _18754_/Q sky130_fd_sc_hd__dfrtp_4
Xclkbuf_leaf_117_HCLK clkbuf_opt_0_HCLK/A vssd1 vssd1 vccd1 vccd1 _19609_/CLK sky130_fd_sc_hd__clkbuf_16
X_17705_ _15435_/X _19772_/Q _18546_/D vssd1 vssd1 vccd1 vccd1 _17705_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14917_ _18099_/Q _14909_/A _14713_/X _14910_/A vssd1 vssd1 vccd1 vccd1 _18099_/D
+ sky130_fd_sc_hd__a22o_1
X_18685_ _18686_/CLK _18685_/D repeater252/X vssd1 vssd1 vccd1 vccd1 _18685_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_63_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13690__B1 _13680_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15897_ _15897_/A vssd1 vssd1 vccd1 vccd1 _16634_/A sky130_fd_sc_hd__buf_2
XANTENNA__17342__S _17566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_224_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17636_ _15695_/Y _19053_/Q _17664_/S vssd1 vssd1 vccd1 vccd1 _18616_/D sky130_fd_sc_hd__mux2_1
X_14848_ _18145_/Q _14845_/X _14802_/X _14847_/X vssd1 vssd1 vccd1 vccd1 _18145_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_224_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16466__B _16469_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17567_ _17566_/X _11153_/Y _17567_/S vssd1 vssd1 vccd1 vccd1 _17567_/X sky130_fd_sc_hd__mux2_1
X_14779_ _18180_/Q _14772_/A _14727_/X _14773_/A vssd1 vssd1 vccd1 vccd1 _18180_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_189_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_136_HCLK_A clkbuf_4_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19306_ _20115_/CLK _19306_/D repeater238/X vssd1 vssd1 vccd1 vccd1 _19306_/Q sky130_fd_sc_hd__dfrtp_1
X_16518_ _19036_/Q vssd1 vssd1 vccd1 vccd1 _16518_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17803__S0 _17918_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17498_ _17497_/X _19875_/Q _19497_/Q vssd1 vssd1 vccd1 vccd1 _17498_/X sky130_fd_sc_hd__mux2_1
XFILLER_220_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16449_ _19763_/Q vssd1 vssd1 vccd1 vccd1 _16449_/Y sky130_fd_sc_hd__inv_2
X_19237_ _19282_/CLK _19237_/D repeater216/X vssd1 vssd1 vccd1 vccd1 _19237_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_31_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16931__A1 hold196/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19168_ _19208_/CLK _19168_/D hold363/X vssd1 vssd1 vccd1 vccd1 _19168_/Q sky130_fd_sc_hd__dfrtp_2
X_18119_ _18145_/CLK _18119_/D vssd1 vssd1 vccd1 vccd1 _18119_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19099_ _19585_/CLK _19099_/D repeater252/X vssd1 vssd1 vccd1 vccd1 _19099_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_145_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09096__A hold332/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19427__RESET_B repeater271/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15826__A _15826_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14170__A1 _19111_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17517__S _17517_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20012_ _20013_/CLK _20012_/D repeater242/X vssd1 vssd1 vccd1 vccd1 _20012_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_87_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09823_ _19963_/Q vssd1 vssd1 vccd1 vccd1 _09871_/A sky130_fd_sc_hd__inv_2
XFILLER_101_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09754_ _09754_/A _09761_/A vssd1 vssd1 vccd1 vccd1 _09755_/A sky130_fd_sc_hd__or2_2
XFILLER_228_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09685_ _19411_/Q vssd1 vssd1 vccd1 vccd1 _09685_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16657__A _19084_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13681__B1 _13680_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17252__S _17482_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15186__B1 _10451_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_58_HCLK_A clkbuf_4_12_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10460_ _19824_/Q _19823_/Q _10460_/C vssd1 vssd1 vccd1 vccd1 _10462_/A sky130_fd_sc_hd__or3_1
XFILLER_148_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_182_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09119_ _13494_/A _15321_/B vssd1 vssd1 vccd1 vccd1 _09120_/A sky130_fd_sc_hd__or2_1
X_10391_ _17748_/X vssd1 vssd1 vccd1 vccd1 _10404_/A sky130_fd_sc_hd__inv_2
XFILLER_109_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19850__RESET_B repeater258/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12130_ _12130_/A _12130_/B _12130_/C vssd1 vssd1 vccd1 vccd1 _15895_/A sky130_fd_sc_hd__or3_4
XFILLER_191_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_190_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17427__S _19498_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12061_ _11991_/X _19328_/Q _12061_/S vssd1 vssd1 vccd1 vccd1 _19328_/D sky130_fd_sc_hd__mux2_1
XFILLER_151_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11012_ _11012_/A vssd1 vssd1 vccd1 vccd1 _19657_/D sky130_fd_sc_hd__inv_2
XFILLER_132_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15820_ _17937_/Q _16096_/B vssd1 vssd1 vccd1 vccd1 _15820_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__13256__A _18751_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15751_ _18515_/Q vssd1 vssd1 vccd1 vccd1 _15751_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12963_ _18948_/Q _12890_/B _12962_/X _12891_/B vssd1 vssd1 vccd1 vccd1 _18948_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_246_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17162__S _17385_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14702_ _18225_/Q _14698_/X _14699_/X _14701_/X vssd1 vssd1 vccd1 vccd1 _18225_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_45_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18470_ _18473_/CLK _18470_/D vssd1 vssd1 vccd1 vccd1 _18470_/Q sky130_fd_sc_hd__dfxtp_1
X_11914_ _11914_/A vssd1 vssd1 vccd1 vccd1 _11914_/X sky130_fd_sc_hd__clkbuf_2
X_15682_ _15686_/B vssd1 vssd1 vccd1 vccd1 _15688_/B sky130_fd_sc_hd__inv_2
XPHY_4440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12894_ _19287_/Q vssd1 vssd1 vccd1 vccd1 _12894_/Y sky130_fd_sc_hd__inv_2
XPHY_4451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17421_ _15768_/Y _14168_/Y _17546_/S vssd1 vssd1 vccd1 vccd1 _17421_/X sky130_fd_sc_hd__mux2_1
XPHY_4462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14633_ _18265_/Q _14630_/X _09168_/X _14632_/X vssd1 vssd1 vccd1 vccd1 _18265_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18757__CLK _19900_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11845_ _12372_/A vssd1 vssd1 vccd1 vccd1 _15774_/A sky130_fd_sc_hd__buf_4
XPHY_4484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output104_A _16151_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17352_ _17351_/X _09714_/Y _17517_/S vssd1 vssd1 vccd1 vccd1 _17352_/X sky130_fd_sc_hd__mux2_1
XFILLER_214_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14564_ _18302_/Q _14558_/X _14509_/X _14560_/X vssd1 vssd1 vccd1 vccd1 _18302_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_60_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11776_ hold202/X _11771_/X _19472_/Q _11772_/X vssd1 vssd1 vccd1 vccd1 hold204/A
+ sky130_fd_sc_hd__o22a_1
XPHY_3794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16303_ _16303_/A vssd1 vssd1 vccd1 vccd1 _16303_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__11986__B1 _11924_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13515_ _18759_/Q vssd1 vssd1 vccd1 vccd1 _13704_/A sky130_fd_sc_hd__inv_2
X_10727_ _19768_/Q _10720_/X _10421_/X _10722_/X vssd1 vssd1 vccd1 vccd1 _19768_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_158_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17283_ _17473_/A0 _16503_/Y _17473_/S vssd1 vssd1 vccd1 vccd1 _17283_/X sky130_fd_sc_hd__mux2_1
XANTENNA__15177__B1 _10715_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16913__A1 _20113_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14495_ _18344_/Q _14491_/X _12717_/X _14493_/X vssd1 vssd1 vccd1 vccd1 _18344_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_202_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19022_ _19608_/CLK _19022_/D hold357/X vssd1 vssd1 vccd1 vccd1 _19022_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__13188__C1 _13176_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16234_ _16234_/A vssd1 vssd1 vccd1 vccd1 _16688_/A sky130_fd_sc_hd__buf_2
X_13446_ _13431_/D _13346_/B _13442_/Y _13445_/X vssd1 vssd1 vccd1 vccd1 _18859_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_186_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10658_ _10658_/A _18488_/D _10658_/C vssd1 vssd1 vccd1 vccd1 _10658_/X sky130_fd_sc_hd__or3_4
XFILLER_70_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16165_ _18406_/Q vssd1 vssd1 vccd1 vccd1 _16165_/Y sky130_fd_sc_hd__inv_2
X_13377_ _20100_/Q vssd1 vssd1 vccd1 vccd1 _13377_/Y sky130_fd_sc_hd__inv_2
X_10589_ _19798_/Q _10589_/B _10589_/C vssd1 vssd1 vccd1 vccd1 _10942_/A sky130_fd_sc_hd__nor3_4
XFILLER_182_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12335__A _12335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19591__RESET_B hold346/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16677__B1 _17060_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15116_ _17981_/Q _15110_/X _14929_/X _15112_/X vssd1 vssd1 vccd1 vccd1 _17981_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_170_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12328_ _12335_/A vssd1 vssd1 vccd1 vccd1 _12328_/X sky130_fd_sc_hd__buf_1
XFILLER_126_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16096_ _18245_/Q _16096_/B vssd1 vssd1 vccd1 vccd1 _16096_/Y sky130_fd_sc_hd__nor2_1
XFILLER_141_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17337__S _17459_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19924_ _19927_/CLK _19924_/D repeater230/X vssd1 vssd1 vccd1 vccd1 _19924_/Q sky130_fd_sc_hd__dfrtp_1
X_15047_ _15048_/A vssd1 vssd1 vccd1 vccd1 _15047_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_79_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12259_ _12298_/A vssd1 vssd1 vccd1 vccd1 _12276_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_69_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12163__B1 _12032_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19855_ _19855_/CLK _19855_/D repeater265/X vssd1 vssd1 vccd1 vccd1 _19855_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_110_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11910__B1 _11909_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18806_ _18856_/CLK _18806_/D repeater231/X vssd1 vssd1 vccd1 vccd1 _18806_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_84_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12070__A _12121_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19786_ _20057_/CLK _19786_/D repeater203/X vssd1 vssd1 vccd1 vccd1 _19786_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_228_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16998_ _16997_/X _09460_/Y _17385_/S vssd1 vssd1 vccd1 vccd1 _16998_/X sky130_fd_sc_hd__mux2_1
XFILLER_209_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18737_ _20051_/CLK _18737_/D repeater206/X vssd1 vssd1 vccd1 vccd1 _18737_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_243_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13663__B1 hold239/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15949_ _18075_/Q vssd1 vssd1 vccd1 vccd1 _15949_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17072__S _17548_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09470_ _09470_/A _09612_/A vssd1 vssd1 vccd1 vccd1 _09471_/B sky130_fd_sc_hd__or2_1
XFILLER_52_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18668_ _19812_/CLK _18668_/D repeater222/X vssd1 vssd1 vccd1 vccd1 _18668_/Q sky130_fd_sc_hd__dfstp_1
X_17619_ _20053_/Q _19727_/Q _17621_/S vssd1 vssd1 vccd1 vccd1 _17619_/X sky130_fd_sc_hd__mux2_1
X_18599_ _19865_/CLK _18599_/D repeater267/X vssd1 vssd1 vccd1 vccd1 _18599_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_211_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09095__B1 _09094_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14725__A _14793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10952__A1 hold148/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17247__S _17518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12154__B1 _12100_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17093__A0 _15768_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11901__B1 _09058_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09806_ _19976_/Q _09809_/A _09803_/A _09731_/X vssd1 vssd1 vccd1 vccd1 _19976_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_59_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16840__A0 _17473_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09737_ _09668_/C _09757_/B _09668_/A vssd1 vssd1 vccd1 vccd1 _09738_/C sky130_fd_sc_hd__o21a_1
XFILLER_39_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09668_ _09668_/A _09807_/B _09668_/C vssd1 vssd1 vccd1 vccd1 _09669_/A sky130_fd_sc_hd__or3_1
XFILLER_27_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09599_ _20017_/Q _09598_/Y _09585_/X _09478_/B vssd1 vssd1 vccd1 vccd1 _20017_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17710__S _18546_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11630_ _19555_/Q _11629_/Y _11626_/B _11563_/X vssd1 vssd1 vccd1 vccd1 _19555_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11968__B1 _09067_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11561_ _11561_/A _11639_/B _11561_/C vssd1 vssd1 vccd1 vccd1 _11562_/A sky130_fd_sc_hd__or3_1
XPHY_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13300_ _13289_/Y _17758_/X _13287_/X _13299_/X vssd1 vssd1 vccd1 vccd1 _18869_/D
+ sky130_fd_sc_hd__o22ai_1
XANTENNA__13709__A1 _18761_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10512_ _19545_/Q _19530_/Q _19529_/Q _10521_/C vssd1 vssd1 vccd1 vccd1 _10526_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_155_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14280_ _18463_/Q _14272_/X _14279_/X _14275_/X vssd1 vssd1 vccd1 vccd1 _18463_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_rebuffer38_A _19418_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11492_ _11523_/A vssd1 vssd1 vccd1 vccd1 _11528_/A sky130_fd_sc_hd__buf_2
XPHY_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13231_ _13231_/A vssd1 vssd1 vccd1 vccd1 _13231_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_40_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19405__CLK _19984_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10443_ _19836_/Q _10441_/X _09075_/X _10442_/X vssd1 vssd1 vccd1 vccd1 _19836_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_156_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12393__B1 _12392_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13162_ _13180_/A vssd1 vssd1 vccd1 vccd1 _13162_/X sky130_fd_sc_hd__clkbuf_2
X_10374_ _10374_/A vssd1 vssd1 vccd1 vccd1 _19857_/D sky130_fd_sc_hd__inv_2
XFILLER_123_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17157__S _17535_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12113_ _19306_/Q _12106_/X _12032_/X _12108_/X vssd1 vssd1 vccd1 vccd1 _19306_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_124_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11994__A _15774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17970_ _20123_/CLK _17970_/D vssd1 vssd1 vccd1 vccd1 _17970_/Q sky130_fd_sc_hd__dfxtp_1
X_13093_ _19166_/Q vssd1 vssd1 vccd1 vccd1 _16468_/A sky130_fd_sc_hd__inv_2
XANTENNA__12145__B1 _12083_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16921_ _16920_/X _15664_/Y _17318_/S vssd1 vssd1 vccd1 vccd1 _16921_/X sky130_fd_sc_hd__mux2_1
X_12044_ _12044_/A vssd1 vssd1 vccd1 vccd1 _12044_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_49_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12696__A1 _18968_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16996__S _17318_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13893__B1 _19222_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17084__A0 _15768_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19640_ _19849_/CLK _19640_/D repeater258/X vssd1 vssd1 vccd1 vccd1 _19640_/Q sky130_fd_sc_hd__dfstp_1
X_16852_ _16851_/X _13380_/Y _17535_/S vssd1 vssd1 vccd1 vccd1 _16852_/X sky130_fd_sc_hd__mux2_1
XFILLER_120_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18913__RESET_B repeater188/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15803_ _18090_/Q vssd1 vssd1 vccd1 vccd1 _15803_/Y sky130_fd_sc_hd__inv_2
XFILLER_225_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19571_ _19576_/CLK _19571_/D repeater282/X vssd1 vssd1 vccd1 vccd1 _19571_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_77_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16783_ _16782_/X _09710_/Y _17512_/S vssd1 vssd1 vccd1 vccd1 _16783_/X sky130_fd_sc_hd__mux2_1
X_13995_ _18679_/Q vssd1 vssd1 vccd1 vccd1 _14010_/A sky130_fd_sc_hd__inv_2
XFILLER_19_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18522_ _19814_/CLK _18522_/D repeater223/X vssd1 vssd1 vccd1 vccd1 _18522_/Q sky130_fd_sc_hd__dfrtp_1
X_15734_ _19724_/Q _15733_/Y _15384_/A vssd1 vssd1 vccd1 vccd1 _18477_/D sky130_fd_sc_hd__o21ai_1
XFILLER_46_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12946_ _19279_/Q _12878_/A _19267_/Q _13003_/A vssd1 vssd1 vccd1 vccd1 _12946_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__17387__A1 _19266_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15665_ _18609_/Q _15661_/A _15661_/B _15664_/Y _15661_/Y vssd1 vssd1 vccd1 vccd1
+ _15666_/B sky130_fd_sc_hd__o32a_1
X_18453_ _18460_/CLK _18453_/D vssd1 vssd1 vccd1 vccd1 _18453_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12877_ _12877_/A _12877_/B vssd1 vssd1 vccd1 vccd1 _12991_/A sky130_fd_sc_hd__or2_1
XPHY_4270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17404_ _17403_/X _17874_/X _17568_/S vssd1 vssd1 vccd1 vccd1 _17404_/X sky130_fd_sc_hd__mux2_2
X_14616_ _14617_/A vssd1 vssd1 vccd1 vccd1 _14616_/X sky130_fd_sc_hd__clkbuf_2
X_18384_ _19637_/CLK _18384_/D vssd1 vssd1 vccd1 vccd1 _18384_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11828_ _19440_/Q _11800_/A _10868_/X _11801_/A vssd1 vssd1 vccd1 vccd1 _19440_/D
+ sky130_fd_sc_hd__a22o_1
X_15596_ _18593_/Q vssd1 vssd1 vccd1 vccd1 _15598_/A sky130_fd_sc_hd__inv_2
XANTENNA__17139__A1 _18974_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11959__B1 hold317/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17335_ _17334_/X _13872_/Y _17545_/S vssd1 vssd1 vccd1 vccd1 _17335_/X sky130_fd_sc_hd__mux2_1
XANTENNA__18662__D hold312/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14547_ _14547_/A vssd1 vssd1 vccd1 vccd1 _14548_/A sky130_fd_sc_hd__inv_2
XFILLER_202_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11759_ hold156/X _11757_/X _19485_/Q _11758_/X vssd1 vssd1 vccd1 vccd1 hold158/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_41_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17266_ _17265_/X _09474_/A _17414_/S vssd1 vssd1 vccd1 vccd1 _17266_/X sky130_fd_sc_hd__mux2_2
X_14478_ _14479_/A vssd1 vssd1 vccd1 vccd1 _14478_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_leaf_41_HCLK_A clkbuf_opt_1_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16217_ _19029_/Q _17473_/S vssd1 vssd1 vccd1 vccd1 _16217_/Y sky130_fd_sc_hd__nand2_1
X_19005_ _19595_/CLK _19005_/D hold346/A vssd1 vssd1 vccd1 vccd1 _19005_/Q sky130_fd_sc_hd__dfrtp_1
X_13429_ _13429_/A _13429_/B _13429_/C _13429_/D vssd1 vssd1 vccd1 vccd1 _13430_/D
+ sky130_fd_sc_hd__or4_4
X_17197_ _15768_/Y _11253_/Y _17546_/S vssd1 vssd1 vccd1 vccd1 _17197_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16148_ _16238_/A vssd1 vssd1 vccd1 vccd1 _16148_/X sky130_fd_sc_hd__buf_2
XFILLER_154_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17311__A1 _17839_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17067__S _17529_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08970_ _08970_/A _08970_/B _08970_/C _08970_/D vssd1 vssd1 vccd1 vccd1 _13285_/A
+ sky130_fd_sc_hd__and4_4
X_16079_ _18021_/Q vssd1 vssd1 vccd1 vccd1 _16079_/Y sky130_fd_sc_hd__inv_2
XFILLER_170_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_216_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19907_ _20006_/CLK _19907_/D repeater241/X vssd1 vssd1 vccd1 vccd1 _19907_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_229_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19838_ _19841_/CLK _19838_/D repeater271/X vssd1 vssd1 vccd1 vccd1 _19838_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_84_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16822__A0 _15963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10162__A2 _10155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput1 input1/A vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_1
X_19769_ _19822_/CLK _19769_/D repeater228/X vssd1 vssd1 vccd1 vccd1 _19769_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_232_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09522_ _19322_/Q vssd1 vssd1 vccd1 vccd1 _09522_/Y sky130_fd_sc_hd__inv_2
XFILLER_232_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09453_ _19381_/Q vssd1 vssd1 vccd1 vccd1 _09453_/Y sky130_fd_sc_hd__inv_2
XFILLER_80_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17530__S _17530_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09068__B1 _09067_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09384_ _10082_/A _19370_/Q _10009_/A _19394_/Q vssd1 vssd1 vccd1 vccd1 _09384_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_101_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19428__CLK _19976_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16889__A0 _15768_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19442__RESET_B repeater193/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12127__B1 _11922_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold297_A HWDATA[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10090_ _10088_/A _10088_/B _10079_/A _10088_/Y vssd1 vssd1 vccd1 vccd1 _19916_/D
+ sky130_fd_sc_hd__a211oi_4
XFILLER_133_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17705__S _18546_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16813__A0 _15768_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_207_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12800_ _12798_/Y _18829_/Q _12799_/Y _18815_/Q vssd1 vssd1 vccd1 vccd1 _12800_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_228_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13780_ _18732_/Q vssd1 vssd1 vccd1 vccd1 _13830_/A sky130_fd_sc_hd__inv_2
X_10992_ _10992_/A vssd1 vssd1 vccd1 vccd1 _10993_/B sky130_fd_sc_hd__inv_2
XFILLER_43_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12731_ _14816_/A vssd1 vssd1 vccd1 vccd1 _12731_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_42_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17440__S _17513_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15450_ _15450_/A _15450_/B vssd1 vssd1 vccd1 vccd1 _15450_/X sky130_fd_sc_hd__or2_1
XANTENNA__09059__B1 _09058_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12662_ _12698_/A vssd1 vssd1 vccd1 vccd1 _12699_/A sky130_fd_sc_hd__inv_2
XPHY_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14401_ _18397_/Q _14394_/X _14326_/X _14396_/X vssd1 vssd1 vccd1 vccd1 _18397_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11613_ _19561_/Q _11612_/Y _11588_/A _11575_/B vssd1 vssd1 vccd1 vccd1 _19561_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15381_ _18639_/Q _18637_/Q vssd1 vssd1 vccd1 vccd1 _17585_/S sky130_fd_sc_hd__nor2_1
XPHY_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11405__A2 _19128_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12593_ _19035_/Q _12590_/X _12356_/X _12591_/X vssd1 vssd1 vccd1 vccd1 _19035_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17120_ _17119_/X _15497_/Y _17513_/S vssd1 vssd1 vccd1 vccd1 _17120_/X sky130_fd_sc_hd__mux2_1
XPHY_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14332_ _18434_/Q _14319_/A _14314_/X _14320_/A vssd1 vssd1 vccd1 vccd1 _18434_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_7_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11544_ _19578_/Q _11617_/A _11504_/A _11541_/A vssd1 vssd1 vccd1 vccd1 _19578_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17051_ _17050_/X _11379_/Y _17548_/S vssd1 vssd1 vccd1 vccd1 _17051_/X sky130_fd_sc_hd__mux2_1
XFILLER_51_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14263_ _18471_/Q _14258_/X _12720_/X _14260_/X vssd1 vssd1 vccd1 vccd1 _18471_/D
+ sky130_fd_sc_hd__a22o_1
X_11475_ _11475_/A _11514_/A vssd1 vssd1 vccd1 vccd1 _11476_/B sky130_fd_sc_hd__or2_2
XFILLER_183_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16002_ _16238_/A vssd1 vssd1 vccd1 vccd1 _16002_/X sky130_fd_sc_hd__buf_2
XANTENNA__12366__B1 _12234_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13214_ _18888_/Q _13213_/Y _13214_/B1 _13176_/X vssd1 vssd1 vccd1 vccd1 _18888_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_143_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10426_ _19843_/Q _10417_/X _10425_/X _10419_/Y vssd1 vssd1 vccd1 vccd1 _19843_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__20088__RESET_B repeater204/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14194_ _19104_/Q vssd1 vssd1 vccd1 vccd1 _14194_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13145_ _19161_/Q vssd1 vssd1 vccd1 vccd1 _13145_/Y sky130_fd_sc_hd__inv_2
X_10357_ _10357_/A vssd1 vssd1 vccd1 vccd1 _10358_/B sky130_fd_sc_hd__inv_2
XFILLER_151_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12118__B1 _11909_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17953_ _18260_/CLK _17953_/D vssd1 vssd1 vccd1 vccd1 _17953_/Q sky130_fd_sc_hd__dfxtp_1
X_13076_ _13076_/A _13187_/A vssd1 vssd1 vccd1 vccd1 _13077_/B sky130_fd_sc_hd__or2_2
XFILLER_239_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10288_ _15716_/A _18643_/Q vssd1 vssd1 vccd1 vccd1 _17630_/S sky130_fd_sc_hd__or2_4
XANTENNA__17057__A0 _17473_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16904_ _16468_/Y _19270_/Q _17541_/S vssd1 vssd1 vccd1 vccd1 _16904_/X sky130_fd_sc_hd__mux2_1
X_12027_ _19346_/Q _12023_/X _12026_/X _12024_/X vssd1 vssd1 vccd1 vccd1 _19346_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_239_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17884_ _17880_/X _17881_/X _17882_/X _17883_/X _19633_/Q _19634_/Q vssd1 vssd1 vccd1
+ vccd1 _17884_/X sky130_fd_sc_hd__mux4_2
XFILLER_66_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16804__A0 _17486_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19623_ _19920_/CLK _19623_/D repeater229/X vssd1 vssd1 vccd1 vccd1 _19623_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_93_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16835_ _17486_/A0 _13092_/Y _17543_/S vssd1 vssd1 vccd1 vccd1 _16835_/X sky130_fd_sc_hd__mux2_1
XFILLER_54_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19554_ _19582_/CLK _19554_/D hold348/A vssd1 vssd1 vccd1 vccd1 _19554_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_65_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16766_ _15963_/X _12752_/Y _17534_/S vssd1 vssd1 vccd1 vccd1 _16766_/X sky130_fd_sc_hd__mux2_1
X_13978_ _18696_/Q vssd1 vssd1 vccd1 vccd1 _14026_/A sky130_fd_sc_hd__inv_2
XANTENNA__09298__B1 _09105_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14291__B1 _14273_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18505_ _19812_/CLK _18505_/D repeater222/X vssd1 vssd1 vccd1 vccd1 _18505_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_62_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15717_ _19876_/Q vssd1 vssd1 vccd1 vccd1 _15717_/Y sky130_fd_sc_hd__inv_2
X_12929_ _19290_/Q vssd1 vssd1 vccd1 vccd1 _12929_/Y sky130_fd_sc_hd__inv_2
X_16697_ _17002_/X _16687_/X _17008_/X _16688_/X _16696_/X vssd1 vssd1 vccd1 vccd1
+ _16698_/C sky130_fd_sc_hd__o221a_1
X_19485_ _19510_/CLK hold158/X repeater260/X vssd1 vssd1 vccd1 vccd1 _19485_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__16568__C1 _16567_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17350__S _17518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19953__RESET_B repeater245/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10852__B1 _10425_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18436_ _18795_/CLK _18436_/D vssd1 vssd1 vccd1 vccd1 _18436_/Q sky130_fd_sc_hd__dfxtp_1
X_15648_ _18606_/Q vssd1 vssd1 vccd1 vccd1 _15648_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16474__B _17473_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_221_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18367_ _19637_/CLK _18367_/D vssd1 vssd1 vccd1 vccd1 _18367_/Q sky130_fd_sc_hd__dfxtp_1
X_15579_ _18589_/Q vssd1 vssd1 vccd1 vccd1 _15581_/A sky130_fd_sc_hd__inv_2
XFILLER_14_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17318_ _17317_/X _15602_/A _17318_/S vssd1 vssd1 vccd1 vccd1 _17318_/X sky130_fd_sc_hd__mux2_1
XFILLER_119_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18298_ _18431_/CLK _18298_/D vssd1 vssd1 vccd1 vccd1 _18298_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17249_ _16585_/Y _19279_/Q _17541_/S vssd1 vssd1 vccd1 vccd1 _17249_/X sky130_fd_sc_hd__mux2_1
XANTENNA__16740__C1 _16739_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12357__B1 _12356_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13619__A _18757_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12523__A hold268/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12109__B1 _12107_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18835__RESET_B repeater239/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08953_ _19860_/Q vssd1 vssd1 vccd1 vccd1 _10361_/A sky130_fd_sc_hd__inv_2
XANTENNA__17048__A0 _17047_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17525__S _17537_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16649__B _16668_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09289__B1 _09079_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14282__B1 _13676_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_225_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09505_ _19323_/Q vssd1 vssd1 vccd1 vccd1 _16720_/A sky130_fd_sc_hd__inv_2
XFILLER_213_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16559__C1 _16558_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_225_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19694__RESET_B repeater208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17260__S _17548_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09436_ _19382_/Q vssd1 vssd1 vccd1 vccd1 _09436_/Y sky130_fd_sc_hd__inv_2
XFILLER_169_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09367_ _20010_/Q vssd1 vssd1 vccd1 vccd1 _09471_/A sky130_fd_sc_hd__inv_2
X_09298_ _20041_/Q _09293_/X _09105_/X _09294_/X vssd1 vssd1 vccd1 vccd1 _20041_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_165_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11260_ _19609_/Q _11258_/Y _11476_/A _19010_/Q vssd1 vssd1 vccd1 vccd1 _11260_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10211_ _10956_/B vssd1 vssd1 vccd1 vccd1 _10211_/X sky130_fd_sc_hd__buf_1
XANTENNA__13529__A _13529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20110__RESET_B repeater217/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11191_ _11191_/A vssd1 vssd1 vccd1 vccd1 _11191_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__17992__CLK _18169_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18576__RESET_B repeater269/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10142_ _16983_/X _10136_/X _19900_/Q _10138_/X vssd1 vssd1 vccd1 vccd1 _19900_/D
+ sky130_fd_sc_hd__o22a_1
XANTENNA__17039__A0 _15768_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13848__B1 _13845_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17435__S _17565_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18505__RESET_B repeater222/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10073_ _10038_/A _10038_/B _10079_/A _10071_/Y vssd1 vssd1 vccd1 vccd1 _19922_/D
+ sky130_fd_sc_hd__a211oi_2
X_14950_ _18082_/Q _14940_/A _14949_/X _14941_/A vssd1 vssd1 vccd1 vccd1 _18082_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_87_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13901_ _13925_/A vssd1 vssd1 vccd1 vccd1 _13901_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_101_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14881_ _18122_/Q _14872_/A _14868_/X _14873_/A vssd1 vssd1 vccd1 vccd1 _18122_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_248_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16620_ _16620_/A _16621_/B vssd1 vssd1 vccd1 vccd1 _16620_/Y sky130_fd_sc_hd__nor2_1
XFILLER_47_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13832_ _13832_/A _13832_/B vssd1 vssd1 vccd1 vccd1 _13833_/A sky130_fd_sc_hd__or2_1
XFILLER_28_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_150_HCLK clkbuf_4_1_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19859_/CLK sky130_fd_sc_hd__clkbuf_16
X_16551_ _19039_/Q _16622_/B vssd1 vssd1 vccd1 vccd1 _16551_/Y sky130_fd_sc_hd__nand2_1
XFILLER_46_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13763_ _18745_/Q _13753_/B _13753_/Y _13760_/X vssd1 vssd1 vccd1 vccd1 _13763_/X
+ sky130_fd_sc_hd__o211a_1
X_10975_ _10975_/A vssd1 vssd1 vccd1 vccd1 _10976_/B sky130_fd_sc_hd__inv_2
XFILLER_189_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17170__S _17534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15502_ _18570_/Q _15498_/A _15501_/Y _15498_/Y vssd1 vssd1 vccd1 vccd1 _15503_/B
+ sky130_fd_sc_hd__o22a_1
X_12714_ _14802_/A vssd1 vssd1 vccd1 vccd1 _12714_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_188_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16482_ _15199_/A _16475_/X _16492_/A _16476_/X _16481_/X vssd1 vssd1 vccd1 vccd1
+ _16482_/Y sky130_fd_sc_hd__o221ai_4
X_19270_ _19282_/CLK _19270_/D repeater216/X vssd1 vssd1 vccd1 vccd1 _19270_/Q sky130_fd_sc_hd__dfrtp_1
X_13694_ _12313_/X _10345_/X _13694_/S vssd1 vssd1 vccd1 vccd1 _18766_/D sky130_fd_sc_hd__mux2_1
XANTENNA__17762__A1 _13491_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19743__CLK _20070_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15433_ _19624_/Q _11169_/B _11170_/B vssd1 vssd1 vccd1 vccd1 _15433_/X sky130_fd_sc_hd__a21bo_1
X_18221_ _20076_/CLK _18221_/D vssd1 vssd1 vccd1 vccd1 _18221_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12645_ _19003_/Q _12643_/X hold239/X _12644_/X vssd1 vssd1 vccd1 vccd1 _19003_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_repeater167_A _17522_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12587__B1 hold281/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15364_ _15364_/A _17587_/X vssd1 vssd1 vccd1 vccd1 _18503_/D sky130_fd_sc_hd__and2_1
XFILLER_30_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18152_ _18169_/CLK _18152_/D vssd1 vssd1 vccd1 vccd1 _18152_/Q sky130_fd_sc_hd__dfxtp_1
X_12576_ _12576_/A vssd1 vssd1 vccd1 vccd1 _12576_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__12051__A2 _12016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17514__A1 _15479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14315_ _18442_/Q _14304_/A _14314_/X _14305_/A vssd1 vssd1 vccd1 vccd1 _18442_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17103_ _17102_/X _19134_/Q _17548_/S vssd1 vssd1 vccd1 vccd1 _17103_/X sky130_fd_sc_hd__mux2_1
X_11527_ _11468_/B _11527_/A2 _11468_/A vssd1 vssd1 vccd1 vccd1 _11528_/C sky130_fd_sc_hd__o21a_1
XPHY_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18083_ _18260_/CLK _18083_/D vssd1 vssd1 vccd1 vccd1 _18083_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14245__D _14245_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15295_ _15318_/A _15295_/B vssd1 vssd1 vccd1 vccd1 _17755_/S sky130_fd_sc_hd__nor2_2
XFILLER_183_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12339__B1 _12102_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17034_ _17033_/X _12894_/Y _17487_/S vssd1 vssd1 vccd1 vccd1 _17034_/X sky130_fd_sc_hd__mux2_1
XFILLER_183_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output96_A _16691_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold309 HWDATA[25] vssd1 vssd1 vccd1 vccd1 input55/A sky130_fd_sc_hd__dlygate4sd3_1
X_14246_ _11926_/A _18663_/Q _14246_/S vssd1 vssd1 vccd1 vccd1 _18663_/D sky130_fd_sc_hd__mux2_1
X_11458_ _11566_/B vssd1 vssd1 vccd1 vccd1 _11592_/A sky130_fd_sc_hd__inv_2
XFILLER_7_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17278__A0 _17473_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10409_ _10409_/A vssd1 vssd1 vccd1 vccd1 _14681_/A sky130_fd_sc_hd__buf_1
X_14177_ _19095_/Q vssd1 vssd1 vccd1 vccd1 _14177_/Y sky130_fd_sc_hd__inv_2
X_11389_ _11389_/A _11389_/B _11389_/C _11389_/D vssd1 vssd1 vccd1 vccd1 _11457_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_113_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13128_ _19173_/Q vssd1 vssd1 vccd1 vccd1 _13128_/Y sky130_fd_sc_hd__inv_2
X_18985_ _19608_/CLK _18985_/D hold273/X vssd1 vssd1 vccd1 vccd1 _18985_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__17345__S _17566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17936_ _19545_/CLK _17936_/D vssd1 vssd1 vccd1 vccd1 _17936_/Q sky130_fd_sc_hd__dfxtp_1
X_13059_ _18887_/Q vssd1 vssd1 vccd1 vccd1 _13060_/A sky130_fd_sc_hd__inv_2
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_239_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16469__B _16469_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12511__B1 _12410_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_239_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater148 _17486_/A0 vssd1 vssd1 vccd1 vccd1 _17473_/A0 sky130_fd_sc_hd__clkbuf_16
X_17867_ _16185_/Y _16186_/Y _16187_/Y _16188_/Y _17908_/S0 _18759_/Q vssd1 vssd1
+ vccd1 vccd1 _17867_/X sky130_fd_sc_hd__mux4_1
XFILLER_38_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrepeater159 _17490_/S vssd1 vssd1 vccd1 vccd1 _17544_/S sky130_fd_sc_hd__buf_8
XFILLER_226_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19606_ _19609_/CLK _19606_/D hold359/X vssd1 vssd1 vccd1 vccd1 _19606_/Q sky130_fd_sc_hd__dfrtp_1
X_16818_ _16817_/X _13545_/A _17536_/S vssd1 vssd1 vccd1 vccd1 _16818_/X sky130_fd_sc_hd__mux2_1
XFILLER_242_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17798_ _18296_/Q _18288_/Q _18280_/Q _18448_/Q _17923_/S0 _19646_/Q vssd1 vssd1
+ vccd1 vccd1 _17798_/X sky130_fd_sc_hd__mux4_2
XFILLER_54_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19537_ _19540_/CLK _19537_/D repeater220/X vssd1 vssd1 vccd1 vccd1 _19537_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__12814__A1 _19231_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16749_ _16201_/Y _16294_/Y _16113_/Y _16200_/X _16748_/X vssd1 vssd1 vccd1 vccd1
+ _16750_/B sky130_fd_sc_hd__o221a_2
XFILLER_235_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17080__S _17517_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19468_ _19470_/CLK _19468_/D repeater274/X vssd1 vssd1 vccd1 vccd1 _19468_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17753__A1 _11153_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09221_ _18650_/Q _09214_/B _09220_/Y _18651_/Q _09214_/Y vssd1 vssd1 vccd1 vccd1
+ _18651_/D sky130_fd_sc_hd__a32o_1
X_18419_ _18435_/CLK _18419_/D vssd1 vssd1 vccd1 vccd1 _18419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19399_ _19997_/CLK _19399_/D repeater271/X vssd1 vssd1 vccd1 vccd1 _19399_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__19034__RESET_B repeater267/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12578__B1 _12401_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09152_ _15322_/A _15322_/C _09156_/B _09125_/D _09151_/Y vssd1 vssd1 vccd1 vccd1
+ _09153_/A sky130_fd_sc_hd__o32a_1
XFILLER_147_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_238_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09083_ _20098_/Q _09069_/X _09082_/X _09072_/X vssd1 vssd1 vccd1 vccd1 _20098_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_190_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_190_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput70 input70/A vssd1 vssd1 vccd1 vccd1 input70/X sky130_fd_sc_hd__buf_2
XFILLER_128_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_31_HCLK _18641_/CLK vssd1 vssd1 vccd1 vccd1 _20090_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_162_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09985_ _19950_/Q _09987_/A _09968_/X _09985_/C1 vssd1 vssd1 vccd1 vccd1 _19950_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_130_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17255__S _17547_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15564__A _15571_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08936_ _19857_/Q vssd1 vssd1 vccd1 vccd1 _10323_/A sky130_fd_sc_hd__inv_2
XFILLER_88_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12502__B1 _12394_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17441__A0 _17486_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18640__CLK _19780_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19804__RESET_B repeater222/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10760_ _10765_/B _19750_/Q vssd1 vssd1 vccd1 vccd1 _10761_/A sky130_fd_sc_hd__or2b_1
XFILLER_16_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09419_ _19931_/Q vssd1 vssd1 vccd1 vccd1 _10047_/A sky130_fd_sc_hd__inv_2
XFILLER_240_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10691_ _12257_/A _15858_/D vssd1 vssd1 vccd1 vccd1 _10718_/A sky130_fd_sc_hd__or2_2
XFILLER_200_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11332__A _18981_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12430_ _19131_/Q _12427_/X _12302_/X _12428_/X vssd1 vssd1 vccd1 vccd1 _19131_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_200_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12361_ _12361_/A vssd1 vssd1 vccd1 vccd1 _12361_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_181_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14100_ _14032_/A _14100_/A2 _14033_/Y _14135_/B vssd1 vssd1 vccd1 vccd1 _18702_/D
+ sky130_fd_sc_hd__a211oi_2
X_11312_ _18967_/Q vssd1 vssd1 vccd1 vccd1 _11312_/Y sky130_fd_sc_hd__inv_2
XFILLER_165_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15080_ _18003_/Q _15072_/A _14780_/X _15073_/A vssd1 vssd1 vccd1 vccd1 _18003_/D
+ sky130_fd_sc_hd__a22o_1
X_12292_ _19204_/Q _12290_/X _12035_/X _12291_/X vssd1 vssd1 vccd1 vccd1 _19204_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_5_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14031_ _14031_/A _14031_/B vssd1 vssd1 vccd1 vccd1 _14032_/B sky130_fd_sc_hd__or2_2
X_11243_ _19595_/Q vssd1 vssd1 vccd1 vccd1 _11475_/A sky130_fd_sc_hd__inv_2
XANTENNA__20123__CLK _20123_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11174_ _19626_/Q _11170_/X _18879_/Q _11173_/X vssd1 vssd1 vccd1 vccd1 _18546_/D
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__19296__CLK _20013_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17165__S _17535_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10125_ _15509_/B _10125_/B vssd1 vssd1 vccd1 vccd1 _15547_/B sky130_fd_sc_hd__or2_1
X_18770_ _20058_/CLK _18770_/D repeater271/X vssd1 vssd1 vccd1 vccd1 _18770_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_95_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15982_ _10707_/Y _15854_/X _15981_/Y _15867_/B vssd1 vssd1 vccd1 vccd1 _15982_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__15691__C1 _15643_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17721_ _19679_/Q _19692_/Q _18510_/Q vssd1 vssd1 vccd1 vccd1 _17721_/X sky130_fd_sc_hd__mux2_1
XFILLER_76_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10056_ _19933_/Q _10055_/Y _10009_/B _10055_/A _10053_/X vssd1 vssd1 vccd1 vccd1
+ _19933_/D sky130_fd_sc_hd__o221a_1
X_14933_ _20076_/Q vssd1 vssd1 vccd1 vccd1 _14933_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_102_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output134_A _15731_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17652_ _15627_/Y _19037_/Q _17655_/S vssd1 vssd1 vccd1 vccd1 _18600_/D sky130_fd_sc_hd__mux2_1
XFILLER_224_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10411__A _10842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14864_ _18134_/Q _14858_/X _14707_/X _14860_/X vssd1 vssd1 vccd1 vccd1 _18134_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_208_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19545__RESET_B repeater221/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16603_ _16818_/X _16394_/X _16878_/X _15898_/X vssd1 vssd1 vccd1 vccd1 _16603_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_35_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13815_ _13909_/D _13815_/B vssd1 vssd1 vccd1 vccd1 _13941_/A sky130_fd_sc_hd__or2_1
XFILLER_90_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17583_ _15392_/X _19524_/Q _17584_/S vssd1 vssd1 vccd1 vccd1 _17583_/X sky130_fd_sc_hd__mux2_1
X_14795_ hold264/X vssd1 vssd1 vccd1 vccd1 hold263/A sky130_fd_sc_hd__buf_2
XFILLER_217_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19322_ _19324_/CLK _19322_/D repeater213/X vssd1 vssd1 vccd1 vccd1 _19322_/Q sky130_fd_sc_hd__dfrtp_4
X_16534_ _19452_/Q vssd1 vssd1 vccd1 vccd1 _16534_/Y sky130_fd_sc_hd__inv_2
X_13746_ _13746_/A _15192_/B vssd1 vssd1 vccd1 vccd1 _15191_/A sky130_fd_sc_hd__or2_1
X_10958_ _10958_/A _11005_/A vssd1 vssd1 vccd1 vccd1 _11001_/A sky130_fd_sc_hd__or2_1
XFILLER_189_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19253_ _19324_/CLK _19253_/D repeater237/X vssd1 vssd1 vccd1 vccd1 _19253_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_189_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16465_ _15846_/A _16448_/X _15859_/A _16457_/X _16464_/X vssd1 vssd1 vccd1 vccd1
+ _16465_/Y sky130_fd_sc_hd__o221ai_4
X_13677_ _18775_/Q _13671_/X _13676_/X _13672_/X vssd1 vssd1 vccd1 vccd1 _18775_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_189_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10889_ _19695_/Q _10878_/A _10866_/X _10879_/A vssd1 vssd1 vccd1 vccd1 _19695_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_31_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17830__S1 _18750_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18204_ _18460_/CLK _18204_/D vssd1 vssd1 vccd1 vccd1 _18204_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15416_ _18540_/Q _13227_/B _13228_/B vssd1 vssd1 vccd1 vccd1 _15416_/X sky130_fd_sc_hd__a21bo_1
X_12628_ _19014_/Q _12622_/X _12398_/X _12623_/X vssd1 vssd1 vccd1 vccd1 _19014_/D
+ sky130_fd_sc_hd__a22o_1
X_19184_ _19293_/CLK _19184_/D repeater187/X vssd1 vssd1 vccd1 vccd1 _19184_/Q sky130_fd_sc_hd__dfrtp_1
X_16396_ _11742_/A _16389_/X _16391_/X _16393_/X _16395_/X vssd1 vssd1 vccd1 vccd1
+ _16396_/X sky130_fd_sc_hd__o2111a_1
XPHY_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_54_HCLK clkbuf_opt_2_HCLK/A vssd1 vssd1 vccd1 vccd1 _19772_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__16752__B _19741_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15347_ _15347_/A _17595_/X vssd1 vssd1 vccd1 vccd1 _18495_/D sky130_fd_sc_hd__and2_1
X_18135_ _20124_/CLK _18135_/D vssd1 vssd1 vccd1 vccd1 _18135_/Q sky130_fd_sc_hd__dfxtp_1
X_12559_ _12598_/A vssd1 vssd1 vccd1 vccd1 _12576_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_129_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18498__RESET_B repeater203/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15278_ _19724_/Q _15278_/B _18513_/Q _18479_/D vssd1 vssd1 vccd1 vccd1 _15278_/X
+ sky130_fd_sc_hd__or4_4
X_18066_ _19851_/CLK _18066_/D vssd1 vssd1 vccd1 vccd1 _18066_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__18513__CLK _19780_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold128 hold352/X vssd1 vssd1 vccd1 vccd1 hold351/A sky130_fd_sc_hd__dlygate4sd3_1
X_14229_ _18499_/Q _14229_/B vssd1 vssd1 vccd1 vccd1 _14230_/B sky130_fd_sc_hd__or2_1
Xhold139 input16/X vssd1 vssd1 vccd1 vccd1 hold139/X sky130_fd_sc_hd__dlygate4sd3_1
X_17017_ _17016_/X _13886_/Y _17545_/S vssd1 vssd1 vccd1 vccd1 _17017_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17897__S1 _18759_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_159_HCLK_A clkbuf_4_0_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17075__S _17493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09770_ _19995_/Q _09769_/Y _09763_/X _09752_/B vssd1 vssd1 vccd1 vccd1 _19995_/D
+ sky130_fd_sc_hd__o211a_1
X_18968_ _19208_/CLK _18968_/D hold363/X vssd1 vssd1 vccd1 vccd1 _18968_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_86_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17919_ _17915_/X _17916_/X _17917_/X _17918_/X _18751_/Q _18752_/Q vssd1 vssd1 vccd1
+ vccd1 _17919_/X sky130_fd_sc_hd__mux4_2
XFILLER_67_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18899_ _19352_/CLK _18899_/D repeater188/X vssd1 vssd1 vccd1 vccd1 _18899_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__09813__C _09813_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_242_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_179_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17821__S1 _18750_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09204_ _08977_/C _09203_/X _09200_/X vssd1 vssd1 vccd1 vccd1 _20069_/D sky130_fd_sc_hd__a21oi_1
XFILLER_210_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09135_ _13494_/A vssd1 vssd1 vccd1 vccd1 _15322_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__11774__A1 hold206/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18850__RESET_B repeater232/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09066_ hold271/X vssd1 vssd1 vccd1 vccd1 _12032_/A sky130_fd_sc_hd__buf_4
XFILLER_163_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17888__S1 _18759_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16465__A1 _15846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09968_ _09968_/A vssd1 vssd1 vccd1 vccd1 _09968_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_134_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_18_HCLK_A clkbuf_4_3_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08919_ _08919_/A vssd1 vssd1 vccd1 vccd1 _09198_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_246_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20088_ _20089_/CLK _20088_/D repeater204/X vssd1 vssd1 vccd1 vccd1 _20088_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_100_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11829__A2 _11800_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09899_ _19941_/Q _09896_/Y _09850_/A _19333_/Q _09898_/X vssd1 vssd1 vccd1 vccd1
+ _09899_/X sky130_fd_sc_hd__a221o_1
XFILLER_18_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17713__S _18546_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11930_ _19399_/Q vssd1 vssd1 vccd1 vccd1 _15512_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_58_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_6_HCLK_A clkbuf_4_2_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11861_ _13630_/A _11861_/B _17610_/X _17614_/X vssd1 vssd1 vccd1 vccd1 _11862_/A
+ sky130_fd_sc_hd__or4b_4
XFILLER_150_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13600_ _13536_/A _13600_/A2 _13588_/X _13598_/Y vssd1 vssd1 vccd1 vccd1 _18812_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_60_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10812_ _17616_/X _10808_/X _19731_/Q _10810_/X vssd1 vssd1 vccd1 vccd1 _19731_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_72_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14580_ _14793_/A vssd1 vssd1 vccd1 vccd1 _14580_/X sky130_fd_sc_hd__clkbuf_2
XPHY_3943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11792_ _19466_/Q _11784_/X _09027_/X _11787_/X vssd1 vssd1 vccd1 vccd1 _19466_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_77_HCLK clkbuf_opt_4_HCLK/A vssd1 vssd1 vccd1 vccd1 _19255_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_3965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13531_ _13531_/A _13607_/A vssd1 vssd1 vccd1 vccd1 _13532_/B sky130_fd_sc_hd__or2_2
XPHY_3976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10743_ _10743_/A vssd1 vssd1 vccd1 vccd1 _10743_/X sky130_fd_sc_hd__buf_1
XPHY_3987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17812__S1 _18750_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11062__A _19632_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16250_ _17379_/X _16235_/X _16237_/Y _16242_/X _16249_/X vssd1 vssd1 vccd1 vccd1
+ _16250_/X sky130_fd_sc_hd__o2111a_2
X_13462_ _13462_/A vssd1 vssd1 vccd1 vccd1 _13483_/A sky130_fd_sc_hd__buf_2
XFILLER_174_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10674_ _17737_/X _10669_/X _19788_/Q _10670_/X vssd1 vssd1 vccd1 vccd1 _19788_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_41_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14400__B1 hold324/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15201_ _15233_/A _15201_/B vssd1 vssd1 vccd1 vccd1 _15201_/X sky130_fd_sc_hd__or2_1
X_12413_ hold277/X vssd1 vssd1 vccd1 vccd1 _12413_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__11997__A _12187_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16181_ _18270_/Q vssd1 vssd1 vccd1 vccd1 _16181_/Y sky130_fd_sc_hd__inv_2
X_13393_ _13390_/Y _18857_/Q _13391_/Y _18863_/Q _13392_/X vssd1 vssd1 vccd1 vccd1
+ _13402_/B sky130_fd_sc_hd__o221a_1
XFILLER_154_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15132_ _17969_/Q _15123_/A _14949_/X _15124_/A vssd1 vssd1 vccd1 vccd1 _17969_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_182_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12344_ hold234/X vssd1 vssd1 vccd1 vccd1 _12344_/X sky130_fd_sc_hd__buf_4
XANTENNA__18591__RESET_B repeater269/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16999__S _17386_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15063_ _18016_/Q _15059_/X _14806_/A _15061_/X vssd1 vssd1 vccd1 vccd1 _18016_/D
+ sky130_fd_sc_hd__a22o_1
X_19940_ _19976_/CLK _19940_/D hold371/X vssd1 vssd1 vccd1 vccd1 _19940_/Q sky130_fd_sc_hd__dfrtp_1
X_12275_ _19215_/Q _12269_/X _12092_/X _12270_/X vssd1 vssd1 vccd1 vccd1 _19215_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_135_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14014_ _14014_/A _14014_/B vssd1 vssd1 vccd1 vccd1 _14129_/A sky130_fd_sc_hd__or2_1
XFILLER_141_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11226_ _19584_/Q vssd1 vssd1 vccd1 vccd1 _11465_/A sky130_fd_sc_hd__inv_2
XANTENNA__09186__A2 _09164_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19871_ _20070_/CLK _19871_/D repeater207/X vssd1 vssd1 vccd1 vccd1 _19871_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17879__S1 _18761_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18822_ _18827_/CLK _18822_/D repeater217/X vssd1 vssd1 vccd1 vccd1 _18822_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_110_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11157_ _19612_/Q _19611_/Q vssd1 vssd1 vccd1 vccd1 _11158_/B sky130_fd_sc_hd__or2_1
XFILLER_150_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14467__B1 _14441_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10108_ _10101_/A _10101_/B _19906_/Q _10030_/A _10053_/X vssd1 vssd1 vccd1 vccd1
+ _19906_/D sky130_fd_sc_hd__o221a_1
XFILLER_95_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19726__RESET_B repeater207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18753_ _18869_/CLK _18753_/D repeater195/X vssd1 vssd1 vccd1 vccd1 _18753_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_49_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11088_ _19639_/Q _12545_/A _12053_/B vssd1 vssd1 vccd1 vccd1 _14255_/A sky130_fd_sc_hd__or3_1
X_15965_ _19440_/Q vssd1 vssd1 vccd1 vccd1 _15965_/Y sky130_fd_sc_hd__inv_2
XFILLER_191_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17405__A0 _17473_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17704_ _17985_/Q _19756_/Q _18548_/Q vssd1 vssd1 vccd1 vccd1 _17704_/X sky130_fd_sc_hd__mux2_1
X_10039_ _10039_/A _10071_/A vssd1 vssd1 vccd1 vccd1 _10040_/B sky130_fd_sc_hd__or2_2
X_14916_ _18100_/Q _14909_/A _14711_/X _14910_/A vssd1 vssd1 vccd1 vccd1 _18100_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_208_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18684_ _18686_/CLK _18684_/D repeater252/X vssd1 vssd1 vccd1 vccd1 _18684_/Q sky130_fd_sc_hd__dfrtp_1
X_15896_ _16530_/A vssd1 vssd1 vccd1 vccd1 _15896_/X sky130_fd_sc_hd__buf_2
XFILLER_63_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17635_ _15699_/X _19054_/Q _17664_/S vssd1 vssd1 vccd1 vccd1 _18617_/D sky130_fd_sc_hd__mux2_1
X_14847_ _14847_/A vssd1 vssd1 vccd1 vccd1 _14847_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_224_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18066__CLK _19851_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17566_ _17565_/X _10212_/Y _17566_/S vssd1 vssd1 vccd1 vccd1 _17566_/X sky130_fd_sc_hd__mux2_1
X_14778_ _18181_/Q _14771_/X _14725_/X _14773_/X vssd1 vssd1 vccd1 vccd1 _18181_/D
+ sky130_fd_sc_hd__a22o_1
X_19305_ _20035_/CLK _19305_/D repeater242/X vssd1 vssd1 vccd1 vccd1 _19305_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_16_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16517_ _19450_/Q vssd1 vssd1 vccd1 vccd1 _16517_/Y sky130_fd_sc_hd__inv_2
XFILLER_232_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13729_ _13729_/A vssd1 vssd1 vccd1 vccd1 _14975_/B sky130_fd_sc_hd__buf_1
XFILLER_204_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17803__S1 _18750_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17497_ _15960_/X _19879_/Q _19498_/Q vssd1 vssd1 vccd1 vccd1 _17497_/X sky130_fd_sc_hd__mux2_1
XFILLER_176_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19236_ _19282_/CLK _19236_/D repeater215/X vssd1 vssd1 vccd1 vccd1 _19236_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__18679__RESET_B repeater252/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16448_ _15205_/Y _15840_/X _16442_/X _16447_/X vssd1 vssd1 vccd1 vccd1 _16448_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_158_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16392__B1 _17341_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19167_ _19214_/CLK _19167_/D hold367/X vssd1 vssd1 vccd1 vccd1 _19167_/Q sky130_fd_sc_hd__dfrtp_4
X_16379_ _16371_/Y _15867_/B _16374_/X _16378_/X vssd1 vssd1 vccd1 vccd1 _16379_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_144_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18118_ _18142_/CLK _18118_/D vssd1 vssd1 vccd1 vccd1 _18118_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19098_ _19585_/CLK _19098_/D repeater252/X vssd1 vssd1 vccd1 vccd1 _19098_/Q sky130_fd_sc_hd__dfrtp_4
X_18049_ _18959_/CLK _18049_/D vssd1 vssd1 vccd1 vccd1 _18049_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12705__B1 _12541_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20011_ _20013_/CLK _20011_/D repeater240/X vssd1 vssd1 vccd1 vccd1 _20011_/Q sky130_fd_sc_hd__dfrtp_1
X_09822_ _19964_/Q vssd1 vssd1 vccd1 vccd1 _09872_/A sky130_fd_sc_hd__inv_2
XFILLER_101_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14458__B1 _14417_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16003__A _16633_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19467__RESET_B repeater274/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09753_ _09753_/A _09765_/A _09753_/C vssd1 vssd1 vccd1 vccd1 _09761_/A sky130_fd_sc_hd__or3_4
XFILLER_101_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17533__S _17539_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15842__A _16055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09684_ _19427_/Q vssd1 vssd1 vccd1 vccd1 _09684_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_199_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18559__CLK _19992_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16383__B1 _16382_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_6_HCLK clkbuf_4_2_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _18954_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_183_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09118_ _20087_/Q vssd1 vssd1 vccd1 vccd1 _13494_/A sky130_fd_sc_hd__inv_2
XFILLER_182_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10390_ _19850_/Q vssd1 vssd1 vccd1 vccd1 _14477_/B sky130_fd_sc_hd__buf_1
XFILLER_135_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17708__S _18546_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09049_ hold310/X vssd1 vssd1 vccd1 vccd1 _09049_/X sky130_fd_sc_hd__buf_4
XANTENNA__10226__A _19836_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10970__A2 _17614_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12060_ _15881_/B _12066_/A vssd1 vssd1 vccd1 vccd1 _12061_/S sky130_fd_sc_hd__or2_1
XFILLER_104_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11011_ _11006_/B _11010_/Y _10978_/X _10989_/A _10957_/A vssd1 vssd1 vccd1 vccd1
+ _11012_/A sky130_fd_sc_hd__o32a_1
XANTENNA__12441__A _12457_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14449__B1 _14405_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_142_HCLK_A clkbuf_4_3_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17443__S _17543_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15750_ _18663_/Q _18476_/Q vssd1 vssd1 vccd1 vccd1 _15750_/X sky130_fd_sc_hd__and2_2
X_12962_ _13060_/B vssd1 vssd1 vccd1 vccd1 _12962_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_246_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14701_ _14701_/A vssd1 vssd1 vccd1 vccd1 _14701_/X sky130_fd_sc_hd__clkbuf_2
X_11913_ _19408_/Q _11905_/X _10877_/X _11906_/X vssd1 vssd1 vccd1 vccd1 _19408_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_246_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15681_ _18613_/Q _15681_/B vssd1 vssd1 vccd1 vccd1 _15686_/B sky130_fd_sc_hd__or2_1
XFILLER_18_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12893_ _18950_/Q vssd1 vssd1 vccd1 vccd1 _12893_/Y sky130_fd_sc_hd__inv_2
XPHY_4430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14368__A _14368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17420_ _17419_/X _13063_/A _17488_/S vssd1 vssd1 vccd1 vccd1 _17420_/X sky130_fd_sc_hd__mux2_1
XPHY_4463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16610__B2 _15898_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11844_ _15867_/A _16055_/A vssd1 vssd1 vccd1 vccd1 _12372_/A sky130_fd_sc_hd__or2_4
X_14632_ _14632_/A vssd1 vssd1 vccd1 vccd1 _14632_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_221_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14563_ _18303_/Q _14558_/X _14537_/X _14560_/X vssd1 vssd1 vccd1 vccd1 _18303_/D
+ sky130_fd_sc_hd__a22o_1
X_17351_ _17486_/A0 _09891_/Y _17543_/S vssd1 vssd1 vccd1 vccd1 _17351_/X sky130_fd_sc_hd__mux2_1
XPHY_3773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11775_ hold199/X _11771_/X _19473_/Q _11772_/X vssd1 vssd1 vccd1 vccd1 hold201/A
+ sky130_fd_sc_hd__o22a_1
XPHY_3784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17797__S0 _17923_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16302_ _19706_/Q vssd1 vssd1 vccd1 vccd1 _16302_/Y sky130_fd_sc_hd__inv_2
X_10726_ _19769_/Q _10720_/X _10418_/X _10722_/X vssd1 vssd1 vccd1 vccd1 _19769_/D
+ sky130_fd_sc_hd__a22o_1
X_13514_ _18763_/Q _14628_/B _13506_/A vssd1 vssd1 vccd1 vccd1 _13516_/A sky130_fd_sc_hd__o21ai_1
XFILLER_202_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16374__B1 _16373_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17282_ _17281_/X _13537_/A _17386_/S vssd1 vssd1 vccd1 vccd1 _17282_/X sky130_fd_sc_hd__mux2_2
X_14494_ _18345_/Q _14491_/X _12714_/X _14493_/X vssd1 vssd1 vccd1 vccd1 _18345_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_146_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19021_ _19609_/CLK _19021_/D hold357/X vssd1 vssd1 vccd1 vccd1 _19021_/Q sky130_fd_sc_hd__dfrtp_2
X_13445_ _13445_/A vssd1 vssd1 vccd1 vccd1 _13445_/X sky130_fd_sc_hd__buf_2
X_16233_ _15253_/Y _15840_/X _16226_/Y _15836_/X _16232_/X vssd1 vssd1 vccd1 vccd1
+ _16233_/X sky130_fd_sc_hd__o221a_1
XANTENNA__18701__RESET_B hold351/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15199__A _15199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10657_ _18488_/Q vssd1 vssd1 vccd1 vccd1 _10658_/C sky130_fd_sc_hd__inv_2
XFILLER_9_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12935__B1 _12933_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13376_ _13373_/Y _18855_/Q _20109_/Q _13429_/A _13375_/X vssd1 vssd1 vccd1 vccd1
+ _13376_/X sky130_fd_sc_hd__a221o_1
XFILLER_166_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16164_ _18342_/Q vssd1 vssd1 vccd1 vccd1 _16164_/Y sky130_fd_sc_hd__inv_2
X_10588_ _10589_/C _10589_/B _19798_/Q vssd1 vssd1 vccd1 vccd1 _10614_/B sky130_fd_sc_hd__and3b_1
XFILLER_182_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17874__A0 _17870_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19978__RESET_B repeater192/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12327_ _12334_/A vssd1 vssd1 vccd1 vccd1 _12327_/X sky130_fd_sc_hd__buf_1
X_15115_ _17982_/Q _15110_/X _14927_/X _15112_/X vssd1 vssd1 vccd1 vccd1 _17982_/D
+ sky130_fd_sc_hd__a22o_1
X_16095_ _18229_/Q vssd1 vssd1 vccd1 vccd1 _16095_/Y sky130_fd_sc_hd__inv_2
X_19923_ _19927_/CLK _19923_/D repeater230/X vssd1 vssd1 vccd1 vccd1 _19923_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__19907__RESET_B repeater241/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15046_ _15094_/A _19850_/Q _15058_/C vssd1 vssd1 vccd1 vccd1 _15048_/A sky130_fd_sc_hd__or3_4
X_12258_ _12372_/A _12487_/B vssd1 vssd1 vccd1 vccd1 _12298_/A sky130_fd_sc_hd__or2_2
XFILLER_141_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11209_ _11460_/A _18993_/Q _19606_/Q _11208_/Y vssd1 vssd1 vccd1 vccd1 _11209_/X
+ sky130_fd_sc_hd__o22a_1
X_19854_ _19855_/CLK _19854_/D repeater265/X vssd1 vssd1 vccd1 vccd1 _19854_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_69_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12189_ _12205_/A vssd1 vssd1 vccd1 vccd1 _12189_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_68_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18487__SET_B repeater222/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10713__A2 _10704_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18805_ _18856_/CLK _18805_/D repeater231/X vssd1 vssd1 vccd1 vccd1 _18805_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__19560__RESET_B repeater269/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19785_ _20057_/CLK _19785_/D repeater203/X vssd1 vssd1 vccd1 vccd1 _19785_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_96_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16997_ _15963_/X _09535_/Y _17534_/S vssd1 vssd1 vccd1 vccd1 _16997_/X sky130_fd_sc_hd__mux2_1
XFILLER_84_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17353__S _17518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18736_ _20035_/CLK _18736_/D repeater244/X vssd1 vssd1 vccd1 vccd1 _18736_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_209_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15948_ _18131_/Q vssd1 vssd1 vccd1 vccd1 _15948_/Y sky130_fd_sc_hd__inv_2
XFILLER_225_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_64_HCLK_A clkbuf_opt_4_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18667_ _19812_/CLK _18667_/D repeater222/X vssd1 vssd1 vccd1 vccd1 _18667_/Q sky130_fd_sc_hd__dfstp_1
X_15879_ _19025_/Q vssd1 vssd1 vccd1 vccd1 _15879_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17618_ _20054_/Q _19728_/Q _17621_/S vssd1 vssd1 vccd1 vccd1 _17618_/X sky130_fd_sc_hd__mux2_1
X_18598_ _19865_/CLK _18598_/D repeater267/X vssd1 vssd1 vccd1 vccd1 _18598_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__14612__B1 hold320/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09095__A1 _20095_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17549_ _15860_/Y _18871_/Q _17550_/S vssd1 vssd1 vccd1 vccd1 _17549_/X sky130_fd_sc_hd__mux2_1
XFILLER_211_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16493__A _16493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17788__S0 _17923_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18851__CLK _18866_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19977__CLK _19984_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19219_ _19221_/CLK _19219_/D hold365/X vssd1 vssd1 vccd1 vccd1 _19219_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_118_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17528__S _17534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_247_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09805_ _09805_/A vssd1 vssd1 vccd1 vccd1 _09809_/A sky130_fd_sc_hd__inv_2
XANTENNA__17263__S _17524_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09736_ _09736_/A vssd1 vssd1 vccd1 vccd1 _09757_/B sky130_fd_sc_hd__inv_2
XFILLER_228_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09667_ _09753_/C _09754_/A _09667_/C _09757_/A vssd1 vssd1 vccd1 vccd1 _09668_/C
+ sky130_fd_sc_hd__or4_4
XFILLER_215_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09598_ _09598_/A vssd1 vssd1 vccd1 vccd1 _09598_/Y sky130_fd_sc_hd__inv_2
XPHY_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14603__B1 _14600_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17779__S0 _19647_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11560_ _11584_/C _11585_/A _11560_/C _11590_/A vssd1 vssd1 vccd1 vccd1 _11561_/C
+ sky130_fd_sc_hd__or4_4
XPHY_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10511_ _10511_/A _10514_/D vssd1 vssd1 vccd1 vccd1 _10521_/C sky130_fd_sc_hd__or2_1
XPHY_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11491_ _19609_/Q _11489_/Y _11227_/Y _11489_/A _11490_/X vssd1 vssd1 vccd1 vccd1
+ _19609_/D sky130_fd_sc_hd__o221a_1
XPHY_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12436__A _15867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13230_ _13230_/A vssd1 vssd1 vccd1 vccd1 _17584_/S sky130_fd_sc_hd__clkbuf_8
X_10442_ _10452_/A vssd1 vssd1 vccd1 vccd1 _10442_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_107_HCLK clkbuf_4_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _18718_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_164_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15747__A _19671_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17438__S _17568_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13161_ _13202_/A vssd1 vssd1 vccd1 vccd1 _13180_/A sky130_fd_sc_hd__inv_1
XFILLER_151_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10373_ _10367_/B _10372_/Y _10368_/X _10354_/X _10323_/A vssd1 vssd1 vccd1 vccd1
+ _10374_/A sky130_fd_sc_hd__o32a_1
XFILLER_3_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12112_ _19307_/Q _12106_/X _12030_/X _12108_/X vssd1 vssd1 vccd1 vccd1 _19307_/D
+ sky130_fd_sc_hd__a22o_1
X_13092_ _19189_/Q vssd1 vssd1 vccd1 vccd1 _13092_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11994__B _11998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16920_ _17473_/A0 _16632_/Y _17547_/S vssd1 vssd1 vccd1 vccd1 _16920_/X sky130_fd_sc_hd__mux2_1
X_12043_ _12043_/A vssd1 vssd1 vccd1 vccd1 _12043_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_172_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16851_ _15963_/X _12772_/Y _17534_/S vssd1 vssd1 vccd1 vccd1 _16851_/X sky130_fd_sc_hd__mux2_1
XANTENNA__16578__A _16688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17173__S _17543_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15802_ _18122_/Q vssd1 vssd1 vccd1 vccd1 _15802_/Y sky130_fd_sc_hd__inv_2
X_19570_ _19576_/CLK _19570_/D repeater282/X vssd1 vssd1 vccd1 vccd1 _19570_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_120_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16782_ _17473_/A0 _09900_/Y _17522_/S vssd1 vssd1 vccd1 vccd1 _16782_/X sky130_fd_sc_hd__mux2_1
XFILLER_207_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13994_ _18680_/Q vssd1 vssd1 vccd1 vccd1 _14011_/A sky130_fd_sc_hd__inv_2
XFILLER_74_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18521_ _19825_/CLK _18521_/D repeater223/X vssd1 vssd1 vccd1 vccd1 _18521_/Q sky130_fd_sc_hd__dfrtp_1
X_15733_ _18477_/Q vssd1 vssd1 vccd1 vccd1 _15733_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16728__D _16728_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12945_ _19267_/Q vssd1 vssd1 vccd1 vccd1 _12945_/Y sky130_fd_sc_hd__inv_2
XFILLER_233_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18953__RESET_B repeater257/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18452_ _18869_/CLK _18452_/D vssd1 vssd1 vccd1 vccd1 _18452_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_233_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15664_ _18609_/Q vssd1 vssd1 vccd1 vccd1 _15664_/Y sky130_fd_sc_hd__inv_2
XPHY_4260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12876_ _12876_/A _12994_/A vssd1 vssd1 vccd1 vccd1 _12877_/B sky130_fd_sc_hd__or2_1
XPHY_4271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17403_ _17402_/X _16173_/X _17567_/S vssd1 vssd1 vccd1 vccd1 _17403_/X sky130_fd_sc_hd__mux2_1
XFILLER_233_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14615_ _14642_/A _14668_/B _15145_/C vssd1 vssd1 vccd1 vccd1 _14617_/A sky130_fd_sc_hd__or3_4
XPHY_4293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18383_ _19637_/CLK _18383_/D vssd1 vssd1 vccd1 vccd1 _18383_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11827_ _19441_/Q _11821_/X _10866_/X _11822_/X vssd1 vssd1 vccd1 vccd1 _19441_/D
+ sky130_fd_sc_hd__a22o_1
X_15595_ _15598_/B _15594_/Y _15590_/X vssd1 vssd1 vccd1 vccd1 _15595_/X sky130_fd_sc_hd__o21a_1
XANTENNA__14070__A1 _19084_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17334_ _17333_/X _14050_/Y _17544_/S vssd1 vssd1 vccd1 vccd1 _17334_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12081__B1 _12080_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11758_ _11772_/A vssd1 vssd1 vccd1 vccd1 _11758_/X sky130_fd_sc_hd__clkbuf_2
X_14546_ _14547_/A vssd1 vssd1 vccd1 vccd1 _14546_/X sky130_fd_sc_hd__clkbuf_2
XPHY_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10709_ _15404_/A _10704_/B _10707_/Y _10708_/Y _10716_/S vssd1 vssd1 vccd1 vccd1
+ _10710_/A sky130_fd_sc_hd__o32a_1
XPHY_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17265_ _17264_/X _09435_/Y _17413_/S vssd1 vssd1 vccd1 vccd1 _17265_/X sky130_fd_sc_hd__mux2_1
X_11689_ _15823_/A _13252_/D vssd1 vssd1 vccd1 vccd1 _11691_/A sky130_fd_sc_hd__or2_2
X_14477_ _14490_/A _14477_/B _15009_/C vssd1 vssd1 vccd1 vccd1 _14479_/A sky130_fd_sc_hd__or3_4
X_19004_ _19595_/CLK _19004_/D hold346/A vssd1 vssd1 vccd1 vccd1 _19004_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_128_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16216_ _19443_/Q _17517_/S vssd1 vssd1 vccd1 vccd1 _16216_/Y sky130_fd_sc_hd__nand2_1
X_13428_ _13428_/A _13428_/B _13428_/C _13428_/D vssd1 vssd1 vccd1 vccd1 _13430_/C
+ sky130_fd_sc_hd__or4_4
XFILLER_162_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17196_ _17195_/X _11391_/Y _17548_/S vssd1 vssd1 vccd1 vccd1 _17196_/X sky130_fd_sc_hd__mux2_1
XFILLER_161_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17348__S _17474_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13359_ _20102_/Q _18848_/Q _13358_/Y _13333_/C vssd1 vssd1 vccd1 vccd1 _13359_/X
+ sky130_fd_sc_hd__o22a_1
X_16147_ _17420_/X _15997_/X _17423_/X _15998_/X _16146_/X vssd1 vssd1 vccd1 vccd1
+ _16147_/X sky130_fd_sc_hd__o221a_2
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16078_ _18141_/Q vssd1 vssd1 vccd1 vccd1 _16078_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19059__RESET_B repeater257/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19906_ _20006_/CLK _19906_/D repeater236/X vssd1 vssd1 vccd1 vccd1 _19906_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_142_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15029_ _18038_/Q _15023_/X _15000_/X _15025_/X vssd1 vssd1 vccd1 vccd1 _18038_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_216_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19837_ _19846_/CLK _19837_/D repeater272/X vssd1 vssd1 vccd1 vccd1 _19837_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_111_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11895__B1 hold317/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15086__B1 hold247/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16488__A _17568_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17083__S _17474_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19768_ _19771_/CLK _19768_/D repeater228/X vssd1 vssd1 vccd1 vccd1 _19768_/Q sky130_fd_sc_hd__dfstp_1
Xinput2 input2/A vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_1
XFILLER_56_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09521_ _19294_/Q vssd1 vssd1 vccd1 vccd1 _09521_/Y sky130_fd_sc_hd__inv_2
XFILLER_225_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18719_ _18727_/CLK _18719_/D repeater253/X vssd1 vssd1 vccd1 vccd1 _18719_/Q sky130_fd_sc_hd__dfrtp_1
X_19699_ _20051_/CLK _19699_/D repeater202/X vssd1 vssd1 vccd1 vccd1 _19699_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_232_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09452_ _19927_/Q vssd1 vssd1 vccd1 vccd1 _10043_/A sky130_fd_sc_hd__inv_2
XFILLER_25_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18694__RESET_B hold351/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09383_ _19934_/Q vssd1 vssd1 vccd1 vccd1 _10009_/A sky130_fd_sc_hd__inv_2
XFILLER_178_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12256__A _12370_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19829__RESET_B repeater271/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16670__B _16718_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17258__S _17545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19482__RESET_B repeater260/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11886__B1 _09030_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15077__B1 _14791_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11350__A2 _11328_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14824__B1 _14749_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09719_ _19984_/Q _09717_/Y _09740_/A _19413_/Q _09718_/X vssd1 vssd1 vccd1 vccd1
+ _09727_/B sky130_fd_sc_hd__o221a_1
X_10991_ _10991_/A vssd1 vssd1 vccd1 vccd1 _19663_/D sky130_fd_sc_hd__inv_2
XFILLER_215_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12730_ _14816_/A _12710_/A _12729_/X _12711_/A vssd1 vssd1 vccd1 vccd1 _18953_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_243_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12661_ _12677_/A vssd1 vssd1 vccd1 vccd1 _12661_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_42_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14052__A1 _19079_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11612_ _11612_/A vssd1 vssd1 vccd1 vccd1 _11612_/Y sky130_fd_sc_hd__inv_2
X_14400_ _18398_/Q _14394_/X hold324/X _14396_/X vssd1 vssd1 vccd1 vccd1 _18398_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15380_ _19796_/Q _10655_/X _19796_/Q _10655_/X vssd1 vssd1 vccd1 vccd1 _15380_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_12592_ _19036_/Q _12590_/X _12353_/X _12591_/X vssd1 vssd1 vccd1 vccd1 _19036_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11989__B _11998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11543_ _11543_/A vssd1 vssd1 vccd1 vccd1 _11617_/A sky130_fd_sc_hd__buf_2
XPHY_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14331_ _18435_/Q _14319_/A _14312_/X _14320_/A vssd1 vssd1 vccd1 vccd1 _18435_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11810__B1 _09058_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15001__B1 _15000_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17050_ _17049_/X _11312_/Y _17459_/S vssd1 vssd1 vccd1 vccd1 _17050_/X sky130_fd_sc_hd__mux2_1
X_14262_ _18472_/Q _14258_/X _12717_/X _14260_/X vssd1 vssd1 vccd1 vccd1 _18472_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_144_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11474_ _11474_/A _11474_/B vssd1 vssd1 vccd1 vccd1 _11514_/A sky130_fd_sc_hd__or2_1
XFILLER_183_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16001_ _17488_/X _15997_/X _17491_/X _15998_/X _16000_/X vssd1 vssd1 vccd1 vccd1
+ _16001_/X sky130_fd_sc_hd__o221a_2
X_13213_ _13213_/A vssd1 vssd1 vccd1 vccd1 _13213_/Y sky130_fd_sc_hd__inv_2
XFILLER_171_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17168__S _17547_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10425_ _12238_/A vssd1 vssd1 vccd1 vccd1 _10425_/X sky130_fd_sc_hd__buf_4
X_14193_ _14193_/A _14193_/B _14193_/C _14192_/X vssd1 vssd1 vccd1 vccd1 _14193_/X
+ sky130_fd_sc_hd__or4b_4
XANTENNA__17924__S0 _19647_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13144_ _13144_/A _13144_/B _13144_/C _13144_/D vssd1 vssd1 vccd1 vccd1 _13160_/C
+ sky130_fd_sc_hd__and4_1
X_10356_ _10356_/A vssd1 vssd1 vccd1 vccd1 _19862_/D sky130_fd_sc_hd__inv_2
XFILLER_152_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17952_ _20090_/CLK _17952_/D vssd1 vssd1 vccd1 vccd1 _17952_/Q sky130_fd_sc_hd__dfxtp_1
X_13075_ _13075_/A _13075_/B vssd1 vssd1 vccd1 vccd1 _13187_/A sky130_fd_sc_hd__or2_1
XFILLER_97_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10287_ _19874_/Q vssd1 vssd1 vccd1 vccd1 _15716_/A sky130_fd_sc_hd__inv_2
XANTENNA__16800__S _17542_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_239_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16903_ _16902_/X _18812_/Q _17386_/S vssd1 vssd1 vccd1 vccd1 _16903_/X sky130_fd_sc_hd__mux2_2
X_12026_ hold233/X vssd1 vssd1 vccd1 vccd1 _12026_/X sky130_fd_sc_hd__buf_4
XANTENNA__20057__RESET_B repeater204/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17883_ _16090_/Y _16091_/Y _16092_/Y _16093_/Y _17913_/S0 _19632_/Q vssd1 vssd1
+ vccd1 vccd1 _17883_/X sky130_fd_sc_hd__mux4_2
XFILLER_239_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19622_ _19920_/CLK _19622_/D repeater229/X vssd1 vssd1 vccd1 vccd1 _19622_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_93_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16834_ _16833_/X _12829_/Y _17386_/S vssd1 vssd1 vccd1 vccd1 _16834_/X sky130_fd_sc_hd__mux2_1
XFILLER_93_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19553_ _19582_/CLK _19553_/D repeater274/X vssd1 vssd1 vccd1 vccd1 _19553_/Q sky130_fd_sc_hd__dfrtp_1
X_16765_ _16764_/X _13553_/A _17386_/S vssd1 vssd1 vccd1 vccd1 _16765_/X sky130_fd_sc_hd__mux2_1
X_13977_ _18697_/Q vssd1 vssd1 vccd1 vccd1 _14027_/A sky130_fd_sc_hd__inv_2
XFILLER_207_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18504_ _19812_/CLK hold254/X repeater222/X vssd1 vssd1 vccd1 vccd1 _18505_/D sky130_fd_sc_hd__dfrtp_1
XFILLER_62_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15716_ _15716_/A _19871_/Q vssd1 vssd1 vccd1 vccd1 _15716_/Y sky130_fd_sc_hd__nor2_1
X_19484_ _19506_/CLK hold167/X repeater260/X vssd1 vssd1 vccd1 vccd1 _19484_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_46_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12928_ _12925_/Y _18945_/Q _12926_/Y _18939_/Q _12927_/X vssd1 vssd1 vccd1 vccd1
+ _12941_/A sky130_fd_sc_hd__o221a_1
XFILLER_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16696_ _16971_/X _16637_/X _17032_/X _16638_/X vssd1 vssd1 vccd1 vccd1 _16696_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_18_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18435_ _18435_/CLK _18435_/D vssd1 vssd1 vccd1 vccd1 _18435_/Q sky130_fd_sc_hd__dfxtp_1
X_15647_ _15666_/A _15647_/B vssd1 vssd1 vccd1 vccd1 _15647_/Y sky130_fd_sc_hd__nor2_1
XPHY_4090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12859_ _12859_/A _12859_/B _13021_/C vssd1 vssd1 vccd1 vccd1 _13001_/C sky130_fd_sc_hd__or3_1
XFILLER_21_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18366_ _18441_/CLK _18366_/D vssd1 vssd1 vccd1 vccd1 _18366_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15578_ _15610_/A _15578_/B vssd1 vssd1 vccd1 vccd1 _17664_/S sky130_fd_sc_hd__nor2_8
XFILLER_147_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17317_ _17473_/A0 _16370_/Y _17473_/S vssd1 vssd1 vccd1 vccd1 _17317_/X sky130_fd_sc_hd__mux2_1
XANTENNA__19993__RESET_B repeater192/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14529_ _19644_/Q _14545_/B _14571_/C vssd1 vssd1 vccd1 vccd1 _14532_/A sky130_fd_sc_hd__or3_4
XFILLER_147_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18297_ _18435_/CLK _18297_/D vssd1 vssd1 vccd1 vccd1 _18297_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12076__A hold289/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19922__RESET_B repeater230/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17248_ _16589_/Y _15514_/Y _17513_/S vssd1 vssd1 vccd1 vccd1 _17248_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16740__B1 _16837_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12357__A1 _19168_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17078__S _17487_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17179_ _17486_/A0 _13132_/Y _17543_/S vssd1 vssd1 vccd1 vccd1 _17179_/X sky130_fd_sc_hd__mux2_1
XANTENNA__17915__S0 _17918_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08952_ _18775_/Q vssd1 vssd1 vccd1 vccd1 _08952_/Y sky130_fd_sc_hd__inv_2
XFILLER_130_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18875__RESET_B repeater210/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18804__RESET_B repeater231/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17541__S _17541_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09504_ _19308_/Q vssd1 vssd1 vccd1 vccd1 _16547_/A sky130_fd_sc_hd__inv_2
XFILLER_25_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12293__B1 _12038_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_225_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16665__B _16668_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_225_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09435_ _19376_/Q vssd1 vssd1 vccd1 vccd1 _09435_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09366_ _20011_/Q vssd1 vssd1 vccd1 vccd1 _09472_/A sky130_fd_sc_hd__inv_2
XANTENNA__12045__B1 _11978_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09297_ _20042_/Q _09293_/X _09101_/X _09294_/X vssd1 vssd1 vccd1 vccd1 _20042_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19663__RESET_B repeater270/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19695__CLK _20051_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17906__S0 _17908_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10210_ _19653_/Q vssd1 vssd1 vccd1 vccd1 _10956_/B sky130_fd_sc_hd__inv_2
XFILLER_97_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11190_ _17714_/X _11184_/X _19617_/Q _11185_/X vssd1 vssd1 vccd1 vccd1 _19617_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17716__S _18546_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10141_ _16984_/X _10136_/X _19901_/Q _10138_/X vssd1 vssd1 vccd1 vccd1 _19901_/D
+ sky130_fd_sc_hd__o22a_1
X_10072_ _19923_/Q _10071_/Y _10057_/X _10040_/B vssd1 vssd1 vccd1 vccd1 _19923_/D
+ sky130_fd_sc_hd__o211a_1
X_13900_ _14003_/B vssd1 vssd1 vccd1 vccd1 _13925_/A sky130_fd_sc_hd__clkbuf_2
X_14880_ _18123_/Q _14872_/A _14713_/X _14873_/A vssd1 vssd1 vccd1 vccd1 _18123_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_47_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18545__RESET_B repeater232/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13831_ _13831_/A _13906_/A vssd1 vssd1 vccd1 vccd1 _13832_/B sky130_fd_sc_hd__or2_2
XFILLER_35_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17451__S _17536_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16550_ _19453_/Q _16622_/B vssd1 vssd1 vccd1 vccd1 _16550_/Y sky130_fd_sc_hd__nand2_1
XFILLER_189_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10974_ _19667_/Q _10973_/Y _10970_/X vssd1 vssd1 vccd1 vccd1 _19667_/D sky130_fd_sc_hd__o21a_1
X_13762_ _18747_/Q _13287_/X _13748_/A _13761_/X vssd1 vssd1 vccd1 vccd1 _18747_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_43_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15501_ _18570_/Q vssd1 vssd1 vccd1 vccd1 _15501_/Y sky130_fd_sc_hd__inv_2
XFILLER_71_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_189_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12713_ _18958_/Q vssd1 vssd1 vccd1 vccd1 _14806_/A sky130_fd_sc_hd__clkbuf_2
X_16481_ _16481_/A _16481_/B _16481_/C vssd1 vssd1 vccd1 vccd1 _16481_/X sky130_fd_sc_hd__and3_2
XFILLER_204_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13693_ _16435_/B _15169_/A vssd1 vssd1 vccd1 vccd1 _13694_/S sky130_fd_sc_hd__or2_1
XANTENNA__13280__A _13280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18220_ _18268_/CLK _18220_/D vssd1 vssd1 vccd1 vccd1 _18220_/Q sky130_fd_sc_hd__dfxtp_1
X_15432_ _19623_/Q _11168_/B _11169_/B vssd1 vssd1 vccd1 vccd1 _15432_/X sky130_fd_sc_hd__a21bo_1
XFILLER_188_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12644_ _12651_/A vssd1 vssd1 vccd1 vccd1 _12644_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_169_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18151_ _18165_/CLK _18151_/D vssd1 vssd1 vccd1 vccd1 _18151_/Q sky130_fd_sc_hd__dfxtp_1
X_15363_ _18503_/Q _14233_/B _17600_/S vssd1 vssd1 vccd1 vccd1 _15363_/X sky130_fd_sc_hd__a21o_1
X_12575_ _19047_/Q _12569_/X _12398_/X _12570_/X vssd1 vssd1 vccd1 vccd1 _19047_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16591__A _16688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17102_ _16466_/Y _18968_/Q _17459_/S vssd1 vssd1 vccd1 vccd1 _17102_/X sky130_fd_sc_hd__mux2_1
X_14314_ _14405_/A vssd1 vssd1 vccd1 vccd1 _14314_/X sky130_fd_sc_hd__buf_2
X_11526_ _19589_/Q _11528_/B _11521_/X _11470_/B vssd1 vssd1 vccd1 vccd1 _19589_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18082_ _18260_/CLK _18082_/D vssd1 vssd1 vccd1 vccd1 _18082_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15294_ _15294_/A vssd1 vssd1 vccd1 vccd1 _17756_/S sky130_fd_sc_hd__inv_2
XPHY_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17033_ _17486_/A0 _13136_/Y _17543_/S vssd1 vssd1 vccd1 vccd1 _17033_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11457_ _11457_/A _11457_/B _11457_/C _11457_/D vssd1 vssd1 vccd1 vccd1 _11566_/B
+ sky130_fd_sc_hd__and4_1
X_14245_ _14245_/A _15821_/B _14245_/C _14245_/D vssd1 vssd1 vccd1 vccd1 _14246_/S
+ sky130_fd_sc_hd__or4_4
XFILLER_183_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10408_ _10989_/A vssd1 vssd1 vccd1 vccd1 _10408_/X sky130_fd_sc_hd__buf_1
X_14176_ _19113_/Q vssd1 vssd1 vccd1 vccd1 _16617_/A sky130_fd_sc_hd__inv_2
X_11388_ _11576_/A _19143_/Q _11571_/A _19138_/Q _11387_/X vssd1 vssd1 vccd1 vccd1
+ _11389_/D sky130_fd_sc_hd__o221a_1
XANTENNA_output89_A _16614_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10339_ _10332_/A _10336_/X _10332_/B _10336_/B vssd1 vssd1 vccd1 vccd1 _19866_/D
+ sky130_fd_sc_hd__o22ai_1
X_13127_ _13113_/X _13127_/B _13127_/C _13127_/D vssd1 vssd1 vccd1 vccd1 _13160_/B
+ sky130_fd_sc_hd__and4b_1
X_18984_ _19608_/CLK _18984_/D hold355/X vssd1 vssd1 vccd1 vccd1 _18984_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_98_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17935_ _18465_/CLK _17935_/D vssd1 vssd1 vccd1 vccd1 _17935_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13058_ _18888_/Q vssd1 vssd1 vccd1 vccd1 _13061_/A sky130_fd_sc_hd__inv_2
XANTENNA__12511__A1 _19078_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12009_ _12016_/A vssd1 vssd1 vccd1 vccd1 _12009_/X sky130_fd_sc_hd__buf_1
XFILLER_66_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17866_ _16181_/Y _16182_/Y _16183_/Y _16184_/Y _17908_/S0 _18759_/Q vssd1 vssd1
+ vccd1 vccd1 _17866_/X sky130_fd_sc_hd__mux4_2
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater149 _15963_/X vssd1 vssd1 vccd1 vccd1 _17486_/A0 sky130_fd_sc_hd__clkbuf_16
X_16817_ _16816_/X _13373_/Y _17535_/S vssd1 vssd1 vccd1 vccd1 _16817_/X sky130_fd_sc_hd__mux2_1
X_19605_ _19609_/CLK _19605_/D hold359/X vssd1 vssd1 vccd1 vccd1 _19605_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_66_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17797_ _18328_/Q _18008_/Q _18312_/Q _18304_/Q _17923_/S0 _19646_/Q vssd1 vssd1
+ vccd1 vccd1 _17797_/X sky130_fd_sc_hd__mux4_2
XFILLER_242_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17361__S _17487_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19536_ _19540_/CLK _19536_/D repeater221/X vssd1 vssd1 vccd1 vccd1 _19536_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_207_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12275__B1 _12092_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16748_ _16042_/Y _18757_/Q _18869_/Q _15956_/Y vssd1 vssd1 vccd1 vccd1 _16748_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_34_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10825__A1 _10448_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19467_ _19470_/CLK _19467_/D repeater274/X vssd1 vssd1 vccd1 vccd1 _19467_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_222_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16679_ _18985_/Q vssd1 vssd1 vccd1 vccd1 _16679_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09220_ _18651_/Q vssd1 vssd1 vccd1 vccd1 _09220_/Y sky130_fd_sc_hd__inv_2
XFILLER_210_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18418_ _18795_/CLK _18418_/D vssd1 vssd1 vccd1 vccd1 _18418_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12027__B1 _12026_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_119_HCLK_A clkbuf_opt_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19398_ _19905_/CLK _19398_/D repeater191/X vssd1 vssd1 vccd1 vccd1 _19398_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_21_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09151_ _09151_/A _09151_/B vssd1 vssd1 vccd1 vccd1 _09151_/Y sky130_fd_sc_hd__nor2_1
X_18349_ _18959_/CLK _18349_/D vssd1 vssd1 vccd1 vccd1 _18349_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09082_ _10446_/A vssd1 vssd1 vccd1 vccd1 _09082_/X sky130_fd_sc_hd__buf_4
XFILLER_238_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_190_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput60 input60/A vssd1 vssd1 vccd1 vccd1 input60/X sky130_fd_sc_hd__clkbuf_8
Xinput71 input71/A vssd1 vssd1 vccd1 vccd1 input71/X sky130_fd_sc_hd__buf_2
XFILLER_190_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17536__S _17536_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15845__A _15858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09984_ _09984_/A vssd1 vssd1 vccd1 vccd1 _09987_/A sky130_fd_sc_hd__inv_2
XFILLER_107_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_3_1_0_HCLK clkbuf_3_1_0_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_3_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_08935_ _19862_/Q _18782_/Q _10328_/A _08934_/Y vssd1 vssd1 vccd1 vccd1 _08935_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_96_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17271__S _17523_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12266__B1 _12076_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_199_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14196__A _19112_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09418_ _19393_/Q vssd1 vssd1 vccd1 vccd1 _09418_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19844__RESET_B repeater270/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12018__B1 hold314/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10690_ _10819_/A _12370_/B _13279_/C vssd1 vssd1 vccd1 vccd1 _15858_/D sky130_fd_sc_hd__or3_4
XANTENNA__13215__C1 _13176_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_240_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09349_ _20028_/Q vssd1 vssd1 vccd1 vccd1 _09488_/A sky130_fd_sc_hd__inv_2
XFILLER_12_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12360_ _19165_/Q _12352_/X _12296_/X _12354_/X vssd1 vssd1 vccd1 vccd1 _19165_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11241__B2 _18997_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11311_ _18965_/Q vssd1 vssd1 vccd1 vccd1 _11311_/Y sky130_fd_sc_hd__inv_2
XFILLER_148_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12291_ _12300_/A vssd1 vssd1 vccd1 vccd1 _12291_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_180_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12444__A _12458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14030_ _14030_/A _14030_/B vssd1 vssd1 vccd1 vccd1 _14031_/B sky130_fd_sc_hd__or2_1
XFILLER_180_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11242_ _19588_/Q vssd1 vssd1 vccd1 vccd1 _11468_/A sky130_fd_sc_hd__inv_2
XANTENNA__11544__A2 _11617_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17446__S _17534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11173_ _11173_/A _18526_/D _11173_/C vssd1 vssd1 vccd1 vccd1 _11173_/X sky130_fd_sc_hd__or3_4
XANTENNA__18797__RESET_B repeater258/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10124_ _18573_/Q _18574_/Q _10124_/C _15537_/A vssd1 vssd1 vccd1 vccd1 _10125_/B
+ sky130_fd_sc_hd__or4_1
XANTENNA__18726__RESET_B repeater253/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15981_ _19757_/Q vssd1 vssd1 vccd1 vccd1 _15981_/Y sky130_fd_sc_hd__inv_2
X_17720_ _15420_/Y _19521_/Q _18546_/D vssd1 vssd1 vccd1 vccd1 _17720_/X sky130_fd_sc_hd__mux2_1
X_10055_ _10055_/A vssd1 vssd1 vccd1 vccd1 _10055_/Y sky130_fd_sc_hd__inv_2
X_14932_ _18093_/Q _14920_/X _14931_/X _14923_/X vssd1 vssd1 vccd1 vccd1 _18093_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_75_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_248_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17651_ _15631_/X _19038_/Q _17655_/S vssd1 vssd1 vccd1 vccd1 _18601_/D sky130_fd_sc_hd__mux2_1
XFILLER_75_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14863_ _18135_/Q _14858_/X _14705_/X _14860_/X vssd1 vssd1 vccd1 vccd1 _18135_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_output127_A _15779_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16640__C1 _16639_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16602_ _19043_/Q vssd1 vssd1 vccd1 vccd1 _16602_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17181__S _17542_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13814_ _13964_/A _13912_/A vssd1 vssd1 vccd1 vccd1 _13815_/B sky130_fd_sc_hd__or2_2
X_17582_ _15395_/X _19525_/Q _17584_/S vssd1 vssd1 vccd1 vccd1 _17582_/X sky130_fd_sc_hd__mux2_1
X_14794_ _18173_/Q _14785_/X _14793_/X _14787_/X vssd1 vssd1 vccd1 vccd1 _18173_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_91_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19321_ _19324_/CLK _19321_/D repeater213/X vssd1 vssd1 vccd1 vccd1 _19321_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_204_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16533_ _16504_/X _16527_/X _16529_/X _16532_/X vssd1 vssd1 vccd1 vccd1 _16533_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_90_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13745_ _18747_/Q vssd1 vssd1 vccd1 vccd1 _13745_/Y sky130_fd_sc_hd__inv_2
XFILLER_232_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10957_ _10957_/A _11009_/A vssd1 vssd1 vccd1 vccd1 _11005_/A sky130_fd_sc_hd__or2_1
XFILLER_16_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19252_ _19324_/CLK _19252_/D repeater237/X vssd1 vssd1 vccd1 vccd1 _19252_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_43_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13206__C1 _13202_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16464_ _11742_/A _16458_/X _16460_/X _16462_/X _16463_/X vssd1 vssd1 vccd1 vccd1
+ _16464_/X sky130_fd_sc_hd__o2111a_1
X_13676_ hold331/X vssd1 vssd1 vccd1 vccd1 _13676_/X sky130_fd_sc_hd__buf_2
XFILLER_189_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10888_ _19696_/Q _10875_/X _10863_/X _10879_/X vssd1 vssd1 vccd1 vccd1 _19696_/D
+ sky130_fd_sc_hd__a22o_1
X_18203_ _18460_/CLK _18203_/D vssd1 vssd1 vccd1 vccd1 _18203_/Q sky130_fd_sc_hd__dfxtp_1
X_15415_ _15419_/A _17573_/X vssd1 vssd1 vccd1 vccd1 _18539_/D sky130_fd_sc_hd__and2_1
XPHY_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12627_ _19015_/Q _12622_/X _12396_/X _12623_/X vssd1 vssd1 vccd1 vccd1 _19015_/D
+ sky130_fd_sc_hd__a22o_1
X_19183_ _19293_/CLK _19183_/D repeater187/X vssd1 vssd1 vccd1 vccd1 _19183_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16395_ _17320_/X _16148_/X _17329_/X _16394_/X vssd1 vssd1 vccd1 vccd1 _16395_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18134_ _18137_/CLK _18134_/D vssd1 vssd1 vccd1 vccd1 _18134_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15346_ _18495_/Q _14225_/B _14226_/B vssd1 vssd1 vccd1 vccd1 _15346_/X sky130_fd_sc_hd__a21bo_1
XPHY_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12558_ _12659_/A _12558_/B vssd1 vssd1 vccd1 vccd1 _12598_/A sky130_fd_sc_hd__or2_4
XPHY_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11509_ _19599_/Q _11508_/Y _11504_/X _11480_/B vssd1 vssd1 vccd1 vccd1 _19599_/D
+ sky130_fd_sc_hd__o211a_1
X_18065_ _18465_/CLK _18065_/D vssd1 vssd1 vccd1 vccd1 _18065_/Q sky130_fd_sc_hd__dfxtp_1
X_15277_ _10909_/A _18635_/Q _15229_/B _15276_/X vssd1 vssd1 vccd1 vccd1 _15277_/Y
+ sky130_fd_sc_hd__a31oi_4
XFILLER_144_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12489_ _12505_/A vssd1 vssd1 vccd1 vccd1 _12489_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__14182__B1 _19112_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold129 hold354/X vssd1 vssd1 vccd1 vccd1 hold353/A sky130_fd_sc_hd__dlygate4sd3_1
X_17016_ _17015_/X _14073_/Y _17490_/S vssd1 vssd1 vccd1 vccd1 _17016_/X sky130_fd_sc_hd__mux2_2
X_14228_ _18498_/Q _14228_/B vssd1 vssd1 vccd1 vccd1 _14229_/B sky130_fd_sc_hd__or2_1
XFILLER_99_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20072__RESET_B repeater207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17356__S _17530_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14159_ _19107_/Q vssd1 vssd1 vccd1 vccd1 _16543_/A sky130_fd_sc_hd__inv_2
XANTENNA__20001__RESET_B repeater192/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18967_ _19137_/CLK _18967_/D hold348/X vssd1 vssd1 vccd1 vccd1 _18967_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_112_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12496__B1 _12384_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17918_ _17935_/Q _18457_/Q _18465_/Q _18065_/Q _17918_/S0 _18750_/Q vssd1 vssd1
+ vccd1 vccd1 _17918_/X sky130_fd_sc_hd__mux4_2
XFILLER_85_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18898_ _18908_/CLK _18898_/D repeater188/X vssd1 vssd1 vccd1 vccd1 _18898_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_239_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17849_ _17845_/X _17846_/X _17847_/X _17848_/X _18760_/Q _18761_/Q vssd1 vssd1 vccd1
+ vccd1 _17849_/X sky130_fd_sc_hd__mux4_2
XFILLER_66_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14237__B2 _17600_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17091__S _17487_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13913__A _19125_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_240_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19519_ _19859_/CLK hold219/X repeater262/X vssd1 vssd1 vccd1 vccd1 _19519_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_240_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09203_ _09203_/A _09205_/A _09205_/B vssd1 vssd1 vccd1 vccd1 _09203_/X sky130_fd_sc_hd__or3_2
XFILLER_194_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09134_ _09113_/A _09131_/X _09136_/B _09133_/X vssd1 vssd1 vccd1 vccd1 _20089_/D
+ sky130_fd_sc_hd__o2bb2a_1
X_09065_ _20104_/Q _09053_/X _09064_/X _09055_/X vssd1 vssd1 vccd1 vccd1 _20104_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_162_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_140_HCLK clkbuf_4_3_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19846_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_104_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17266__S _17414_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19733__CLK _20051_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09967_ _09967_/A vssd1 vssd1 vccd1 vccd1 _09967_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08918_ _20123_/Q _20124_/Q vssd1 vssd1 vccd1 vccd1 _08919_/A sky130_fd_sc_hd__nor2_1
X_20087_ _20090_/CLK _20087_/D repeater205/X vssd1 vssd1 vccd1 vccd1 _20087_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_hold272_A HWDATA[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_246_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09898_ _19952_/Q _19344_/Q _09860_/A _09897_/Y vssd1 vssd1 vccd1 vccd1 _09898_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_4601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12239__B1 _12238_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11860_ _13642_/B vssd1 vssd1 vccd1 vccd1 _11861_/B sky130_fd_sc_hd__inv_2
XPHY_4634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10811_ _17615_/X _10808_/X _19732_/Q _10810_/X vssd1 vssd1 vccd1 vccd1 _19732_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_60_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11791_ _19467_/Q _11784_/X _09025_/X _11787_/X vssd1 vssd1 vccd1 vccd1 _19467_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_214_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12439__A _15769_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13530_ _13530_/A _13530_/B vssd1 vssd1 vccd1 vccd1 _13607_/A sky130_fd_sc_hd__or2_1
XFILLER_25_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10742_ _10742_/A vssd1 vssd1 vccd1 vccd1 _10743_/A sky130_fd_sc_hd__inv_2
XPHY_3988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13461_ _13428_/D _13336_/B _13459_/Y _13437_/X vssd1 vssd1 vccd1 vccd1 _18849_/D
+ sky130_fd_sc_hd__a211oi_2
X_10673_ _17736_/X _10669_/X _19789_/Q _10670_/X vssd1 vssd1 vccd1 vccd1 _19789_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_158_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_102_HCLK_A clkbuf_4_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15200_ _15201_/B vssd1 vssd1 vccd1 vccd1 _16957_/S sky130_fd_sc_hd__inv_2
X_12412_ _12427_/A vssd1 vssd1 vccd1 vccd1 _12412_/X sky130_fd_sc_hd__buf_1
X_16180_ _17973_/Q vssd1 vssd1 vccd1 vccd1 _16180_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12411__B1 _12410_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13392_ _20111_/Q _13428_/B _20113_/Q _13431_/D vssd1 vssd1 vccd1 vccd1 _13392_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_138_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15131_ _17970_/Q _15123_/A _14935_/X _15124_/A vssd1 vssd1 vccd1 vccd1 _17970_/D
+ sky130_fd_sc_hd__a22o_1
X_12343_ _19174_/Q _12341_/X _12107_/X _12342_/X vssd1 vssd1 vccd1 vccd1 _19174_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_181_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15062_ _18017_/Q _15059_/X _14802_/A _15061_/X vssd1 vssd1 vccd1 vccd1 _18017_/D
+ sky130_fd_sc_hd__a22o_1
X_12274_ _19216_/Q _12269_/X _12090_/X _12270_/X vssd1 vssd1 vccd1 vccd1 _19216_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18907__RESET_B repeater188/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11225_ _19005_/Q vssd1 vssd1 vccd1 vccd1 _11225_/Y sky130_fd_sc_hd__inv_2
X_14013_ _14013_/A _14013_/B vssd1 vssd1 vccd1 vccd1 _14014_/B sky130_fd_sc_hd__or2_2
XANTENNA__17176__S _17543_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19870_ _19905_/CLK _19870_/D repeater210/X vssd1 vssd1 vccd1 vccd1 _19870_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__10725__B1 _10451_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11156_ _18547_/Q vssd1 vssd1 vccd1 vccd1 _11175_/A sky130_fd_sc_hd__inv_2
X_18821_ _18827_/CLK _18821_/D repeater231/X vssd1 vssd1 vccd1 vccd1 _18821_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__18560__RESET_B repeater193/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10107_ _10107_/A _10107_/B _10107_/C vssd1 vssd1 vccd1 vccd1 _19907_/D sky130_fd_sc_hd__nor3_1
XFILLER_0_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18752_ _19900_/CLK _18752_/D repeater195/X vssd1 vssd1 vccd1 vccd1 _18752_/Q sky130_fd_sc_hd__dfrtp_2
X_11087_ _15222_/A _19225_/Q _15232_/C vssd1 vssd1 vccd1 vccd1 _12545_/A sky130_fd_sc_hd__or3_4
X_15964_ _19402_/Q vssd1 vssd1 vccd1 vccd1 _15964_/Y sky130_fd_sc_hd__inv_2
X_17703_ _19815_/Q _19757_/Q _18548_/Q vssd1 vssd1 vccd1 vccd1 _17703_/X sky130_fd_sc_hd__mux2_1
X_10038_ _10038_/A _10038_/B vssd1 vssd1 vccd1 vccd1 _10071_/A sky130_fd_sc_hd__or2_1
XFILLER_49_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14915_ _18101_/Q _14908_/X _14709_/X _14910_/X vssd1 vssd1 vccd1 vccd1 _18101_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_208_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18683_ _18686_/CLK _18683_/D repeater252/X vssd1 vssd1 vccd1 vccd1 _18683_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_236_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15895_ _15895_/A vssd1 vssd1 vccd1 vccd1 _16530_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_75_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16613__C1 _16612_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17634_ _15702_/Y _19055_/Q _17664_/S vssd1 vssd1 vccd1 vccd1 _18618_/D sky130_fd_sc_hd__mux2_1
X_14846_ _14846_/A vssd1 vssd1 vccd1 vccd1 _14847_/A sky130_fd_sc_hd__inv_2
XFILLER_236_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_21_HCLK clkbuf_4_3_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20036_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_189_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17565_ _17564_/X _16747_/A _17565_/S vssd1 vssd1 vccd1 vccd1 _17565_/X sky130_fd_sc_hd__mux2_1
XFILLER_63_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14777_ _18182_/Q _14771_/X _14723_/X _14773_/X vssd1 vssd1 vccd1 vccd1 _18182_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_189_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11989_ _15881_/B _11998_/A vssd1 vssd1 vccd1 vccd1 _11990_/S sky130_fd_sc_hd__or2_1
XFILLER_90_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19304_ _20035_/CLK _19304_/D repeater242/X vssd1 vssd1 vccd1 vccd1 _19304_/Q sky130_fd_sc_hd__dfrtp_4
X_16516_ _16504_/X _16507_/X _16511_/X _16515_/X vssd1 vssd1 vccd1 vccd1 _16516_/Y
+ sky130_fd_sc_hd__o211ai_4
X_13728_ _14366_/A _14366_/B _17763_/X _13291_/Y _13727_/X vssd1 vssd1 vccd1 vccd1
+ _18756_/D sky130_fd_sc_hd__a41o_1
X_17496_ _17495_/X _20037_/Q _19497_/Q vssd1 vssd1 vccd1 vccd1 _17496_/X sky130_fd_sc_hd__mux2_1
XFILLER_232_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19235_ _19282_/CLK _19235_/D repeater216/X vssd1 vssd1 vccd1 vccd1 _19235_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_176_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16447_ _16443_/Y _15971_/A _15336_/A _15973_/X _16446_/X vssd1 vssd1 vccd1 vccd1
+ _16447_/X sky130_fd_sc_hd__o221a_1
X_13659_ _18787_/Q _13656_/X hold233/X _13658_/X vssd1 vssd1 vccd1 vccd1 _18787_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16392__B2 _15999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19166_ _19214_/CLK _19166_/D hold367/X vssd1 vssd1 vccd1 vccd1 _19166_/Q sky130_fd_sc_hd__dfrtp_2
X_16378_ _16375_/Y _15971_/A _15330_/A _15973_/X _16377_/X vssd1 vssd1 vccd1 vccd1
+ _16378_/X sky130_fd_sc_hd__o221a_1
XFILLER_185_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_163_HCLK clkbuf_4_0_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19506_/CLK sky130_fd_sc_hd__clkbuf_16
X_18117_ _18145_/CLK _18117_/D vssd1 vssd1 vccd1 vccd1 _18117_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12953__A1 _12952_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15329_ _18480_/Q vssd1 vssd1 vccd1 vccd1 _15832_/A sky130_fd_sc_hd__inv_2
X_19097_ _19585_/CLK _19097_/D hold365/X vssd1 vssd1 vccd1 vccd1 _19097_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_24_HCLK_A clkbuf_4_9_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_87_HCLK_A clkbuf_4_13_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18048_ _18473_/CLK _18048_/D vssd1 vssd1 vccd1 vccd1 _18048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17086__S _17545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10716__A0 _10715_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20010_ _20091_/CLK _20010_/D repeater240/X vssd1 vssd1 vccd1 vccd1 _20010_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_98_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09821_ _19965_/Q vssd1 vssd1 vccd1 vccd1 _09873_/A sky130_fd_sc_hd__inv_2
XFILLER_113_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19999_ _20003_/CLK _19999_/D repeater185/X vssd1 vssd1 vccd1 vccd1 _19999_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12469__B1 hold256/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09752_ _09752_/A _09752_/B vssd1 vssd1 vccd1 vccd1 _09765_/A sky130_fd_sc_hd__or2_2
XFILLER_228_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09683_ _09640_/A _19401_/Q _19972_/Q _09680_/Y _09682_/X vssd1 vssd1 vccd1 vccd1
+ _09689_/C sky130_fd_sc_hd__o221a_1
XFILLER_227_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16604__C1 _16603_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19436__RESET_B repeater210/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20113__CLK _20115_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16907__A0 _16906_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12641__B1 _12030_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16673__B _16673_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18160__CLK _18198_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09117_ _17604_/X vssd1 vssd1 vccd1 vccd1 _09162_/A sky130_fd_sc_hd__inv_2
XFILLER_191_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09048_ _20110_/Q _09041_/X hold317/X _09043_/X vssd1 vssd1 vccd1 vccd1 _20110_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_191_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11010_ _19657_/Q _11010_/B vssd1 vssd1 vccd1 vccd1 _11010_/Y sky130_fd_sc_hd__nor2_1
XFILLER_49_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_44_HCLK clkbuf_opt_2_HCLK/A vssd1 vssd1 vccd1 vccd1 _19544_/CLK sky130_fd_sc_hd__clkbuf_16
X_12961_ _12891_/A _12891_/B _12892_/Y _13027_/C vssd1 vssd1 vccd1 vccd1 _18949_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_46_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14700_ _14700_/A vssd1 vssd1 vccd1 vccd1 _14701_/A sky130_fd_sc_hd__inv_2
X_11912_ _19409_/Q _11905_/X _11911_/X _11906_/X vssd1 vssd1 vccd1 vccd1 _19409_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_233_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15680_ _18613_/Q vssd1 vssd1 vccd1 vccd1 _15683_/A sky130_fd_sc_hd__inv_2
XPHY_4420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12892_ _12892_/A vssd1 vssd1 vccd1 vccd1 _12892_/Y sky130_fd_sc_hd__inv_2
XPHY_4431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19177__RESET_B repeater212/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16610__A2 _16394_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14631_ _14631_/A vssd1 vssd1 vccd1 vccd1 _14632_/A sky130_fd_sc_hd__inv_2
XPHY_4453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11843_ _14680_/B vssd1 vssd1 vccd1 vccd1 _16055_/A sky130_fd_sc_hd__clkbuf_4
XPHY_4464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17350_ _17349_/X _15467_/A _17518_/S vssd1 vssd1 vccd1 vccd1 _17350_/X sky130_fd_sc_hd__mux2_1
XPHY_4497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12632__B1 _12404_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14562_ _18304_/Q _14558_/X _14535_/X _14560_/X vssd1 vssd1 vccd1 vccd1 _18304_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11774_ hold206/X _11771_/X _19474_/Q _11772_/X vssd1 vssd1 vccd1 vccd1 hold208/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_201_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16301_ _19690_/Q vssd1 vssd1 vccd1 vccd1 _16301_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16583__B _16583_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_241_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17797__S1 _19646_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13513_ _14628_/B _18758_/Q _14641_/B _13704_/B _17759_/X vssd1 vssd1 vccd1 vccd1
+ _13513_/Y sky130_fd_sc_hd__o221ai_1
X_10725_ _19770_/Q _10720_/X _10451_/X _10722_/X vssd1 vssd1 vccd1 vccd1 _19770_/D
+ sky130_fd_sc_hd__a22o_1
X_17281_ _17280_/X _16501_/Y _17385_/S vssd1 vssd1 vccd1 vccd1 _17281_/X sky130_fd_sc_hd__mux2_1
X_14493_ _14493_/A vssd1 vssd1 vccd1 vccd1 _14493_/X sky130_fd_sc_hd__clkbuf_2
X_19020_ _19609_/CLK _19020_/D hold357/X vssd1 vssd1 vccd1 vccd1 _19020_/Q sky130_fd_sc_hd__dfrtp_1
X_16232_ _16227_/Y _16053_/X _16228_/Y _15828_/A _16231_/X vssd1 vssd1 vccd1 vccd1
+ _16232_/X sky130_fd_sc_hd__o221a_1
XFILLER_158_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11801__A _11801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13444_ _18860_/Q _13442_/Y _13348_/B _13443_/X vssd1 vssd1 vccd1 vccd1 _18860_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__19779__CLK _19780_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10656_ _19672_/Q vssd1 vssd1 vccd1 vccd1 _10658_/A sky130_fd_sc_hd__inv_2
XFILLER_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16163_ _18350_/Q vssd1 vssd1 vccd1 vccd1 _16163_/Y sky130_fd_sc_hd__inv_2
X_10587_ _19797_/Q vssd1 vssd1 vccd1 vccd1 _10589_/B sky130_fd_sc_hd__inv_2
X_13375_ _20093_/Q _18839_/Q _13374_/Y _13322_/B vssd1 vssd1 vccd1 vccd1 _13375_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_182_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16803__S _17482_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14137__B1 _18681_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15114_ _17983_/Q _15110_/X _14925_/X _15112_/X vssd1 vssd1 vccd1 vccd1 _17983_/D
+ sky130_fd_sc_hd__a22o_1
X_12326_ _19185_/Q _12318_/X _12080_/X _12321_/X vssd1 vssd1 vccd1 vccd1 _19185_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_5_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16094_ _19845_/Q vssd1 vssd1 vccd1 vccd1 _16094_/Y sky130_fd_sc_hd__inv_2
XFILLER_126_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19922_ _19927_/CLK _19922_/D repeater230/X vssd1 vssd1 vccd1 vccd1 _19922_/Q sky130_fd_sc_hd__dfrtp_1
X_15045_ _18026_/Q _15036_/A _15020_/X _15037_/A vssd1 vssd1 vccd1 vccd1 _18026_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_181_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12257_ _12257_/A _15911_/A vssd1 vssd1 vccd1 vccd1 _12487_/B sky130_fd_sc_hd__or2_2
XFILLER_141_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11208_ _19020_/Q vssd1 vssd1 vccd1 vccd1 _11208_/Y sky130_fd_sc_hd__inv_2
X_12188_ _12228_/A vssd1 vssd1 vccd1 vccd1 _12205_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_19853_ _19865_/CLK _19853_/D repeater267/X vssd1 vssd1 vccd1 vccd1 _19853_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_69_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18804_ _18856_/CLK _18804_/D repeater231/X vssd1 vssd1 vccd1 vccd1 _18804_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__19947__RESET_B hold371/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11139_ _11139_/A vssd1 vssd1 vccd1 vccd1 _11139_/Y sky130_fd_sc_hd__inv_2
XFILLER_205_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19784_ _20057_/CLK _19784_/D repeater203/X vssd1 vssd1 vccd1 vccd1 _19784_/Q sky130_fd_sc_hd__dfrtp_1
X_16996_ _16673_/Y _15675_/Y _17318_/S vssd1 vssd1 vccd1 vccd1 _16996_/X sky130_fd_sc_hd__mux2_2
XFILLER_68_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15947_ _18219_/Q vssd1 vssd1 vccd1 vccd1 _15947_/Y sky130_fd_sc_hd__inv_2
X_18735_ _19224_/CLK _18735_/D repeater186/X vssd1 vssd1 vccd1 vccd1 _18735_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_225_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13463__A _13483_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18666_ _19544_/CLK _18666_/D repeater222/X vssd1 vssd1 vccd1 vccd1 _18666_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_224_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15878_ _19400_/Q _15878_/B vssd1 vssd1 vccd1 vccd1 _15878_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__18183__CLK _18198_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17617_ _20055_/Q _19729_/Q _17621_/S vssd1 vssd1 vccd1 vccd1 _17617_/X sky130_fd_sc_hd__mux2_1
X_14829_ _18155_/Q _14821_/A _14780_/X _14822_/A vssd1 vssd1 vccd1 vccd1 _18155_/D
+ sky130_fd_sc_hd__a22o_1
X_18597_ _19157_/CLK _18597_/D repeater267/X vssd1 vssd1 vccd1 vccd1 _18597_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_51_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17548_ _17547_/X _15861_/Y _17548_/S vssd1 vssd1 vccd1 vccd1 _17548_/X sky130_fd_sc_hd__mux2_1
XFILLER_205_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17788__S1 _19646_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17479_ _17478_/X _09849_/A _17518_/S vssd1 vssd1 vccd1 vccd1 _17479_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11711__A _11731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14376__B1 _14312_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19218_ _19221_/CLK _19218_/D hold365/X vssd1 vssd1 vccd1 vccd1 _19218_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_146_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14193__D_N _14192_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19149_ _19576_/CLK _19149_/D repeater281/X vssd1 vssd1 vccd1 vccd1 _19149_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_157_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_246_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_67_HCLK clkbuf_opt_3_HCLK/A vssd1 vssd1 vccd1 vccd1 _19927_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__17544__S _17544_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09804_ _19977_/Q _09803_/Y _09790_/B _09731_/X vssd1 vssd1 vccd1 vccd1 _19977_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_101_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19617__RESET_B repeater230/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16668__B _16668_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09735_ _19364_/Q _09735_/B vssd1 vssd1 vccd1 vccd1 _09736_/A sky130_fd_sc_hd__or2_1
XFILLER_86_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09666_ _09739_/B _09666_/B _09666_/C vssd1 vssd1 vccd1 vccd1 _09757_/A sky130_fd_sc_hd__or3_4
XFILLER_243_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09597_ _09478_/A _09478_/B _09595_/Y _09587_/X vssd1 vssd1 vccd1 vccd1 _20018_/D
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__16684__A _16684_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11417__B2 _19146_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold235_A HWDATA[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17779__S1 _19648_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20104__RESET_B repeater233/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10510_ _11651_/A _11649_/A _10736_/A _11653_/A vssd1 vssd1 vccd1 vccd1 _10537_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_195_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11490_ _11504_/A vssd1 vssd1 vccd1 vccd1 _11490_/X sky130_fd_sc_hd__clkbuf_2
XPHY_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10441_ _10450_/A vssd1 vssd1 vccd1 vccd1 _10441_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__17719__S _18546_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17305__A0 _15768_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10372_ _19857_/Q _10372_/B vssd1 vssd1 vccd1 vccd1 _10372_/Y sky130_fd_sc_hd__nor2_1
X_13160_ _13160_/A _13160_/B _13160_/C _13160_/D vssd1 vssd1 vccd1 vccd1 _13202_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_200_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20009__CLK _20013_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12111_ _19308_/Q _12106_/X _12028_/X _12108_/X vssd1 vssd1 vccd1 vccd1 _19308_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18056__CLK _18169_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13091_ _18918_/Q vssd1 vssd1 vccd1 vccd1 _13091_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_70_HCLK_A clkbuf_opt_2_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12042_ _19338_/Q _12034_/X _11975_/X _12036_/X vssd1 vssd1 vccd1 vccd1 _19338_/D
+ sky130_fd_sc_hd__a22o_1
Xhold290 HWDATA[29] vssd1 vssd1 vccd1 vccd1 input59/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17454__S _17488_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16850_ _16849_/X _13868_/Y _17545_/S vssd1 vssd1 vccd1 vccd1 _16850_/X sky130_fd_sc_hd__mux2_1
X_15801_ _18242_/Q _16096_/B vssd1 vssd1 vccd1 vccd1 _15801_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__19358__RESET_B hold370/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16781_ _16780_/X _20033_/Q _17414_/S vssd1 vssd1 vccd1 vccd1 _16781_/X sky130_fd_sc_hd__mux2_1
XFILLER_77_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13993_ _18681_/Q vssd1 vssd1 vccd1 vccd1 _14012_/B sky130_fd_sc_hd__inv_2
X_18520_ _19814_/CLK _18520_/D repeater223/X vssd1 vssd1 vccd1 vccd1 _18520_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_207_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15732_ _20037_/Q vssd1 vssd1 vccd1 vccd1 _15732_/Y sky130_fd_sc_hd__clkinv_4
X_12944_ _19274_/Q _12965_/C _12942_/Y _18931_/Q _12943_/X vssd1 vssd1 vccd1 vccd1
+ _12944_/X sky130_fd_sc_hd__a221o_1
XANTENNA__10700__A _18879_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18451_ _18460_/CLK _18451_/D vssd1 vssd1 vccd1 vccd1 _18451_/Q sky130_fd_sc_hd__dfxtp_1
X_15663_ _15666_/A _15663_/B vssd1 vssd1 vccd1 vccd1 _15663_/Y sky130_fd_sc_hd__nor2_1
XFILLER_45_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12875_ _12964_/C _12875_/B vssd1 vssd1 vccd1 vccd1 _12994_/A sky130_fd_sc_hd__or2_1
XFILLER_34_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17402_ _17401_/X _10200_/Y _17566_/S vssd1 vssd1 vccd1 vccd1 _17402_/X sky130_fd_sc_hd__mux2_1
XPHY_4272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14614_ _18763_/Q _14628_/B _15195_/B vssd1 vssd1 vccd1 vccd1 _15145_/C sky130_fd_sc_hd__or3_4
XPHY_4283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18382_ _18441_/CLK _18382_/D vssd1 vssd1 vccd1 vccd1 _18382_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12605__B1 _12536_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11826_ _19442_/Q _11821_/X _10863_/X _11822_/X vssd1 vssd1 vccd1 vccd1 _19442_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15594_ _15594_/A _15594_/B vssd1 vssd1 vccd1 vccd1 _15594_/Y sky130_fd_sc_hd__nor2_1
XPHY_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17333_ _15768_/Y _14195_/Y _17546_/S vssd1 vssd1 vccd1 vccd1 _17333_/X sky130_fd_sc_hd__mux2_1
XFILLER_230_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14545_ _14598_/A _14545_/B _14598_/C vssd1 vssd1 vccd1 vccd1 _14547_/A sky130_fd_sc_hd__or3_4
XPHY_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11757_ _11771_/A vssd1 vssd1 vccd1 vccd1 _11757_/X sky130_fd_sc_hd__clkbuf_2
XPHY_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10708_ hold336/X vssd1 vssd1 vccd1 vccd1 _10708_/Y sky130_fd_sc_hd__inv_2
X_17264_ _15963_/X _09541_/Y _17534_/S vssd1 vssd1 vccd1 vccd1 _17264_/X sky130_fd_sc_hd__mux2_1
XPHY_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14476_ _14476_/A _15318_/B vssd1 vssd1 vccd1 vccd1 _15009_/C sky130_fd_sc_hd__or2_2
X_11688_ _11671_/X _11672_/Y _18628_/Q _19529_/Q _11668_/X vssd1 vssd1 vccd1 vccd1
+ _19529_/D sky130_fd_sc_hd__a32o_1
XFILLER_201_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19003_ _19208_/CLK _19003_/D hold363/X vssd1 vssd1 vccd1 vccd1 _19003_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_128_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16215_ _16215_/A _16469_/B vssd1 vssd1 vccd1 vccd1 _16215_/Y sky130_fd_sc_hd__nor2_1
X_13427_ _18866_/Q _13435_/A _13426_/X _13354_/B vssd1 vssd1 vccd1 vccd1 _18866_/D
+ sky130_fd_sc_hd__o211a_1
X_10639_ _10638_/Y _10598_/A _10617_/X _10589_/B _10618_/A vssd1 vssd1 vccd1 vccd1
+ _10640_/A sky130_fd_sc_hd__o32a_1
X_17195_ _17194_/X _11317_/Y _17459_/S vssd1 vssd1 vccd1 vccd1 _17195_/X sky130_fd_sc_hd__mux2_1
XFILLER_143_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16146_ _17426_/X _15904_/A _17433_/X _15999_/X vssd1 vssd1 vccd1 vccd1 _16146_/X
+ sky130_fd_sc_hd__o22a_1
X_13358_ _20102_/Q vssd1 vssd1 vccd1 vccd1 _13358_/Y sky130_fd_sc_hd__inv_2
XFILLER_182_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12309_ _12309_/A _12316_/B vssd1 vssd1 vccd1 vccd1 _12310_/S sky130_fd_sc_hd__or2_1
X_16077_ _15846_/X _16058_/X _15859_/X _16065_/X _16076_/X vssd1 vssd1 vccd1 vccd1
+ _16077_/Y sky130_fd_sc_hd__o221ai_4
X_13289_ _18869_/Q vssd1 vssd1 vccd1 vccd1 _13289_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19905_ _19905_/CLK _19905_/D repeater191/X vssd1 vssd1 vccd1 vccd1 _19905_/Q sky130_fd_sc_hd__dfrtp_1
X_15028_ _18039_/Q _15023_/X _14998_/X _15025_/X vssd1 vssd1 vccd1 vccd1 _18039_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_170_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17364__S _17544_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19836_ _20058_/CLK _19836_/D repeater271/X vssd1 vssd1 vccd1 vccd1 _19836_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_96_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16488__B _17567_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19099__RESET_B repeater252/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19767_ _19771_/CLK _19767_/D repeater189/X vssd1 vssd1 vccd1 vccd1 _19767_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_37_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput3 input3/A vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_1
X_16979_ _16473_/Y _15477_/Y _17524_/S vssd1 vssd1 vccd1 vccd1 _16979_/X sky130_fd_sc_hd__mux2_1
X_09520_ _09494_/A _19324_/Q _20034_/Q _09517_/Y _09519_/X vssd1 vssd1 vccd1 vccd1
+ _09528_/B sky130_fd_sc_hd__o221a_1
XANTENNA__19028__RESET_B repeater269/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_237_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18718_ _18718_/CLK _18718_/D repeater253/X vssd1 vssd1 vccd1 vccd1 _18718_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_232_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19698_ _19720_/CLK _19698_/D repeater201/X vssd1 vssd1 vccd1 vccd1 _19698_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_36_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19944__CLK _19976_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09451_ _19907_/Q _09446_/Y _10083_/A _19371_/Q _09450_/X vssd1 vssd1 vccd1 vccd1
+ _09463_/B sky130_fd_sc_hd__o221a_1
XFILLER_225_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18649_ _20050_/CLK _18649_/D repeater197/X vssd1 vssd1 vccd1 vccd1 _18649_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_240_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14597__B1 hold320/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09382_ _19910_/Q vssd1 vssd1 vccd1 vccd1 _10082_/A sky130_fd_sc_hd__inv_2
XFILLER_224_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17539__S _17539_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14521__B1 _14437_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09284__C _11742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17274__S _17490_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19451__RESET_B repeater271/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_1_0_HCLK_A clkbuf_3_1_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14199__A _19119_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09718_ _09742_/A _19415_/Q _09742_/A _19415_/Q vssd1 vssd1 vccd1 vccd1 _09718_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_10990_ _10984_/B _10978_/X _10988_/Y _10989_/X _10963_/A vssd1 vssd1 vccd1 vccd1
+ _10991_/A sky130_fd_sc_hd__o32a_1
XFILLER_71_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09649_ _19986_/Q vssd1 vssd1 vccd1 vccd1 _09742_/A sky130_fd_sc_hd__inv_2
XFILLER_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12660_ _12698_/A vssd1 vssd1 vccd1 vccd1 _12677_/A sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_248_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11611_ _11575_/A _11575_/B _11617_/A _11609_/Y vssd1 vssd1 vccd1 vccd1 _19562_/D
+ sky130_fd_sc_hd__a211oi_2
XPHY_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12591_ _12600_/A vssd1 vssd1 vccd1 vccd1 _12591_/X sky130_fd_sc_hd__clkbuf_2
XPHY_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14330_ _18436_/Q _14319_/A _14329_/X _14320_/A vssd1 vssd1 vccd1 vccd1 _18436_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11542_ _19579_/Q _11541_/Y _11504_/A _11542_/C1 vssd1 vssd1 vccd1 vccd1 _19579_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17449__S _17534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14261_ _18473_/Q _14258_/X _12714_/X _14260_/X vssd1 vssd1 vccd1 vccd1 _18473_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_156_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11473_ _11473_/A _11517_/A vssd1 vssd1 vccd1 vccd1 _11474_/B sky130_fd_sc_hd__or2_1
XPHY_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16000_ _17494_/X _15904_/A _17503_/X _15999_/X vssd1 vssd1 vccd1 vccd1 _16000_/X
+ sky130_fd_sc_hd__o22a_1
X_13212_ _13062_/A _13212_/A2 _13210_/Y _13202_/X vssd1 vssd1 vccd1 vccd1 _18889_/D
+ sky130_fd_sc_hd__a211oi_2
X_10424_ _19844_/Q _10417_/X _10423_/X _10419_/Y vssd1 vssd1 vccd1 vccd1 _19844_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_109_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14192_ _19096_/Q _14006_/A _14191_/Y _18681_/Q vssd1 vssd1 vccd1 vccd1 _14192_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_164_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17924__S1 _19648_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13143_ _19168_/Q _13069_/A _16210_/A _18891_/Q _13142_/X vssd1 vssd1 vccd1 vccd1
+ _13144_/D sky130_fd_sc_hd__o221a_1
X_10355_ _10349_/B _10320_/X _10353_/Y _10354_/X _10328_/A vssd1 vssd1 vccd1 vccd1
+ _10356_/A sky130_fd_sc_hd__o32a_1
XANTENNA__19539__RESET_B repeater221/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14512__B1 hold330/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17951_ _20079_/CLK _17951_/D vssd1 vssd1 vccd1 vccd1 _17951_/Q sky130_fd_sc_hd__dfxtp_1
X_13074_ _13074_/A _13190_/A vssd1 vssd1 vccd1 vccd1 _13075_/B sky130_fd_sc_hd__or2_2
X_10286_ _10286_/A _10286_/B vssd1 vssd1 vccd1 vccd1 _19872_/D sky130_fd_sc_hd__or2_1
XANTENNA__17184__S _17545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16902_ _16469_/Y _20099_/Q _17385_/S vssd1 vssd1 vccd1 vccd1 _16902_/X sky130_fd_sc_hd__mux2_1
X_12025_ _19347_/Q _12023_/X hold276/X _12024_/X vssd1 vssd1 vccd1 vccd1 _19347_/D
+ sky130_fd_sc_hd__a22o_1
X_17882_ _16086_/Y _16087_/Y _16088_/Y _16089_/Y _17913_/S0 _19632_/Q vssd1 vssd1
+ vccd1 vccd1 _17882_/X sky130_fd_sc_hd__mux4_1
XFILLER_239_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19621_ _19920_/CLK _19621_/D repeater229/X vssd1 vssd1 vccd1 vccd1 _19621_/Q sky130_fd_sc_hd__dfrtp_1
X_16833_ _16832_/X _13357_/Y _17385_/S vssd1 vssd1 vccd1 vccd1 _16833_/X sky130_fd_sc_hd__mux2_1
XFILLER_38_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16764_ _16763_/X _13391_/Y _17535_/S vssd1 vssd1 vccd1 vccd1 _16764_/X sky130_fd_sc_hd__mux2_1
X_19552_ _19561_/CLK _19552_/D hold348/A vssd1 vssd1 vccd1 vccd1 _19552_/Q sky130_fd_sc_hd__dfrtp_1
X_13976_ _18698_/Q vssd1 vssd1 vccd1 vccd1 _14028_/A sky130_fd_sc_hd__inv_2
XFILLER_207_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20097__RESET_B repeater233/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18503_ _19795_/CLK _18503_/D repeater226/X vssd1 vssd1 vccd1 vccd1 _18503_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_34_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15715_ _15715_/A _15715_/B vssd1 vssd1 vccd1 vccd1 _18650_/D sky130_fd_sc_hd__nor2_1
XFILLER_207_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12927_ _19284_/Q _12967_/B _19282_/Q _12964_/B vssd1 vssd1 vccd1 vccd1 _12927_/X
+ sky130_fd_sc_hd__o22a_1
X_19483_ _19506_/CLK hold176/X repeater260/X vssd1 vssd1 vccd1 vccd1 _19483_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_61_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16695_ _17095_/X _16683_/X _17079_/X _16684_/X _16694_/X vssd1 vssd1 vccd1 vccd1
+ _16698_/B sky130_fd_sc_hd__o221a_4
XANTENNA__20026__RESET_B repeater239/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18434_ _18795_/CLK _18434_/D vssd1 vssd1 vccd1 vccd1 _18434_/Q sky130_fd_sc_hd__dfxtp_1
X_15646_ _18605_/Q _15649_/C _15645_/Y _15641_/Y vssd1 vssd1 vccd1 vccd1 _15647_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__17860__S0 _17913_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12858_ _18920_/Q vssd1 vssd1 vccd1 vccd1 _13021_/C sky130_fd_sc_hd__inv_2
XPHY_4080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12054__A1 _17614_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18365_ _19515_/CLK _18365_/D vssd1 vssd1 vccd1 vccd1 _18365_/Q sky130_fd_sc_hd__dfxtp_1
X_11809_ _19455_/Q _11807_/X hold276/X _11808_/X vssd1 vssd1 vccd1 vccd1 _19455_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13251__B1 _12543_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15577_ _15610_/A _18588_/Q vssd1 vssd1 vccd1 vccd1 _15577_/Y sky130_fd_sc_hd__nor2_1
X_12789_ _19248_/Q _13548_/A _19244_/Q _13544_/A _12788_/X vssd1 vssd1 vccd1 vccd1
+ _12808_/A sky130_fd_sc_hd__o221a_1
XPHY_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17316_ _16414_/X _18233_/Q _17564_/S vssd1 vssd1 vccd1 vccd1 _17316_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14528_ _18322_/Q _14519_/A _14474_/X _14520_/A vssd1 vssd1 vccd1 vccd1 _18322_/D
+ sky130_fd_sc_hd__a22o_1
X_18296_ _18435_/CLK _18296_/D vssd1 vssd1 vccd1 vccd1 _18296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17359__S _17386_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17247_ _17246_/X _19956_/Q _17518_/S vssd1 vssd1 vccd1 vccd1 _17247_/X sky130_fd_sc_hd__mux2_1
XFILLER_175_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14459_ _18364_/Q _14452_/A _14419_/X _14453_/A vssd1 vssd1 vccd1 vccd1 _18364_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16740__B2 _15896_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17178_ _17177_/X _13072_/A _17542_/S vssd1 vssd1 vccd1 vccd1 _17178_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16129_ _16127_/Y _15973_/A _16128_/Y _16055_/X vssd1 vssd1 vccd1 vccd1 _16129_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__17915__S1 _18750_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19962__RESET_B hold371/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12092__A hold298/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08981__A1 _18870_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08951_ _19865_/Q vssd1 vssd1 vccd1 vccd1 _10331_/A sky130_fd_sc_hd__inv_2
XFILLER_102_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17094__S _17490_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19819_ _19822_/CLK _19819_/D repeater228/X vssd1 vssd1 vccd1 vccd1 _19819_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_244_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09503_ _20022_/Q _09500_/Y _09487_/A _19317_/Q _09502_/X vssd1 vssd1 vccd1 vccd1
+ _09512_/B sky130_fd_sc_hd__o221a_1
XFILLER_213_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09434_ _10013_/A _19366_/Q _19906_/Q _09430_/Y _09433_/X vssd1 vssd1 vccd1 vccd1
+ _09440_/C sky130_fd_sc_hd__o221a_1
XFILLER_24_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18844__RESET_B repeater232/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_212_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17851__S0 _17913_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09365_ _20012_/Q vssd1 vssd1 vccd1 vccd1 _09473_/A sky130_fd_sc_hd__inv_4
XANTENNA__11171__A _19814_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09296_ _20043_/Q _09293_/X _09098_/X _09294_/X vssd1 vssd1 vccd1 vccd1 _20043_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_177_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17269__S _17542_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15578__A _15610_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16731__B2 _16512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14742__B1 _14693_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17906__S1 _18759_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13098__A _19172_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16901__S _17513_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18864__CLK _18866_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10140_ _16985_/X _10136_/X _19902_/Q _10138_/X vssd1 vssd1 vccd1 vccd1 _19902_/D
+ sky130_fd_sc_hd__o22a_1
XANTENNA__19632__RESET_B repeater258/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10071_ _10071_/A vssd1 vssd1 vccd1 vccd1 _10071_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_198_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17732__S _18508_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13830_ _13830_/A _13830_/B _13917_/A vssd1 vssd1 vccd1 vccd1 _13906_/A sky130_fd_sc_hd__or3_1
XANTENNA__10250__A _19516_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_216_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13761_ _13756_/A _13756_/B _13757_/A _13760_/X vssd1 vssd1 vccd1 vccd1 _13761_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_44_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10973_ _10973_/A _10973_/B vssd1 vssd1 vccd1 vccd1 _10973_/Y sky130_fd_sc_hd__nor2_1
XFILLER_204_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15500_ _15498_/Y _15499_/X _15483_/X vssd1 vssd1 vccd1 vccd1 _15500_/X sky130_fd_sc_hd__o21a_1
XFILLER_16_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18244__CLK _19847_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12712_ _14802_/A _12709_/X hold242/X _12711_/X vssd1 vssd1 vccd1 vccd1 _18959_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17842__S0 _17913_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18585__RESET_B repeater272/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16480_ _16979_/X _16638_/A _16990_/X _16688_/A _16479_/Y vssd1 vssd1 vccd1 vccd1
+ _16481_/C sky130_fd_sc_hd__o221a_1
XFILLER_189_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13692_ _15197_/A vssd1 vssd1 vccd1 vccd1 _16435_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_16_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15431_ _19622_/Q _11167_/B _11168_/B vssd1 vssd1 vccd1 vccd1 _15431_/X sky130_fd_sc_hd__a21bo_1
XFILLER_62_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18514__RESET_B repeater208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12643_ _12650_/A vssd1 vssd1 vccd1 vccd1 _12643_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_30_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18150_ _18165_/CLK _18150_/D vssd1 vssd1 vccd1 vccd1 _18150_/Q sky130_fd_sc_hd__dfxtp_1
X_15362_ _15364_/A _17588_/X vssd1 vssd1 vccd1 vccd1 _18502_/D sky130_fd_sc_hd__and2_1
XPHY_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12574_ _19048_/Q _12569_/X _12396_/X _12570_/X vssd1 vssd1 vccd1 vccd1 _19048_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17101_ _17100_/X _09472_/A _17530_/S vssd1 vssd1 vccd1 vccd1 _17101_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11795__B1 _09030_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14313_ _18443_/Q _14304_/A _14312_/X _14305_/A vssd1 vssd1 vccd1 vccd1 _18443_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17179__S _17543_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11525_ _11525_/A vssd1 vssd1 vccd1 vccd1 _11528_/B sky130_fd_sc_hd__inv_2
XPHY_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18081_ _18137_/CLK _18081_/D vssd1 vssd1 vccd1 vccd1 _18081_/Q sky130_fd_sc_hd__dfxtp_1
X_15293_ _15388_/A _15292_/X _10612_/Y _15277_/Y _15220_/Y vssd1 vssd1 vccd1 vccd1
+ _18553_/D sky130_fd_sc_hd__o221ai_1
XFILLER_157_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17032_ _17031_/X _15557_/A _17474_/S vssd1 vssd1 vccd1 vccd1 _17032_/X sky130_fd_sc_hd__mux2_1
X_14244_ _18554_/Q _15334_/A _18664_/Q _18508_/Q vssd1 vssd1 vccd1 vccd1 _18664_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_7_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11456_ _11437_/X _11456_/B _11456_/C _11456_/D vssd1 vssd1 vccd1 vccd1 _11457_/D
+ sky130_fd_sc_hd__and4b_1
X_10407_ _19847_/Q vssd1 vssd1 vccd1 vccd1 _10989_/A sky130_fd_sc_hd__clkbuf_2
X_14175_ _19123_/Q _14032_/A _14171_/Y _18673_/Q _14174_/X vssd1 vssd1 vccd1 vccd1
+ _14184_/B sky130_fd_sc_hd__o221a_1
X_11387_ _11581_/A _19148_/Q _19567_/Q _11386_/Y vssd1 vssd1 vccd1 vccd1 _11387_/X
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__16811__S _17490_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13126_ _13122_/Y _18905_/Q _19164_/Q _13066_/A _13125_/X vssd1 vssd1 vccd1 vccd1
+ _13127_/D sky130_fd_sc_hd__o221a_1
X_10338_ _10338_/A vssd1 vssd1 vccd1 vccd1 _19867_/D sky130_fd_sc_hd__inv_2
X_18983_ _19600_/CLK _18983_/D hold273/X vssd1 vssd1 vccd1 vccd1 _18983_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_112_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17934_ _18465_/CLK _17934_/D vssd1 vssd1 vccd1 vccd1 _17934_/Q sky130_fd_sc_hd__dfxtp_1
X_13057_ _18889_/Q vssd1 vssd1 vccd1 vccd1 _13062_/A sky130_fd_sc_hd__inv_2
XFILLER_112_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10269_ _10263_/X _10268_/B _10267_/Y _19648_/Q _11039_/B vssd1 vssd1 vccd1 vccd1
+ _10269_/X sky130_fd_sc_hd__a32o_1
XFILLER_79_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12008_ _19358_/Q _12000_/X _09027_/X _12003_/X vssd1 vssd1 vccd1 vccd1 _19358_/D
+ sky130_fd_sc_hd__a22o_1
X_17865_ _16177_/Y _16178_/Y _16179_/Y _16180_/Y _17908_/S0 _18759_/Q vssd1 vssd1
+ vccd1 vccd1 _17865_/X sky130_fd_sc_hd__mux4_2
XANTENNA__16789__A1 _18989_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17642__S _17655_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19604_ _19610_/CLK _19604_/D hold343/X vssd1 vssd1 vccd1 vccd1 _19604_/Q sky130_fd_sc_hd__dfrtp_1
X_16816_ _15963_/X _12777_/Y _17534_/S vssd1 vssd1 vccd1 vccd1 _16816_/X sky130_fd_sc_hd__mux2_1
XFILLER_213_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17796_ _18392_/Q _18384_/Q _18376_/Q _18368_/Q _17923_/S0 _19646_/Q vssd1 vssd1
+ vccd1 vccd1 _17796_/X sky130_fd_sc_hd__mux4_2
XFILLER_35_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19535_ _19541_/CLK _19535_/D repeater221/X vssd1 vssd1 vccd1 vccd1 _19535_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_19_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16747_ _16747_/A _16747_/B vssd1 vssd1 vccd1 vccd1 _16747_/Y sky130_fd_sc_hd__nor2_8
X_13959_ _13947_/A _13947_/B _13957_/Y _13919_/X vssd1 vssd1 vccd1 vccd1 _18710_/D
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__14567__A _14780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16678_ _16678_/A _16678_/B _16678_/C _16678_/D vssd1 vssd1 vccd1 vccd1 _16678_/X
+ sky130_fd_sc_hd__or4_4
XANTENNA__17833__S0 _17918_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19466_ _19970_/CLK _19466_/D repeater274/X vssd1 vssd1 vccd1 vccd1 _19466_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_222_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18417_ _19849_/CLK _18417_/D vssd1 vssd1 vccd1 vccd1 _18417_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15629_ _15629_/A vssd1 vssd1 vccd1 vccd1 _15629_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18737__CLK _20051_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19397_ _20091_/CLK _19397_/D repeater236/X vssd1 vssd1 vccd1 vccd1 _19397_/Q sky130_fd_sc_hd__dfrtp_1
X_09150_ _09154_/A _09156_/A _09144_/C _20087_/Q _09138_/A vssd1 vssd1 vccd1 vccd1
+ _09151_/B sky130_fd_sc_hd__o32a_1
XANTENNA__09979__B1 _09968_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18348_ _19630_/CLK _18348_/D vssd1 vssd1 vccd1 vccd1 _18348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10319__B _13285_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17089__S _17548_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18279_ _19847_/CLK _18279_/D vssd1 vssd1 vccd1 vccd1 _18279_/Q sky130_fd_sc_hd__dfxtp_1
X_09081_ hold248/X vssd1 vssd1 vccd1 vccd1 _10446_/A sky130_fd_sc_hd__buf_4
XFILLER_163_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16713__B2 _16002_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13527__A1 _13491_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_238_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput50 input50/A vssd1 vssd1 vccd1 vccd1 input50/X sky130_fd_sc_hd__clkbuf_4
Xinput61 input61/A vssd1 vssd1 vccd1 vccd1 input61/X sky130_fd_sc_hd__buf_4
Xinput72 input72/A vssd1 vssd1 vccd1 vccd1 input72/X sky130_fd_sc_hd__buf_2
XFILLER_238_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15845__B _15858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09983_ _09859_/A _09983_/A2 _09981_/Y _09970_/X vssd1 vssd1 vccd1 vccd1 _19951_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_115_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08934_ _18782_/Q vssd1 vssd1 vccd1 vccd1 _08934_/Y sky130_fd_sc_hd__inv_2
XFILLER_69_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17552__S _19498_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12266__A1 _19222_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17824__S0 _18751_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09417_ _09397_/X _09400_/X _09417_/C _09417_/D vssd1 vssd1 vccd1 vccd1 _09417_/Y
+ sky130_fd_sc_hd__nand4bb_2
XFILLER_25_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_198_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_240_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09348_ _20029_/Q vssd1 vssd1 vccd1 vccd1 _09489_/A sky130_fd_sc_hd__inv_2
XFILLER_200_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09279_ _20050_/Q _09270_/A _09108_/X _09271_/A vssd1 vssd1 vccd1 vccd1 _20050_/D
+ sky130_fd_sc_hd__a22o_1
X_11310_ _11227_/Y _18991_/Q _19587_/Q _11308_/Y _11309_/X vssd1 vssd1 vccd1 vccd1
+ _11315_/C sky130_fd_sc_hd__o221a_1
XFILLER_148_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12290_ _12298_/A vssd1 vssd1 vccd1 vccd1 _12290_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_113_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11241_ _19579_/Q _11236_/Y _11464_/A _18997_/Q _11240_/X vssd1 vssd1 vccd1 vccd1
+ _11248_/C sky130_fd_sc_hd__o221a_1
XFILLER_180_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11172_ _18526_/Q vssd1 vssd1 vccd1 vccd1 _11173_/C sky130_fd_sc_hd__inv_2
XFILLER_134_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10123_ _18577_/Q _18576_/Q _18578_/Q vssd1 vssd1 vccd1 vccd1 _15537_/A sky130_fd_sc_hd__or3_1
XANTENNA__15140__B1 _10698_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15980_ _19522_/Q vssd1 vssd1 vccd1 vccd1 _15980_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10054_ _19934_/Q _10052_/X _10053_/X _10049_/A vssd1 vssd1 vccd1 vccd1 _19934_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA_input33_A HREADY vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14931_ _20077_/Q vssd1 vssd1 vccd1 vccd1 _14931_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_leaf_125_HCLK_A clkbuf_4_4_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17462__S _19498_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15771__A _16721_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17650_ _15634_/Y _19039_/Q _17655_/S vssd1 vssd1 vccd1 vccd1 _18602_/D sky130_fd_sc_hd__mux2_1
X_14862_ _18136_/Q _14858_/X _14703_/X _14860_/X vssd1 vssd1 vccd1 vccd1 _18136_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_208_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_236_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16586__B _16615_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16601_ _19457_/Q vssd1 vssd1 vccd1 vccd1 _16601_/Y sky130_fd_sc_hd__inv_2
X_13813_ _13945_/A _13944_/C _13813_/C _13813_/D vssd1 vssd1 vccd1 vccd1 _13912_/A
+ sky130_fd_sc_hd__or4_4
X_17581_ _15397_/X _19526_/Q _17584_/S vssd1 vssd1 vccd1 vccd1 _17581_/X sky130_fd_sc_hd__mux2_1
XFILLER_91_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14793_ _14793_/A vssd1 vssd1 vccd1 vccd1 _14793_/X sky130_fd_sc_hd__buf_2
XFILLER_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19320_ _19320_/CLK _19320_/D repeater214/X vssd1 vssd1 vccd1 vccd1 _19320_/Q sky130_fd_sc_hd__dfrtp_4
X_16532_ _17161_/X _16512_/X _17149_/X _16513_/X _16531_/X vssd1 vssd1 vccd1 vccd1
+ _16532_/X sky130_fd_sc_hd__o221a_4
XANTENNA__17815__S0 _17918_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13744_ _13737_/A _13259_/B _17764_/X _18749_/Q vssd1 vssd1 vccd1 vccd1 _18749_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_204_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_188_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10956_ _10956_/A _10956_/B _10956_/C _10956_/D vssd1 vssd1 vccd1 vccd1 _11009_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_73_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19251_ _19324_/CLK _19251_/D repeater237/X vssd1 vssd1 vccd1 vccd1 _19251_/Q sky130_fd_sc_hd__dfrtp_4
X_16463_ _17081_/X _16148_/X _16768_/X _16394_/X vssd1 vssd1 vccd1 vccd1 _16463_/X
+ sky130_fd_sc_hd__o22a_1
X_13675_ _18776_/Q _13671_/X _13674_/X _13672_/X vssd1 vssd1 vccd1 vccd1 _18776_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_232_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10887_ _19697_/Q _10875_/X _10861_/X _10879_/X vssd1 vssd1 vccd1 vccd1 _19697_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16806__S _17488_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater172_A _17488_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15414_ _18539_/Q _13226_/B _13227_/B vssd1 vssd1 vccd1 vccd1 _15414_/X sky130_fd_sc_hd__a21bo_1
X_18202_ _18460_/CLK _18202_/D vssd1 vssd1 vccd1 vccd1 _18202_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12626_ _19016_/Q _12622_/X _12394_/X _12623_/X vssd1 vssd1 vccd1 vccd1 _19016_/D
+ sky130_fd_sc_hd__a22o_1
X_19182_ _19293_/CLK _19182_/D repeater187/X vssd1 vssd1 vccd1 vccd1 _19182_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16394_ _16633_/A vssd1 vssd1 vccd1 vccd1 _16394_/X sky130_fd_sc_hd__clkbuf_4
XPHY_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18133_ _18137_/CLK _18133_/D vssd1 vssd1 vccd1 vccd1 _18133_/Q sky130_fd_sc_hd__dfxtp_1
X_15345_ _15347_/A _17596_/X vssd1 vssd1 vccd1 vccd1 _18494_/D sky130_fd_sc_hd__and2_1
X_12557_ _12553_/A _12556_/B _19057_/Q _12556_/Y vssd1 vssd1 vccd1 vccd1 _19057_/D
+ sky130_fd_sc_hd__o22a_1
XPHY_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11508_ _11508_/A vssd1 vssd1 vccd1 vccd1 _11508_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19554__RESET_B hold348/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18064_ _18465_/CLK _18064_/D vssd1 vssd1 vccd1 vccd1 _18064_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10440__B1 _09071_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15276_ _15278_/B _15275_/A _15215_/B _15275_/Y _10933_/A vssd1 vssd1 vccd1 vccd1
+ _15276_/X sky130_fd_sc_hd__o221a_1
XFILLER_144_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12488_ _12528_/A vssd1 vssd1 vccd1 vccd1 _12505_/A sky130_fd_sc_hd__clkbuf_2
X_17015_ _15768_/Y _14180_/Y _17546_/S vssd1 vssd1 vccd1 vccd1 _17015_/X sky130_fd_sc_hd__mux2_1
X_14227_ _18497_/Q _14227_/B vssd1 vssd1 vccd1 vccd1 _14228_/B sky130_fd_sc_hd__or2_1
XANTENNA__17637__S _17655_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11439_ _19144_/Q vssd1 vssd1 vccd1 vccd1 _11439_/Y sky130_fd_sc_hd__inv_2
XFILLER_160_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10155__A _10155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12193__B1 _12069_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14158_ _19095_/Q _14005_/A _14155_/Y _18679_/Q _14157_/X vssd1 vssd1 vccd1 vccd1
+ _14166_/B sky130_fd_sc_hd__o221a_1
XFILLER_152_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13109_ _13109_/A _13109_/B _13109_/C _13109_/D vssd1 vssd1 vccd1 vccd1 _13160_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_140_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14089_ _14050_/Y _18678_/Q _14087_/Y _18688_/Q _14088_/X vssd1 vssd1 vccd1 vccd1
+ _14093_/C sky130_fd_sc_hd__o221a_1
X_18966_ _19137_/CLK _18966_/D hold370/X vssd1 vssd1 vccd1 vccd1 _18966_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12370__A _12370_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17917_ _18361_/Q _18001_/Q _18417_/Q _18401_/Q _17918_/S0 _18750_/Q vssd1 vssd1
+ vccd1 vccd1 _17917_/X sky130_fd_sc_hd__mux4_2
XFILLER_140_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18897_ _18908_/CLK _18897_/D hold373/X vssd1 vssd1 vccd1 vccd1 _18897_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_121_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17372__S _17567_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17848_ _16359_/Y _16360_/Y _16361_/Y _16362_/Y _17908_/S0 _18759_/Q vssd1 vssd1
+ vccd1 vccd1 _17848_/X sky130_fd_sc_hd__mux4_1
XFILLER_27_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_226_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17779_ _17775_/X _17776_/X _17777_/X _17778_/X _19647_/Q _19648_/Q vssd1 vssd1 vccd1
+ vccd1 _17779_/X sky130_fd_sc_hd__mux4_2
XANTENNA_clkbuf_leaf_47_HCLK_A clkbuf_opt_2_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_241_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19518_ _19867_/CLK hold205/X repeater262/X vssd1 vssd1 vccd1 vccd1 _19518_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_240_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17806__S0 _17918_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19449_ _20058_/CLK _19449_/D repeater271/X vssd1 vssd1 vccd1 vccd1 _19449_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_195_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09202_ _09202_/A vssd1 vssd1 vccd1 vccd1 _20070_/D sky130_fd_sc_hd__inv_2
XFILLER_10_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09133_ _15321_/A _09138_/A _09133_/C vssd1 vssd1 vccd1 vccd1 _09133_/X sky130_fd_sc_hd__and3_1
XANTENNA__19295__RESET_B repeater239/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09064_ _12030_/A vssd1 vssd1 vccd1 vccd1 _09064_/X sky130_fd_sc_hd__buf_4
XFILLER_135_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17547__S _17547_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09966_ _09869_/A _09869_/B _09963_/Y _09987_/B vssd1 vssd1 vccd1 vccd1 _19961_/D
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__16870__A0 _15963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08917_ _08917_/A vssd1 vssd1 vccd1 vccd1 _16986_/S sky130_fd_sc_hd__clkinv_4
X_20086_ _20124_/CLK _20086_/D repeater205/X vssd1 vssd1 vccd1 vccd1 _20086_/Q sky130_fd_sc_hd__dfrtp_1
X_09897_ _19344_/Q vssd1 vssd1 vccd1 vccd1 _09897_/Y sky130_fd_sc_hd__inv_2
XFILLER_245_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16687__A _16687_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17282__S _17386_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_4_15_0_HCLK_A clkbuf_3_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold265_A HWDATA[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10810_ _10810_/A vssd1 vssd1 vccd1 vccd1 _10810_/X sky130_fd_sc_hd__clkbuf_2
XPHY_3912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11790_ _19468_/Q _11784_/X hold288/X _11787_/X vssd1 vssd1 vccd1 vccd1 _19468_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12439__B _12487_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10741_ _10742_/A vssd1 vssd1 vccd1 vccd1 _10741_/X sky130_fd_sc_hd__clkbuf_2
XPHY_3967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16925__A1 hold148/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_214_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13739__A1 _18752_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13460_ _18850_/Q _13459_/Y _13443_/A _13338_/B vssd1 vssd1 vccd1 vccd1 _18850_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_198_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10672_ _17735_/X _10669_/X _19790_/Q _10670_/X vssd1 vssd1 vccd1 vccd1 _19790_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14654__B _15839_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12411_ _19143_/Q _12400_/X _12410_/X _12402_/X vssd1 vssd1 vccd1 vccd1 _19143_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19408__CLK _19984_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13391_ _20117_/Q vssd1 vssd1 vccd1 vccd1 _13391_/Y sky130_fd_sc_hd__inv_1
XANTENNA__12411__A1 _19143_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10422__B1 _10421_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15130_ _17971_/Q _15123_/A _14933_/X _15124_/A vssd1 vssd1 vccd1 vccd1 _17971_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_126_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12342_ _12362_/A vssd1 vssd1 vccd1 vccd1 _12342_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_138_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_opt_2_HCLK clkbuf_opt_2_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_opt_2_HCLK/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_182_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15061_ _15061_/A vssd1 vssd1 vccd1 vccd1 _15061_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__17457__S _17545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12273_ _19217_/Q _12269_/X _12088_/X _12270_/X vssd1 vssd1 vccd1 vccd1 _19217_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_4_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12175__B1 _11918_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14012_ _14012_/A _14012_/B _14012_/C vssd1 vssd1 vccd1 vccd1 _14013_/B sky130_fd_sc_hd__or3_1
X_11224_ _18995_/Q vssd1 vssd1 vccd1 vccd1 _11224_/Y sky130_fd_sc_hd__inv_2
XANTENNA__09040__B1 _09039_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17102__A1 _18968_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10725__A1 _19770_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18820_ _18827_/CLK _18820_/D repeater231/X vssd1 vssd1 vccd1 vccd1 _18820_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12190__A _12228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11155_ _11155_/A vssd1 vssd1 vccd1 vccd1 _19627_/D sky130_fd_sc_hd__inv_2
XANTENNA__10703__A _18879_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10106_ _10101_/A _10101_/B _10101_/C vssd1 vssd1 vccd1 vccd1 _10107_/B sky130_fd_sc_hd__o21a_1
X_18751_ _19900_/CLK _18751_/D repeater195/X vssd1 vssd1 vccd1 vccd1 _18751_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_122_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11086_ _11086_/A _12246_/B vssd1 vssd1 vccd1 vccd1 _15232_/C sky130_fd_sc_hd__or2_1
X_15963_ _17539_/S _17537_/S _17548_/S _15881_/B vssd1 vssd1 vccd1 vccd1 _15963_/X
+ sky130_fd_sc_hd__or4b_4
XANTENNA__13675__B1 _13674_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16597__A _16597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17192__S _17493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17702_ _19816_/Q _19758_/Q _18548_/Q vssd1 vssd1 vccd1 vccd1 _17702_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10037_ _10037_/A _10074_/A vssd1 vssd1 vccd1 vccd1 _10038_/B sky130_fd_sc_hd__or2_2
X_14914_ _18102_/Q _14908_/X _14707_/X _14910_/X vssd1 vssd1 vccd1 vccd1 _18102_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_209_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18682_ _18686_/CLK _18682_/D repeater252/X vssd1 vssd1 vccd1 vccd1 _18682_/Q sky130_fd_sc_hd__dfrtp_4
X_15894_ _17518_/X _15887_/X _17524_/X _15889_/X _15893_/X vssd1 vssd1 vccd1 vccd1
+ _15918_/B sky130_fd_sc_hd__o221a_1
XFILLER_208_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17633_ _15705_/X _19056_/Q _17664_/S vssd1 vssd1 vccd1 vccd1 _18619_/D sky130_fd_sc_hd__mux2_1
XFILLER_208_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14845_ _14846_/A vssd1 vssd1 vccd1 vccd1 _14845_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_75_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17564_ _15801_/Y _15799_/Y _17564_/S vssd1 vssd1 vccd1 vccd1 _17564_/X sky130_fd_sc_hd__mux2_1
X_14776_ _18183_/Q _14771_/X _14751_/X _14773_/X vssd1 vssd1 vccd1 vccd1 _18183_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_210_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11988_ _12309_/A vssd1 vssd1 vccd1 vccd1 _15881_/B sky130_fd_sc_hd__buf_1
X_19303_ _20035_/CLK _19303_/D repeater242/X vssd1 vssd1 vccd1 vccd1 _19303_/Q sky130_fd_sc_hd__dfrtp_4
X_13727_ _13733_/A _13293_/X _14743_/A vssd1 vssd1 vccd1 vccd1 _13727_/X sky130_fd_sc_hd__o21a_1
X_16515_ _17266_/X _16512_/X _17304_/X _16513_/X _16514_/X vssd1 vssd1 vccd1 vccd1
+ _16515_/X sky130_fd_sc_hd__o221a_4
X_10939_ _19810_/Q _10939_/B _10939_/C _10939_/D vssd1 vssd1 vccd1 vccd1 _10940_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_90_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17495_ _15962_/X _20041_/Q _19498_/Q vssd1 vssd1 vccd1 vccd1 _17495_/X sky130_fd_sc_hd__mux2_1
XANTENNA__19735__RESET_B repeater208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19234_ _20035_/CLK _19234_/D repeater215/X vssd1 vssd1 vccd1 vccd1 _19234_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_189_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16446_ _16444_/Y _15830_/A _16445_/Y _15976_/X vssd1 vssd1 vccd1 vccd1 _16446_/X
+ sky130_fd_sc_hd__o22a_1
X_13658_ _13672_/A vssd1 vssd1 vccd1 vccd1 _13658_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_176_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12609_ _12659_/B _15863_/B vssd1 vssd1 vccd1 vccd1 _12610_/S sky130_fd_sc_hd__or2_1
X_16377_ _15227_/Y _15854_/A _16376_/Y _15976_/X vssd1 vssd1 vccd1 vccd1 _16377_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_31_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19165_ _19208_/CLK _19165_/D hold370/X vssd1 vssd1 vccd1 vccd1 _19165_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_129_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13589_ _13541_/A _13541_/B _13588_/X _13586_/Y vssd1 vssd1 vccd1 vccd1 _18818_/D
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__10413__A0 _10147_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15328_ _19699_/Q vssd1 vssd1 vccd1 vccd1 _15330_/A sky130_fd_sc_hd__inv_2
X_18116_ _19435_/CLK _18116_/D vssd1 vssd1 vccd1 vccd1 _18116_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19096_ _19585_/CLK _19096_/D hold365/X vssd1 vssd1 vccd1 vccd1 _19096_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17341__A1 _17849_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17367__S _17459_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15259_ _15259_/A _15259_/B vssd1 vssd1 vccd1 vccd1 _15259_/Y sky130_fd_sc_hd__nor2_1
XFILLER_145_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18047_ _18959_/CLK _18047_/D vssd1 vssd1 vccd1 vccd1 _18047_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14580__A _14793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12166__B1 _12035_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10716__A1 _19773_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11913__B1 _10877_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09820_ _19966_/Q vssd1 vssd1 vccd1 vccd1 _09874_/A sky130_fd_sc_hd__inv_2
XANTENNA__18688__RESET_B hold359/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19998_ _20003_/CLK _19998_/D repeater192/X vssd1 vssd1 vccd1 vccd1 _19998_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_99_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09751_ _09751_/A _09769_/A vssd1 vssd1 vccd1 vccd1 _09752_/B sky130_fd_sc_hd__or2_1
XANTENNA__18617__RESET_B repeater269/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18949_ _19290_/CLK _18949_/D repeater187/X vssd1 vssd1 vccd1 vccd1 _18949_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__13666__B1 hold250/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09682_ _19993_/Q _09681_/Y _09629_/B _19428_/Q vssd1 vssd1 vccd1 vccd1 _09682_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_39_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11444__A _19128_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_242_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09116_ _20086_/Q vssd1 vssd1 vccd1 vccd1 _15321_/B sky130_fd_sc_hd__inv_2
XFILLER_164_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17277__S _17566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15586__A _15610_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09047_ hold318/X vssd1 vssd1 vccd1 vccd1 hold317/A sky130_fd_sc_hd__buf_4
XFILLER_89_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15894__B2 _15889_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09022__B1 _09021_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17096__A0 _17486_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11904__B1 _09067_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19850__CLK _19851_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09949_ _09990_/A vssd1 vssd1 vccd1 vccd1 _09968_/A sky130_fd_sc_hd__inv_2
XFILLER_86_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12960_ _12960_/A vssd1 vssd1 vccd1 vccd1 _13027_/C sky130_fd_sc_hd__buf_6
X_20069_ _20070_/CLK _20069_/D repeater207/X vssd1 vssd1 vccd1 vccd1 _20069_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_180_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17399__A1 _17869_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_245_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11911_ hold260/X vssd1 vssd1 vccd1 vccd1 _11911_/X sky130_fd_sc_hd__clkbuf_4
X_12891_ _12891_/A _12891_/B vssd1 vssd1 vccd1 vccd1 _12892_/A sky130_fd_sc_hd__or2_1
XPHY_4410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17740__S _18508_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14630_ _14631_/A vssd1 vssd1 vccd1 vccd1 _14630_/X sky130_fd_sc_hd__clkbuf_2
XPHY_4443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10891__B1 _10870_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11842_ _15749_/A _11842_/B _15829_/B _11842_/D vssd1 vssd1 vccd1 vccd1 _14680_/B
+ sky130_fd_sc_hd__or4_4
XPHY_4454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14082__B1 _19081_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_30_HCLK_A _18641_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14561_ _18305_/Q _14558_/X _14531_/X _14560_/X vssd1 vssd1 vccd1 vccd1 _18305_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11773_ hold196/X _11771_/X _19475_/Q _11772_/X vssd1 vssd1 vccd1 vccd1 hold198/A
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12632__A1 _19012_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_93_HCLK_A clkbuf_4_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16300_ _19030_/Q vssd1 vssd1 vccd1 vccd1 _16300_/Y sky130_fd_sc_hd__inv_2
X_13512_ _18758_/Q vssd1 vssd1 vccd1 vccd1 _13704_/B sky130_fd_sc_hd__inv_2
XPHY_3786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10724_ _19771_/Q _10720_/X _10448_/X _10722_/X vssd1 vssd1 vccd1 vccd1 _19771_/D
+ sky130_fd_sc_hd__a22o_1
X_17280_ _15963_/X _12779_/Y _17534_/S vssd1 vssd1 vccd1 vccd1 _17280_/X sky130_fd_sc_hd__mux2_1
XFILLER_159_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14492_ _14492_/A vssd1 vssd1 vccd1 vccd1 _14493_/A sky130_fd_sc_hd__inv_2
XANTENNA__17571__A1 _19772_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16231_ _16229_/Y _16303_/A _16230_/Y _16055_/X vssd1 vssd1 vccd1 vccd1 _16231_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_70_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13443_ _13443_/A vssd1 vssd1 vccd1 vccd1 _13443_/X sky130_fd_sc_hd__clkbuf_2
X_10655_ _19795_/Q _10655_/B vssd1 vssd1 vccd1 vccd1 _10655_/X sky130_fd_sc_hd__or2_2
XANTENNA__12185__A _12187_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16162_ _18150_/Q vssd1 vssd1 vccd1 vccd1 _16162_/Y sky130_fd_sc_hd__inv_2
X_13374_ _20093_/Q vssd1 vssd1 vccd1 vccd1 _13374_/Y sky130_fd_sc_hd__inv_4
XFILLER_167_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10586_ _19800_/Q _19799_/Q _19813_/Q _10590_/D vssd1 vssd1 vccd1 vccd1 _10589_/C
+ sky130_fd_sc_hd__or4_4
X_15113_ _17984_/Q _15110_/X _14921_/X _15112_/X vssd1 vssd1 vccd1 vccd1 _17984_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17187__S _17545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12325_ _19186_/Q _12318_/X _12078_/X _12321_/X vssd1 vssd1 vccd1 vccd1 _19186_/D
+ sky130_fd_sc_hd__a22o_1
X_16093_ _18045_/Q vssd1 vssd1 vccd1 vccd1 _16093_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12148__B1 _12090_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19921_ _19927_/CLK _19921_/D repeater230/X vssd1 vssd1 vccd1 vccd1 _19921_/Q sky130_fd_sc_hd__dfrtp_1
X_15044_ _18027_/Q _15036_/A _15006_/X _15037_/A vssd1 vssd1 vccd1 vccd1 _18027_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_79_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12256_ _12370_/A _12370_/B _12256_/C vssd1 vssd1 vccd1 vccd1 _15911_/A sky130_fd_sc_hd__or3_4
XANTENNA__17087__A0 _15768_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13896__B1 _13845_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11207_ _19579_/Q vssd1 vssd1 vccd1 vccd1 _11460_/A sky130_fd_sc_hd__inv_2
X_19852_ _19859_/CLK _19852_/D repeater262/X vssd1 vssd1 vccd1 vccd1 _19852_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_96_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12187_ _12187_/A _12187_/B vssd1 vssd1 vccd1 vccd1 _12228_/A sky130_fd_sc_hd__or2_4
XFILLER_229_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18803_ _20059_/CLK _18803_/D repeater198/X vssd1 vssd1 vccd1 vccd1 _18803_/Q sky130_fd_sc_hd__dfrtp_2
X_11138_ _15222_/A _11144_/B vssd1 vssd1 vccd1 vccd1 _11139_/A sky130_fd_sc_hd__or2_1
XFILLER_122_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19783_ _20057_/CLK _19783_/D repeater203/X vssd1 vssd1 vccd1 vccd1 _19783_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18710__RESET_B repeater253/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16995_ _16994_/X _13871_/Y _17545_/S vssd1 vssd1 vccd1 vccd1 _16995_/X sky130_fd_sc_hd__mux2_1
XFILLER_95_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18734_ _19224_/CLK _18734_/D repeater186/X vssd1 vssd1 vccd1 vccd1 _18734_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_237_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11069_ _19848_/Q vssd1 vssd1 vccd1 vccd1 _14489_/B sky130_fd_sc_hd__clkbuf_2
X_15946_ _18235_/Q vssd1 vssd1 vccd1 vccd1 _15946_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18665_ _19812_/CLK _18665_/D repeater222/X vssd1 vssd1 vccd1 vccd1 _18665_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_92_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19987__RESET_B repeater193/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_225_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15877_ _19905_/Q vssd1 vssd1 vccd1 vccd1 _15877_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17650__S _17655_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17616_ _20056_/Q _19730_/Q _17621_/S vssd1 vssd1 vccd1 vccd1 _17616_/X sky130_fd_sc_hd__mux2_1
XFILLER_63_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14828_ _18156_/Q _14821_/A hold263/X _14822_/A vssd1 vssd1 vccd1 vccd1 _18156_/D
+ sky130_fd_sc_hd__a22o_1
X_18596_ _19577_/CLK _18596_/D repeater267/X vssd1 vssd1 vccd1 vccd1 _18596_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_17_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_130_HCLK clkbuf_4_4_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19582_/CLK sky130_fd_sc_hd__clkbuf_16
X_17547_ _17546_/X _11324_/Y _17547_/S vssd1 vssd1 vccd1 vccd1 _17547_/X sky130_fd_sc_hd__mux2_1
X_14759_ _14760_/A vssd1 vssd1 vccd1 vccd1 _14759_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_205_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18478__CLK _19780_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17478_ _17477_/X _15964_/Y _17523_/S vssd1 vssd1 vccd1 vccd1 _17478_/X sky130_fd_sc_hd__mux2_1
X_19217_ _19221_/CLK _19217_/D hold365/X vssd1 vssd1 vccd1 vccd1 _19217_/Q sky130_fd_sc_hd__dfrtp_1
X_16429_ _17960_/Q vssd1 vssd1 vccd1 vccd1 _16429_/Y sky130_fd_sc_hd__inv_2
XFILLER_158_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12095__A hold315/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12387__B1 _12386_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19148_ _19597_/CLK _19148_/D repeater281/X vssd1 vssd1 vccd1 vccd1 _19148_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17314__A1 _17844_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17097__S _17523_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19079_ _19115_/CLK _19079_/D hold353/X vssd1 vssd1 vccd1 vccd1 _19079_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_133_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18869__RESET_B repeater195/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12139__B1 _12074_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16825__A0 _17473_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09803_ _09803_/A vssd1 vssd1 vccd1 vccd1 _09803_/Y sky130_fd_sc_hd__inv_2
XFILLER_141_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_219_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09734_ _09734_/A vssd1 vssd1 vccd1 vccd1 _09813_/C sky130_fd_sc_hd__buf_2
XFILLER_28_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09665_ _09751_/A _09750_/A _09753_/A _09752_/A vssd1 vssd1 vccd1 vccd1 _09666_/C
+ sky130_fd_sc_hd__or4_4
XFILLER_39_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17560__S _17565_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_199_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19657__RESET_B repeater270/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09596_ _20019_/Q _09595_/Y _09585_/X _09480_/B vssd1 vssd1 vccd1 vccd1 _20019_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11417__A2 _19132_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17553__A1 _20036_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16904__S _17541_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10440_ _19837_/Q _10433_/X _09071_/X _10435_/X vssd1 vssd1 vccd1 vccd1 _19837_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_148_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10371_ _10371_/A vssd1 vssd1 vccd1 vccd1 _10372_/B sky130_fd_sc_hd__inv_2
XFILLER_136_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12110_ _19309_/Q _12106_/X _12026_/X _12108_/X vssd1 vssd1 vccd1 vccd1 _19309_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_108_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13090_ _13090_/A vssd1 vssd1 vccd1 vccd1 _13090_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_11_HCLK clkbuf_4_2_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _18260_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_156_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17735__S _18508_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12041_ _19339_/Q _12034_/X _11911_/X _12036_/X vssd1 vssd1 vccd1 vccd1 _19339_/D
+ sky130_fd_sc_hd__a22o_1
Xhold280 HWDATA[28] vssd1 vssd1 vccd1 vccd1 input58/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold291 input61/X vssd1 vssd1 vccd1 vccd1 hold291/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10253__A _19498_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16816__A0 _15963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11353__B2 _18969_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_238_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15800_ _16115_/A vssd1 vssd1 vccd1 vccd1 _16096_/B sky130_fd_sc_hd__buf_2
XFILLER_172_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16780_ _16720_/Y _19395_/Q _17413_/S vssd1 vssd1 vccd1 vccd1 _16780_/X sky130_fd_sc_hd__mux2_1
X_13992_ _18682_/Q vssd1 vssd1 vccd1 vccd1 _14012_/A sky130_fd_sc_hd__inv_2
XFILLER_207_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_153_HCLK clkbuf_4_1_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _18795_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_74_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15731_ _19875_/Q vssd1 vssd1 vccd1 vccd1 _15731_/Y sky130_fd_sc_hd__clkinv_4
X_12943_ _19276_/Q _12964_/C _19276_/Q _12964_/C vssd1 vssd1 vccd1 vccd1 _12943_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_46_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17241__A0 _15768_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17470__S _17566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10864__B1 _10863_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18450_ _18460_/CLK _18450_/D vssd1 vssd1 vccd1 vccd1 _18450_/Q sky130_fd_sc_hd__dfxtp_1
X_12874_ _12964_/D _12997_/A vssd1 vssd1 vccd1 vccd1 _12875_/B sky130_fd_sc_hd__or2_2
X_15662_ _15661_/A _15661_/B _15661_/Y vssd1 vssd1 vccd1 vccd1 _15663_/B sky130_fd_sc_hd__a21oi_1
XPHY_4240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19746__CLK _20070_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17401_ _17400_/X _16174_/Y _17565_/S vssd1 vssd1 vccd1 vccd1 _17401_/X sky130_fd_sc_hd__mux2_1
XPHY_4273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11825_ _19443_/Q _11821_/X _10861_/X _11822_/X vssd1 vssd1 vccd1 vccd1 _19443_/D
+ sky130_fd_sc_hd__a22o_1
X_14613_ _14613_/A vssd1 vssd1 vccd1 vccd1 _15195_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_233_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18381_ _19515_/CLK _18381_/D vssd1 vssd1 vccd1 vccd1 _18381_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_output102_A _16735_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15593_ _15593_/A vssd1 vssd1 vccd1 vccd1 _15598_/B sky130_fd_sc_hd__inv_2
XPHY_4284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14395__A _14395_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14544_ _15070_/A vssd1 vssd1 vccd1 vccd1 _14598_/A sky130_fd_sc_hd__buf_1
X_17332_ _17331_/X _13066_/A _17488_/S vssd1 vssd1 vccd1 vccd1 _17332_/X sky130_fd_sc_hd__mux2_1
XPHY_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11756_ hold145/X _11750_/X _19486_/Q _11751_/X vssd1 vssd1 vccd1 vccd1 hold147/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_14_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17544__A1 _14072_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10707_ _19775_/Q vssd1 vssd1 vccd1 vccd1 _10707_/Y sky130_fd_sc_hd__inv_2
XPHY_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14475_ _18354_/Q _14464_/A _14474_/X _14465_/A vssd1 vssd1 vccd1 vccd1 _18354_/D
+ sky130_fd_sc_hd__a22o_1
X_17263_ _17262_/X _09863_/A _17524_/S vssd1 vssd1 vccd1 vccd1 _17263_/X sky130_fd_sc_hd__mux2_2
X_11687_ _10522_/B _11674_/X _10735_/B _11675_/X vssd1 vssd1 vccd1 vccd1 _19530_/D
+ sky130_fd_sc_hd__o22ai_1
XPHY_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16814__S _17490_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater252_A repeater253/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19002_ _19137_/CLK _19002_/D hold348/X vssd1 vssd1 vccd1 vccd1 _19002_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__12369__B1 _12241_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13426_ _13443_/A vssd1 vssd1 vccd1 vccd1 _13426_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_201_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16214_ _16616_/A vssd1 vssd1 vccd1 vccd1 _16469_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_128_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10638_ _18555_/Q vssd1 vssd1 vccd1 vccd1 _10638_/Y sky130_fd_sc_hd__inv_2
X_17194_ _15768_/Y _11225_/Y _17546_/S vssd1 vssd1 vccd1 vccd1 _17194_/X sky130_fd_sc_hd__mux2_1
X_16145_ _17414_/X _16069_/X _17411_/X _16070_/X _16144_/X vssd1 vssd1 vccd1 vccd1
+ _16145_/X sky130_fd_sc_hd__o221a_1
X_13357_ _20122_/Q vssd1 vssd1 vccd1 vccd1 _13357_/Y sky130_fd_sc_hd__inv_2
X_10569_ _10569_/A vssd1 vssd1 vccd1 vccd1 _10615_/A sky130_fd_sc_hd__inv_2
XANTENNA__12643__A _12650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12308_ _19193_/Q _12276_/A _12241_/X _12277_/A vssd1 vssd1 vccd1 vccd1 _19193_/D
+ sky130_fd_sc_hd__a22o_1
X_16076_ _15749_/B _16068_/X _16072_/X _16074_/X _16075_/X vssd1 vssd1 vccd1 vccd1
+ _16076_/X sky130_fd_sc_hd__o2111a_2
X_13288_ _13254_/Y _13278_/X _13268_/Y _13287_/X vssd1 vssd1 vccd1 vccd1 _18870_/D
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__13869__B1 _19210_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17645__S _17655_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15027_ _18040_/Q _15023_/X _14996_/X _15025_/X vssd1 vssd1 vccd1 vccd1 _18040_/D
+ sky130_fd_sc_hd__a22o_1
X_19904_ _20123_/CLK _19904_/D repeater195/X vssd1 vssd1 vccd1 vccd1 _19904_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_130_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12239_ _19228_/Q _12205_/A _12238_/X _12206_/A vssd1 vssd1 vccd1 vccd1 _19228_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_142_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16807__A0 _15963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19835_ _20058_/CLK _19835_/D repeater194/X vssd1 vssd1 vccd1 vccd1 _19835_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__17480__A0 _15963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19766_ _19771_/CLK _19766_/D repeater189/X vssd1 vssd1 vccd1 vccd1 _19766_/Q sky130_fd_sc_hd__dfstp_1
X_16978_ _16977_/X _19146_/Q _17548_/S vssd1 vssd1 vccd1 vccd1 _16978_/X sky130_fd_sc_hd__mux2_1
XANTENNA__14294__B1 _13674_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_237_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput4 input4/A vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_1
X_18717_ _18718_/CLK _18717_/D repeater253/X vssd1 vssd1 vccd1 vccd1 _18717_/Q sky130_fd_sc_hd__dfrtp_1
X_15929_ _18147_/Q vssd1 vssd1 vccd1 vccd1 _15929_/Y sky130_fd_sc_hd__inv_2
X_19697_ _19720_/CLK _19697_/D repeater201/X vssd1 vssd1 vccd1 vccd1 _19697_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_237_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17380__S _17518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09450_ _10039_/A _19383_/Q _19911_/Q _09449_/Y vssd1 vssd1 vccd1 vccd1 _09450_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_18648_ _20050_/CLK _18648_/D repeater200/X vssd1 vssd1 vccd1 vccd1 _18648_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_225_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_240_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09381_ _19372_/Q vssd1 vssd1 vccd1 vccd1 _09381_/Y sky130_fd_sc_hd__inv_2
X_18579_ _19470_/CLK _18579_/D repeater273/X vssd1 vssd1 vccd1 vccd1 _18579_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_178_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09399__A _19390_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_34_HCLK _18641_/CLK vssd1 vssd1 vccd1 vccd1 _20079_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__17299__A0 _15963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16510__A2 _15904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15864__A _15867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_248_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19838__RESET_B repeater271/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14285__B1 _13682_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold178_A HADDR[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09717_ _19413_/Q vssd1 vssd1 vccd1 vccd1 _09717_/Y sky130_fd_sc_hd__inv_2
XFILLER_216_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17223__A0 _15768_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17290__S _17414_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10846__B1 _10446_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19491__RESET_B repeater260/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09648_ _19987_/Q vssd1 vssd1 vccd1 vccd1 _09743_/A sky130_fd_sc_hd__inv_2
XFILLER_216_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19420__RESET_B repeater192/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_215_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09579_ _09488_/A _09579_/A2 _09577_/Y _09604_/B vssd1 vssd1 vccd1 vccd1 _20028_/D
+ sky130_fd_sc_hd__a211oi_4
XPHY_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08939__A2_N _18779_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11610_ _19563_/Q _11609_/Y _11588_/A _11577_/B vssd1 vssd1 vccd1 vccd1 _19563_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12590_ _12598_/A vssd1 vssd1 vccd1 vccd1 _12590_/X sky130_fd_sc_hd__clkbuf_2
XPHY_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11541_ _11541_/A vssd1 vssd1 vccd1 vccd1 _11541_/Y sky130_fd_sc_hd__inv_2
XPHY_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16734__C1 _16733_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10248__A _10954_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14260_ _14260_/A vssd1 vssd1 vccd1 vccd1 _14260_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_rebuffer36_A _19418_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11472_ _11472_/A _11472_/B vssd1 vssd1 vccd1 vccd1 _11517_/A sky130_fd_sc_hd__or2_1
XPHY_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13211_ _18890_/Q _13210_/Y _13180_/A _13211_/C1 vssd1 vssd1 vccd1 vccd1 _18890_/D
+ sky130_fd_sc_hd__o211a_1
X_10423_ _10423_/A vssd1 vssd1 vccd1 vccd1 _10423_/X sky130_fd_sc_hd__buf_4
X_14191_ _19102_/Q vssd1 vssd1 vccd1 vccd1 _14191_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13142_ _19180_/Q _13081_/A _16645_/A _18909_/Q vssd1 vssd1 vccd1 vccd1 _13142_/X
+ sky130_fd_sc_hd__o22a_1
X_10354_ _10354_/A vssd1 vssd1 vccd1 vccd1 _10354_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__19299__CLK _20013_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11079__A _15858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17465__S _17566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15774__A _15774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17950_ _20079_/CLK _17950_/D vssd1 vssd1 vccd1 vccd1 _17950_/Q sky130_fd_sc_hd__dfxtp_1
X_13073_ _13073_/A _13073_/B vssd1 vssd1 vccd1 vccd1 _13190_/A sky130_fd_sc_hd__or2_1
X_10285_ _10181_/A _10759_/C _19872_/Q vssd1 vssd1 vccd1 vccd1 _10286_/B sky130_fd_sc_hd__o21a_1
XANTENNA__16589__B _16622_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16901_ _16900_/X _15561_/Y _17513_/S vssd1 vssd1 vccd1 vccd1 _16901_/X sky130_fd_sc_hd__mux2_1
X_12024_ _12044_/A vssd1 vssd1 vccd1 vccd1 _12024_/X sky130_fd_sc_hd__buf_1
XFILLER_105_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17881_ _16082_/Y _16083_/Y _16084_/Y _16085_/Y _17913_/S0 _19632_/Q vssd1 vssd1
+ vccd1 vccd1 _17881_/X sky130_fd_sc_hd__mux4_2
X_19620_ _19920_/CLK _19620_/D repeater230/X vssd1 vssd1 vccd1 vccd1 _19620_/Q sky130_fd_sc_hd__dfrtp_1
X_16832_ _15963_/X _12734_/Y _17534_/S vssd1 vssd1 vccd1 vccd1 _16832_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11807__A _11821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14276__B1 _14273_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_219_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19551_ _19561_/CLK _19551_/D repeater274/X vssd1 vssd1 vccd1 vccd1 _19551_/Q sky130_fd_sc_hd__dfrtp_1
X_16763_ _15963_/X _12767_/Y _17534_/S vssd1 vssd1 vccd1 vccd1 _16763_/X sky130_fd_sc_hd__mux2_1
XFILLER_76_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16809__S _17536_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13975_ _18699_/Q vssd1 vssd1 vccd1 vccd1 _14029_/A sky130_fd_sc_hd__inv_2
XFILLER_46_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18502_ _19795_/CLK _18502_/D repeater219/X vssd1 vssd1 vccd1 vccd1 _18502_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_202_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15714_ _15714_/A _15715_/B vssd1 vssd1 vccd1 vccd1 _18649_/D sky130_fd_sc_hd__nor2_1
X_19482_ _19506_/CLK hold164/X repeater260/X vssd1 vssd1 vccd1 vccd1 _19482_/Q sky130_fd_sc_hd__dfrtp_1
X_12926_ _19282_/Q vssd1 vssd1 vccd1 vccd1 _12926_/Y sky130_fd_sc_hd__inv_2
X_16694_ _16765_/X _16633_/X _17021_/X _16634_/X vssd1 vssd1 vccd1 vccd1 _16694_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_207_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18433_ _18795_/CLK _18433_/D vssd1 vssd1 vccd1 vccd1 _18433_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__19161__RESET_B hold370/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15645_ _18605_/Q vssd1 vssd1 vccd1 vccd1 _15645_/Y sky130_fd_sc_hd__inv_2
XPHY_4070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17860__S1 _19632_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12857_ _18921_/Q vssd1 vssd1 vccd1 vccd1 _12859_/B sky130_fd_sc_hd__inv_6
XPHY_4081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18364_ _18795_/CLK _18364_/D vssd1 vssd1 vccd1 vccd1 _18364_/Q sky130_fd_sc_hd__dfxtp_1
X_11808_ _11822_/A vssd1 vssd1 vccd1 vccd1 _11808_/X sky130_fd_sc_hd__clkbuf_2
X_12788_ _12786_/Y _18819_/Q _19242_/Q _13542_/A vssd1 vssd1 vccd1 vccd1 _12788_/X
+ sky130_fd_sc_hd__o22a_1
X_15576_ _15702_/A vssd1 vssd1 vccd1 vccd1 _15610_/A sky130_fd_sc_hd__buf_4
XPHY_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_57_HCLK clkbuf_4_12_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20048_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17315_ _16415_/X _19833_/Q _17566_/S vssd1 vssd1 vccd1 vccd1 _17315_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09012__A _10842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11739_ _19500_/Q _11737_/X _16932_/X _11738_/X vssd1 vssd1 vccd1 vccd1 hold222/A
+ sky130_fd_sc_hd__a22o_1
X_14527_ _18323_/Q _14519_/A hold334/X _14520_/A vssd1 vssd1 vccd1 vccd1 _18323_/D
+ sky130_fd_sc_hd__a22o_1
X_18295_ _18435_/CLK _18295_/D vssd1 vssd1 vccd1 vccd1 _18295_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_202_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17246_ _16588_/Y _17246_/A1 _17487_/S vssd1 vssd1 vccd1 vccd1 _17246_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14458_ _18365_/Q _14451_/X _14417_/X _14453_/X vssd1 vssd1 vccd1 vccd1 _18365_/D
+ sky130_fd_sc_hd__a22o_1
X_13409_ _20106_/Q vssd1 vssd1 vccd1 vccd1 _13409_/Y sky130_fd_sc_hd__clkinvlp_2
XFILLER_190_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14389_ _18403_/Q _14381_/A _12731_/X _14382_/A vssd1 vssd1 vccd1 vccd1 _18403_/D
+ sky130_fd_sc_hd__a22o_1
X_17177_ _17176_/X _12951_/Y _17541_/S vssd1 vssd1 vccd1 vccd1 _17177_/X sky130_fd_sc_hd__mux2_1
XFILLER_183_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16128_ _19676_/Q vssd1 vssd1 vccd1 vccd1 _16128_/Y sky130_fd_sc_hd__inv_2
XFILLER_170_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17375__S _17566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08950_ _19855_/Q vssd1 vssd1 vccd1 vccd1 _10321_/D sky130_fd_sc_hd__inv_2
X_16059_ _19767_/Q vssd1 vssd1 vccd1 vccd1 _16059_/Y sky130_fd_sc_hd__inv_2
XFILLER_143_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12514__B1 _12413_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19818_ _19822_/CLK _19818_/D repeater228/X vssd1 vssd1 vccd1 vccd1 _19818_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__11717__A _11731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19749_ _20070_/CLK _19749_/D repeater204/X vssd1 vssd1 vccd1 vccd1 _19749_/Q sky130_fd_sc_hd__dfrtp_2
X_09502_ _20023_/Q _09501_/Y _09478_/A _19308_/Q vssd1 vssd1 vccd1 vccd1 _09502_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_37_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13490__A1 _13483_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17756__A1 _12058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09433_ _19927_/Q _09431_/Y _10009_/B _19393_/Q vssd1 vssd1 vccd1 vccd1 _09433_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_213_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17851__S1 _19632_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09364_ _20013_/Q vssd1 vssd1 vccd1 vccd1 _09474_/B sky130_fd_sc_hd__inv_2
XFILLER_240_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17508__A1 _17904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15859__A _15859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09295_ _20044_/Q _09293_/X _09094_/X _09294_/X vssd1 vssd1 vccd1 vccd1 _20044_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_193_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18813__RESET_B repeater239/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16731__A2 _16493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17285__S _17546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16495__B2 _16683_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13411__A1_N _20108_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold295_A HWDATA[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10070_ _10040_/A _10040_/B _10032_/A _10068_/Y vssd1 vssd1 vccd1 vccd1 _19924_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_130_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14003__A _14003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10250__B _19515_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13760_ _17763_/S _13760_/B vssd1 vssd1 vccd1 vccd1 _13760_/X sky130_fd_sc_hd__or2_2
XFILLER_43_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10972_ _10978_/A vssd1 vssd1 vccd1 vccd1 _10973_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__17747__A1 _11059_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12711_ _12711_/A vssd1 vssd1 vccd1 vccd1 _12711_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_243_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13691_ _18767_/Q _13685_/X _13682_/X _13686_/Y vssd1 vssd1 vccd1 vccd1 _18767_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12458__A _12458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17842__S1 _19632_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15430_ _19621_/Q _11166_/B _11167_/B vssd1 vssd1 vccd1 vccd1 _15430_/X sky130_fd_sc_hd__a21bo_1
XPHY_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12642_ _19004_/Q _12636_/X _12032_/A _12637_/X vssd1 vssd1 vccd1 vccd1 _19004_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_31_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13233__B2 _17584_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14430__B1 _14415_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15361_ _18502_/Q _14232_/B _14233_/B vssd1 vssd1 vccd1 vccd1 _15361_/X sky130_fd_sc_hd__a21bo_1
XFILLER_178_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12573_ _19049_/Q _12569_/X _12394_/X _12570_/X vssd1 vssd1 vccd1 vccd1 _19049_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15769__A _15769_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17100_ _17099_/X _09396_/Y _17413_/S vssd1 vssd1 vccd1 vccd1 _17100_/X sky130_fd_sc_hd__mux2_1
XPHY_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14312_ hold335/X vssd1 vssd1 vccd1 vccd1 _14312_/X sky130_fd_sc_hd__buf_2
X_11524_ _11470_/A _11470_/B _11523_/X _11520_/Y vssd1 vssd1 vccd1 vccd1 _19590_/D
+ sky130_fd_sc_hd__a211oi_2
XPHY_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15292_ _15211_/A _15216_/C _15217_/Y vssd1 vssd1 vccd1 vccd1 _15292_/X sky130_fd_sc_hd__o21a_1
XFILLER_184_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18080_ _18137_/CLK _18080_/D vssd1 vssd1 vccd1 vccd1 _18080_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14243_ _18508_/Q vssd1 vssd1 vccd1 vccd1 _15334_/A sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_148_HCLK_A clkbuf_4_1_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17031_ _17473_/A0 _16692_/Y _17042_/S vssd1 vssd1 vccd1 vccd1 _17031_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11455_ _19573_/Q _11450_/Y _11626_/A _19136_/Q _11454_/X vssd1 vssd1 vccd1 vccd1
+ _11456_/D sky130_fd_sc_hd__o221a_1
XFILLER_194_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10406_ _10404_/A _14378_/B _10404_/Y vssd1 vssd1 vccd1 vccd1 _19848_/D sky130_fd_sc_hd__a21oi_1
X_14174_ _14172_/Y _18700_/Q _14173_/Y _18690_/Q vssd1 vssd1 vccd1 vccd1 _14174_/X
+ sky130_fd_sc_hd__o22a_1
X_11386_ _19147_/Q vssd1 vssd1 vccd1 vccd1 _11386_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17195__S _17459_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13125_ _13123_/Y _18897_/Q _16618_/A _18907_/Q vssd1 vssd1 vccd1 vccd1 _13125_/X
+ sky130_fd_sc_hd__o22a_1
X_10337_ _19867_/Q _10320_/X _10335_/A _08927_/Y _10336_/X vssd1 vssd1 vccd1 vccd1
+ _10338_/A sky130_fd_sc_hd__o32a_1
XFILLER_140_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18982_ _19608_/CLK _18982_/D hold355/X vssd1 vssd1 vccd1 vccd1 _18982_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_3_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17933_ _18465_/CLK _17933_/D vssd1 vssd1 vccd1 vccd1 _17933_/Q sky130_fd_sc_hd__dfxtp_1
X_13056_ _18890_/Q vssd1 vssd1 vccd1 vccd1 _13063_/A sky130_fd_sc_hd__inv_2
X_10268_ _19647_/Q _10268_/B vssd1 vssd1 vccd1 vccd1 _11039_/B sky130_fd_sc_hd__nand2_1
XFILLER_79_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12007_ _19359_/Q _12000_/X _09025_/X _12003_/X vssd1 vssd1 vccd1 vccd1 _19359_/D
+ sky130_fd_sc_hd__a22o_1
X_17864_ _17860_/X _17861_/X _17862_/X _17863_/X _19633_/Q _19634_/Q vssd1 vssd1 vccd1
+ vccd1 _17864_/X sky130_fd_sc_hd__mux4_2
XFILLER_238_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10199_ _19835_/Q _10962_/A _10198_/Y _19662_/Q vssd1 vssd1 vccd1 vccd1 _10209_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_213_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19603_ _19610_/CLK _19603_/D hold343/X vssd1 vssd1 vccd1 vccd1 _19603_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_78_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16815_ _16814_/X _13835_/Y _17545_/S vssd1 vssd1 vccd1 vccd1 _16815_/X sky130_fd_sc_hd__mux2_1
XFILLER_93_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17795_ _18320_/Q _18440_/Q _18432_/Q _18424_/Q _17923_/S0 _19646_/Q vssd1 vssd1
+ vccd1 vccd1 _17795_/X sky130_fd_sc_hd__mux4_1
X_19534_ _19544_/CLK _19534_/D repeater221/X vssd1 vssd1 vccd1 vccd1 _19534_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_53_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16746_ _16174_/Y _16271_/Y _16094_/Y _16173_/X _16745_/X vssd1 vssd1 vccd1 vccd1
+ _16747_/B sky130_fd_sc_hd__o221a_2
X_13958_ _18711_/Q _13957_/Y _13949_/B _13925_/X vssd1 vssd1 vccd1 vccd1 _18711_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_234_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19465_ _19470_/CLK _19465_/D repeater274/X vssd1 vssd1 vccd1 vccd1 _19465_/Q sky130_fd_sc_hd__dfrtp_1
X_12909_ _19286_/Q vssd1 vssd1 vccd1 vccd1 _12909_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17833__S1 _18750_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16677_ _17056_/X _16597_/X _17060_/X _16598_/X vssd1 vssd1 vccd1 vccd1 _16678_/D
+ sky130_fd_sc_hd__a22o_2
X_13889_ _13887_/Y _18707_/Q _13888_/Y _18722_/Q vssd1 vssd1 vccd1 vccd1 _13889_/X
+ sky130_fd_sc_hd__o22a_1
X_18416_ _18416_/CLK _18416_/D vssd1 vssd1 vccd1 vccd1 _18416_/Q sky130_fd_sc_hd__dfxtp_1
X_15628_ _18601_/Q vssd1 vssd1 vccd1 vccd1 _15628_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_222_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19396_ _20091_/CLK _19396_/D repeater236/X vssd1 vssd1 vccd1 vccd1 _19396_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__14421__B1 _14403_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11235__B1 _11487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18347_ _18954_/CLK _18347_/D vssd1 vssd1 vccd1 vccd1 _18347_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15559_ _18583_/Q vssd1 vssd1 vccd1 vccd1 _15559_/Y sky130_fd_sc_hd__inv_2
XFILLER_175_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09080_ _20099_/Q _09069_/X _09079_/X _09072_/X vssd1 vssd1 vccd1 vccd1 _20099_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_187_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18278_ _19847_/CLK _18278_/D vssd1 vssd1 vccd1 vccd1 _18278_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16713__A2 _16513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput40 input40/A vssd1 vssd1 vccd1 vccd1 input40/X sky130_fd_sc_hd__buf_1
X_17229_ _17228_/X _15480_/Y _17524_/S vssd1 vssd1 vccd1 vccd1 _17229_/X sky130_fd_sc_hd__mux2_1
XFILLER_238_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput51 input51/A vssd1 vssd1 vccd1 vccd1 input51/X sky130_fd_sc_hd__clkbuf_4
Xinput62 input62/A vssd1 vssd1 vccd1 vccd1 input62/X sky130_fd_sc_hd__buf_4
Xinput73 input73/A vssd1 vssd1 vccd1 vccd1 input73/X sky130_fd_sc_hd__buf_6
XFILLER_162_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08954__A2 _08952_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09982_ _19952_/Q _09981_/Y _09968_/X _09861_/B vssd1 vssd1 vccd1 vccd1 _19952_/D
+ sky130_fd_sc_hd__o211a_1
X_08933_ _19862_/Q vssd1 vssd1 vccd1 vccd1 _10328_/A sky130_fd_sc_hd__inv_2
XFILLER_115_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14660__B1 _14604_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_225_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17824__S1 _18752_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09416_ _09416_/A _09416_/B _09416_/C _09416_/D vssd1 vssd1 vccd1 vccd1 _09417_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_186_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14412__B1 _14351_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_9_HCLK clkbuf_4_2_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _18268_/CLK sky130_fd_sc_hd__clkbuf_16
X_09347_ _20030_/Q vssd1 vssd1 vccd1 vccd1 _09490_/A sky130_fd_sc_hd__inv_2
XFILLER_139_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11777__A1 hold193/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09278_ _20051_/Q _09270_/A _09105_/X _09271_/A vssd1 vssd1 vccd1 vccd1 _20051_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_166_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16912__S _17524_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11240_ _19600_/Q _16643_/A _11488_/A _19022_/Q vssd1 vssd1 vccd1 vccd1 _11240_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_180_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11171_ _19814_/Q vssd1 vssd1 vccd1 vccd1 _11173_/A sky130_fd_sc_hd__inv_2
XANTENNA__19853__RESET_B repeater267/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12741__A _19250_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10122_ _18572_/Q _18575_/Q _18579_/Q vssd1 vssd1 vccd1 vccd1 _10124_/C sky130_fd_sc_hd__or3_2
XFILLER_110_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17743__S _18508_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10053_ _10053_/A vssd1 vssd1 vccd1 vccd1 _10053_/X sky130_fd_sc_hd__clkbuf_2
X_14930_ _18094_/Q _14920_/X _14929_/X _14923_/X vssd1 vssd1 vccd1 vccd1 _18094_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19337__CLK _20013_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14861_ _18137_/Q _14858_/X _14699_/X _14860_/X vssd1 vssd1 vccd1 vccd1 _18137_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_180_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14100__C1 _14135_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16600_ _16600_/A _16600_/B _16600_/C _16600_/D vssd1 vssd1 vccd1 vccd1 _16600_/X
+ sky130_fd_sc_hd__or4_4
XFILLER_180_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13812_ _13950_/A _13949_/A _13812_/C _13951_/A vssd1 vssd1 vccd1 vccd1 _13813_/D
+ sky130_fd_sc_hd__or4_4
Xclkbuf_4_3_0_HCLK clkbuf_4_3_0_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_3_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_17580_ _15399_/X _19527_/Q _17584_/S vssd1 vssd1 vccd1 vccd1 _17580_/X sky130_fd_sc_hd__mux2_1
XFILLER_63_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14792_ _18174_/Q _14785_/X _14791_/X _14787_/X vssd1 vssd1 vccd1 vccd1 _18174_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_113_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16531_ _17181_/X _16684_/A _17172_/X _16493_/X vssd1 vssd1 vccd1 vccd1 _16531_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_244_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19487__CLK _19510_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10955_ _10978_/A vssd1 vssd1 vccd1 vccd1 _10955_/Y sky130_fd_sc_hd__inv_2
X_13743_ _17764_/X _13262_/B _13742_/X vssd1 vssd1 vccd1 vccd1 _18750_/D sky130_fd_sc_hd__a21oi_1
XFILLER_189_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12188__A _12228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17815__S1 _18750_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19250_ _19324_/CLK _19250_/D repeater237/X vssd1 vssd1 vccd1 vccd1 _19250_/Q sky130_fd_sc_hd__dfrtp_2
X_16462_ _17092_/X _16530_/A _17086_/X _16509_/A _16461_/X vssd1 vssd1 vccd1 vccd1
+ _16462_/X sky130_fd_sc_hd__o221a_2
XFILLER_232_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10886_ _19698_/Q _10875_/X _10885_/X _10879_/X vssd1 vssd1 vccd1 vccd1 _19698_/D
+ sky130_fd_sc_hd__a22o_1
X_13674_ hold325/X vssd1 vssd1 vccd1 vccd1 _13674_/X sky130_fd_sc_hd__buf_2
XFILLER_231_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18201_ _19630_/CLK _18201_/D vssd1 vssd1 vccd1 vccd1 _18201_/Q sky130_fd_sc_hd__dfxtp_1
X_15413_ _15413_/A _17574_/X vssd1 vssd1 vccd1 vccd1 _18538_/D sky130_fd_sc_hd__and2_1
XPHY_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12625_ _19017_/Q _12622_/X _12392_/X _12623_/X vssd1 vssd1 vccd1 vccd1 _19017_/D
+ sky130_fd_sc_hd__a22o_1
X_19181_ _19293_/CLK _19181_/D repeater187/X vssd1 vssd1 vccd1 vccd1 _19181_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16393_ _17332_/X _15997_/X _17335_/X _15998_/X _16392_/X vssd1 vssd1 vccd1 vccd1
+ _16393_/X sky130_fd_sc_hd__o221a_2
XPHY_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_repeater165_A _17543_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18132_ _18198_/CLK _18132_/D vssd1 vssd1 vccd1 vccd1 _18132_/Q sky130_fd_sc_hd__dfxtp_1
X_15344_ _18494_/Q _14224_/B _14225_/B vssd1 vssd1 vccd1 vccd1 _15344_/X sky130_fd_sc_hd__a21bo_1
X_12556_ _12556_/A _12556_/B vssd1 vssd1 vccd1 vccd1 _12556_/Y sky130_fd_sc_hd__nor2_1
XPHY_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11507_ _11480_/A _11480_/B _11506_/X _11503_/Y vssd1 vssd1 vccd1 vccd1 _19600_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_200_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18063_ _18465_/CLK _18063_/D vssd1 vssd1 vccd1 vccd1 _18063_/Q sky130_fd_sc_hd__dfxtp_1
X_15275_ _15275_/A vssd1 vssd1 vccd1 vccd1 _15275_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16822__S _17534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12487_ _12659_/A _12487_/B vssd1 vssd1 vccd1 vccd1 _12528_/A sky130_fd_sc_hd__or2_4
XANTENNA__14706__B2 _14701_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17014_ _17013_/X _09870_/A _17524_/S vssd1 vssd1 vccd1 vccd1 _17014_/X sky130_fd_sc_hd__mux2_2
X_14226_ _18496_/Q _14226_/B vssd1 vssd1 vccd1 vccd1 _14227_/B sky130_fd_sc_hd__or2_1
X_11438_ _19571_/Q vssd1 vssd1 vccd1 vccd1 _11584_/A sky130_fd_sc_hd__inv_2
XFILLER_99_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14157_ _14156_/Y _18688_/Q _19100_/Q _14010_/A vssd1 vssd1 vccd1 vccd1 _14157_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__13747__A _18870_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11369_ _19563_/Q vssd1 vssd1 vccd1 vccd1 _11576_/A sky130_fd_sc_hd__inv_2
XANTENNA__19594__RESET_B hold346/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12651__A _12651_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13108_ _13105_/Y _18894_/Q _19163_/Q _13065_/A _13107_/X vssd1 vssd1 vccd1 vccd1
+ _13109_/D sky130_fd_sc_hd__o221a_1
X_14088_ _19069_/Q _14011_/A _19086_/Q _14027_/A vssd1 vssd1 vccd1 vccd1 _14088_/X
+ sky130_fd_sc_hd__o22a_1
X_18965_ _19208_/CLK _18965_/D hold370/X vssd1 vssd1 vccd1 vccd1 _18965_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_113_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17653__S _17655_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17916_ _18193_/Q _18185_/Q _18177_/Q _18161_/Q _17918_/S0 _18750_/Q vssd1 vssd1
+ vccd1 vccd1 _17916_/X sky130_fd_sc_hd__mux4_2
X_13039_ _18907_/Q vssd1 vssd1 vccd1 vccd1 _13079_/A sky130_fd_sc_hd__inv_2
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18896_ _18908_/CLK _18896_/D hold372/X vssd1 vssd1 vccd1 vccd1 _18896_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__14890__B1 _14812_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17847_ _16355_/Y _16356_/Y _16357_/Y _16358_/Y _17908_/S0 _18759_/Q vssd1 vssd1
+ vccd1 vccd1 _17847_/X sky130_fd_sc_hd__mux4_1
XANTENNA__14578__A _14791_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17778_ _18292_/Q _18284_/Q _18276_/Q _18444_/Q _17923_/S0 _19646_/Q vssd1 vssd1
+ vccd1 vccd1 _17778_/X sky130_fd_sc_hd__mux4_2
XANTENNA__20081__RESET_B repeater204/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19517_ _19867_/CLK hold209/X repeater262/X vssd1 vssd1 vccd1 vccd1 _19517_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_207_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16729_ _19469_/Q vssd1 vssd1 vccd1 vccd1 _16729_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12098__A hold301/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17806__S1 _18750_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_241_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19448_ _20058_/CLK _19448_/D repeater194/X vssd1 vssd1 vccd1 vccd1 _19448_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_168_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16395__B1 _17329_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09201_ _20070_/Q _09199_/A _09198_/X _08978_/A _09200_/X vssd1 vssd1 vccd1 vccd1
+ _09202_/A sky130_fd_sc_hd__o32a_1
X_19379_ _19927_/CLK _19379_/D repeater230/X vssd1 vssd1 vccd1 vccd1 _19379_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_148_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09132_ _20087_/Q vssd1 vssd1 vccd1 vccd1 _15321_/A sky130_fd_sc_hd__buf_1
XANTENNA__11730__A _11730_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09063_ hold257/X vssd1 vssd1 vccd1 vccd1 _12030_/A sky130_fd_sc_hd__buf_4
XFILLER_190_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_131_HCLK_A clkbuf_4_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12184__A1 _19260_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13381__B1 _20099_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12561__A _12598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19264__RESET_B repeater245/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09965_ _19962_/Q _09963_/Y _09871_/B _09964_/X vssd1 vssd1 vccd1 vccd1 _19962_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__11177__A _11191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17563__S _17568_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08916_ _08982_/A _10132_/B vssd1 vssd1 vccd1 vccd1 _08917_/A sky130_fd_sc_hd__or2_4
X_20085_ _20085_/CLK _20085_/D repeater204/X vssd1 vssd1 vccd1 vccd1 _20085_/Q sky130_fd_sc_hd__dfrtp_1
X_09896_ _19333_/Q vssd1 vssd1 vccd1 vccd1 _09896_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11695__B1 _10885_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_hold160_A HADDR[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold258_A HWDATA[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16907__S _17545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10740_ _15826_/A _13252_/D vssd1 vssd1 vccd1 vccd1 _10742_/A sky130_fd_sc_hd__or2_2
XFILLER_214_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10671_ _17734_/X _10669_/X _19791_/Q _10670_/X vssd1 vssd1 vccd1 vccd1 _19791_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_13_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12736__A _19235_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12410_ hold294/X vssd1 vssd1 vccd1 vccd1 _12410_/X sky130_fd_sc_hd__buf_2
XANTENNA__12947__B1 _12945_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_11_0_HCLK clkbuf_3_5_0_HCLK/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_2_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_13390_ _20111_/Q vssd1 vssd1 vccd1 vccd1 _13390_/Y sky130_fd_sc_hd__inv_2
XFILLER_223_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17738__S _18508_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14149__C1 _14112_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12341_ _12361_/A vssd1 vssd1 vccd1 vccd1 _12341_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_181_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10256__A _19627_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15060_ _15060_/A vssd1 vssd1 vccd1 vccd1 _15061_/A sky130_fd_sc_hd__inv_2
XFILLER_181_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12272_ _19218_/Q _12269_/X _12086_/X _12270_/X vssd1 vssd1 vccd1 vccd1 _19218_/D
+ sky130_fd_sc_hd__a22o_1
X_14011_ _14011_/A _14011_/B vssd1 vssd1 vccd1 vccd1 _14012_/C sky130_fd_sc_hd__or2_2
XANTENNA__12175__A1 _19266_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11223_ _11223_/A _11223_/B _11223_/C _11223_/D vssd1 vssd1 vccd1 vccd1 _11223_/X
+ sky130_fd_sc_hd__and4_1
XANTENNA__09040__A1 _20113_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12471__A _12478_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_53_HCLK_A clkbuf_4_9_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11154_ _11150_/X _11152_/X _11022_/X _11153_/Y _17756_/X vssd1 vssd1 vccd1 vccd1
+ _11155_/A sky130_fd_sc_hd__o32a_1
XFILLER_68_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10105_ _10011_/B _10104_/A _19908_/Q _10107_/A _10053_/X vssd1 vssd1 vccd1 vccd1
+ _19908_/D sky130_fd_sc_hd__o221a_1
XANTENNA__17473__S _17473_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18750_ _19900_/CLK _18750_/D repeater199/X vssd1 vssd1 vccd1 vccd1 _18750_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_1_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11085_ _12551_/A _12553_/A _11085_/C vssd1 vssd1 vccd1 vccd1 _12246_/B sky130_fd_sc_hd__or3_1
X_15962_ _16436_/B _18738_/Q vssd1 vssd1 vccd1 vccd1 _15962_/X sky130_fd_sc_hd__and2_1
XFILLER_48_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_237_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17701_ _19817_/Q _19759_/Q _18548_/Q vssd1 vssd1 vccd1 vccd1 _17701_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10036_ _10036_/A _10036_/B vssd1 vssd1 vccd1 vccd1 _10074_/A sky130_fd_sc_hd__or2_1
X_14913_ _18103_/Q _14908_/X _14705_/X _14910_/X vssd1 vssd1 vccd1 vccd1 _18103_/D
+ sky130_fd_sc_hd__a22o_1
X_18681_ _18686_/CLK _18681_/D hold359/X vssd1 vssd1 vccd1 vccd1 _18681_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_102_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output132_A _19876_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15893_ _17536_/X _16493_/A _15892_/Y _15845_/D vssd1 vssd1 vccd1 vccd1 _15893_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_64_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17632_ _15716_/Y _10291_/B _18643_/Q vssd1 vssd1 vccd1 vccd1 _18643_/D sky130_fd_sc_hd__mux2_1
X_14844_ _14990_/A _15034_/B _15094_/C vssd1 vssd1 vccd1 vccd1 _14846_/A sky130_fd_sc_hd__or3_4
XFILLER_64_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17563_ _17562_/X _17909_/X _17568_/S vssd1 vssd1 vccd1 vccd1 _17563_/X sky130_fd_sc_hd__mux2_1
X_14775_ _18184_/Q _14771_/X _14749_/X _14773_/X vssd1 vssd1 vccd1 vccd1 _18184_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_223_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16817__S _17535_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11987_ _19366_/Q _11955_/A _11926_/X _11956_/A vssd1 vssd1 vccd1 vccd1 _19366_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_216_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19302_ _19952_/CLK _19302_/D repeater242/X vssd1 vssd1 vccd1 vccd1 _19302_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_210_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16514_ _17296_/X _15896_/X _17282_/X _16493_/X vssd1 vssd1 vccd1 vccd1 _16514_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_17_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13726_ _18756_/Q vssd1 vssd1 vccd1 vccd1 _14743_/A sky130_fd_sc_hd__clkbuf_2
X_10938_ _17606_/X _10938_/B vssd1 vssd1 vccd1 vccd1 _15298_/D sky130_fd_sc_hd__nand2_1
XFILLER_189_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17494_ _17493_/X _11420_/Y _17548_/S vssd1 vssd1 vccd1 vccd1 _17494_/X sky130_fd_sc_hd__mux2_2
X_19233_ _19314_/CLK _19233_/D repeater214/X vssd1 vssd1 vccd1 vccd1 _19233_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_231_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16445_ _19680_/Q vssd1 vssd1 vccd1 vccd1 _16445_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10869_ _19702_/Q _10856_/A _10868_/X _10857_/A vssd1 vssd1 vccd1 vccd1 _19702_/D
+ sky130_fd_sc_hd__a22o_1
X_13657_ _13671_/A vssd1 vssd1 vccd1 vccd1 _13672_/A sky130_fd_sc_hd__inv_2
XFILLER_158_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12608_ _19025_/Q _12576_/A _12543_/X _12577_/A vssd1 vssd1 vccd1 vccd1 _19025_/D
+ sky130_fd_sc_hd__a22o_1
X_19164_ _19214_/CLK _19164_/D hold367/X vssd1 vssd1 vccd1 vccd1 _19164_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16376_ _19679_/Q vssd1 vssd1 vccd1 vccd1 _16376_/Y sky130_fd_sc_hd__inv_2
XPHY_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13588_ _13588_/A vssd1 vssd1 vccd1 vccd1 _13588_/X sky130_fd_sc_hd__buf_2
XFILLER_191_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18115_ _18142_/CLK _18115_/D vssd1 vssd1 vccd1 vccd1 _18115_/Q sky130_fd_sc_hd__dfxtp_1
X_15327_ _10909_/A _15215_/B _18636_/Q _15326_/Y vssd1 vssd1 vccd1 vccd1 _18636_/D
+ sky130_fd_sc_hd__a31o_1
XANTENNA__17648__S _17655_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12539_ _19063_/Q _12528_/X _12538_/X _12529_/X vssd1 vssd1 vccd1 vccd1 _19063_/D
+ sky130_fd_sc_hd__a22o_1
X_19095_ _19585_/CLK _19095_/D hold365/X vssd1 vssd1 vccd1 vccd1 _19095_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_219_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19502__CLK _19510_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18046_ _18473_/CLK _18046_/D vssd1 vssd1 vccd1 vccd1 _18046_/Q sky130_fd_sc_hd__dfxtp_1
X_15258_ _18634_/Q vssd1 vssd1 vccd1 vccd1 _15259_/B sky130_fd_sc_hd__inv_2
XFILLER_172_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14209_ _19113_/Q _14022_/A _19104_/Q _14013_/A _14208_/X vssd1 vssd1 vccd1 vccd1
+ _14218_/B sky130_fd_sc_hd__o221a_1
XFILLER_153_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15189_ _17930_/Q _14251_/A _10423_/A _14252_/A vssd1 vssd1 vccd1 vccd1 _17930_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10177__B1 _09098_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19997_ _19997_/CLK _19997_/D repeater185/X vssd1 vssd1 vccd1 vccd1 _19997_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17383__S _17413_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09750_ _09750_/A _09750_/B vssd1 vssd1 vccd1 vccd1 _09769_/A sky130_fd_sc_hd__or2_1
XFILLER_140_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18948_ _19290_/CLK _18948_/D repeater211/X vssd1 vssd1 vccd1 vccd1 _18948_/Q sky130_fd_sc_hd__dfrtp_1
X_09681_ _19422_/Q vssd1 vssd1 vccd1 vccd1 _09681_/Y sky130_fd_sc_hd__inv_2
X_18879_ _20048_/CLK _18879_/D repeater191/X vssd1 vssd1 vccd1 vccd1 _18879_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_27_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18657__RESET_B repeater210/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15040__B1 _14998_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09115_ _09127_/A _09133_/C _20087_/Q _09138_/A vssd1 vssd1 vccd1 vccd1 _09139_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_13_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11092__A1_N _11059_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15867__A _15867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09046_ _20111_/Q _09041_/X hold300/X _09043_/X vssd1 vssd1 vccd1 vccd1 _20111_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__15894__A2 _15887_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17293__S _17566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09948_ _09948_/A _09948_/B _09948_/C _09948_/D vssd1 vssd1 vccd1 vccd1 _09990_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_219_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20068_ _20124_/CLK _20068_/D repeater207/X vssd1 vssd1 vccd1 vccd1 _20068_/Q sky130_fd_sc_hd__dfrtp_1
X_09879_ _19970_/Q vssd1 vssd1 vccd1 vccd1 _09879_/Y sky130_fd_sc_hd__inv_2
XFILLER_245_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16210__B _16212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11910_ _19410_/Q _11905_/X _11909_/X _11906_/X vssd1 vssd1 vccd1 vccd1 _19410_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_245_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12890_ _18948_/Q _12890_/B vssd1 vssd1 vccd1 vccd1 _12891_/B sky130_fd_sc_hd__nand2_1
XPHY_4411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11841_ _12313_/A vssd1 vssd1 vccd1 vccd1 _11841_/X sky130_fd_sc_hd__buf_1
XPHY_4444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12093__B1 _12092_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11772_ _11772_/A vssd1 vssd1 vccd1 vccd1 _11772_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14560_ _14560_/A vssd1 vssd1 vccd1 vccd1 _14560_/X sky130_fd_sc_hd__clkbuf_2
XPHY_4488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17020__A1 _09374_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10723_ _19772_/Q _10720_/X _10446_/X _10722_/X vssd1 vssd1 vccd1 vccd1 _19772_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11840__A0 _10147_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13511_ _13511_/A vssd1 vssd1 vccd1 vccd1 _14641_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_213_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14491_ _14492_/A vssd1 vssd1 vccd1 vccd1 _14491_/X sky130_fd_sc_hd__clkbuf_2
XPHY_3798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15031__B1 _15004_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16230_ _19819_/Q vssd1 vssd1 vccd1 vccd1 _16230_/Y sky130_fd_sc_hd__inv_2
X_13442_ _13442_/A vssd1 vssd1 vccd1 vccd1 _13442_/Y sky130_fd_sc_hd__inv_2
X_10654_ _19794_/Q _10654_/B vssd1 vssd1 vccd1 vccd1 _10655_/B sky130_fd_sc_hd__or2_1
XFILLER_158_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12185__B _12372_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_90_HCLK clkbuf_4_12_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20013_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__17468__S _17564_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13373_ _20109_/Q vssd1 vssd1 vccd1 vccd1 _13373_/Y sky130_fd_sc_hd__inv_4
XFILLER_186_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16161_ _18014_/Q vssd1 vssd1 vccd1 vccd1 _16161_/Y sky130_fd_sc_hd__inv_2
X_10585_ _19804_/Q _19803_/Q _10585_/C vssd1 vssd1 vccd1 vccd1 _10590_/D sky130_fd_sc_hd__or3_1
XFILLER_194_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15112_ _15112_/A vssd1 vssd1 vccd1 vccd1 _15112_/X sky130_fd_sc_hd__clkbuf_2
X_12324_ _19187_/Q _12318_/X _12076_/X _12321_/X vssd1 vssd1 vccd1 vccd1 _19187_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_182_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16092_ _18469_/Q vssd1 vssd1 vccd1 vccd1 _16092_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16531__B1 _17172_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19920_ _19920_/CLK _19920_/D repeater230/X vssd1 vssd1 vccd1 vccd1 _19920_/Q sky130_fd_sc_hd__dfrtp_1
X_15043_ _18028_/Q _15036_/A _15004_/X _15037_/A vssd1 vssd1 vccd1 vccd1 _18028_/D
+ sky130_fd_sc_hd__a22o_1
X_12255_ _15232_/A _12252_/S _15232_/B _12254_/Y vssd1 vssd1 vccd1 vccd1 _19225_/D
+ sky130_fd_sc_hd__o22ai_1
XANTENNA__10159__B1 _09090_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11206_ _19606_/Q vssd1 vssd1 vccd1 vccd1 _11486_/A sky130_fd_sc_hd__inv_2
X_19851_ _19851_/CLK _19851_/D repeater258/X vssd1 vssd1 vccd1 vccd1 _19851_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_122_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12186_ _12180_/X _19259_/Q _12186_/S vssd1 vssd1 vccd1 vccd1 _19259_/D sky130_fd_sc_hd__mux2_1
XFILLER_150_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11137_ _19226_/Q _11135_/X _12708_/B _17613_/X vssd1 vssd1 vccd1 vccd1 _11144_/B
+ sky130_fd_sc_hd__a211o_1
X_18802_ _20059_/CLK _18802_/D repeater199/X vssd1 vssd1 vccd1 vccd1 _18802_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_205_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19782_ _20055_/CLK _19782_/D repeater204/X vssd1 vssd1 vccd1 vccd1 _19782_/Q sky130_fd_sc_hd__dfrtp_1
X_16994_ _16993_/X _16657_/Y _17490_/S vssd1 vssd1 vccd1 vccd1 _16994_/X sky130_fd_sc_hd__mux2_2
XFILLER_122_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_237_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18733_ _19224_/CLK _18733_/D repeater186/X vssd1 vssd1 vccd1 vccd1 _18733_/Q sky130_fd_sc_hd__dfrtp_1
X_11068_ _11060_/Y _11067_/X _11060_/Y _11067_/X vssd1 vssd1 vccd1 vccd1 _11076_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_48_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15945_ _18251_/Q vssd1 vssd1 vccd1 vccd1 _15945_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10019_ _10037_/A _10036_/A _10019_/C _10019_/D vssd1 vssd1 vccd1 vccd1 _10021_/B
+ sky130_fd_sc_hd__or4_4
XANTENNA__11545__A _19024_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18664_ _19813_/CLK _18664_/D repeater225/X vssd1 vssd1 vccd1 vccd1 _18664_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_64_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15876_ _19439_/Q vssd1 vssd1 vccd1 vccd1 _15876_/Y sky130_fd_sc_hd__inv_2
XFILLER_221_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17615_ _20057_/Q _19731_/Q _17621_/S vssd1 vssd1 vccd1 vccd1 _17615_/X sky130_fd_sc_hd__mux2_1
XFILLER_224_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14827_ _18157_/Q _14820_/X _14793_/X _14822_/X vssd1 vssd1 vccd1 vccd1 _18157_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_36_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18595_ _19437_/CLK _18595_/D repeater269/X vssd1 vssd1 vccd1 vccd1 _18595_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_63_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17546_ _15862_/Y _11218_/Y _17546_/S vssd1 vssd1 vccd1 vccd1 _17546_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14758_ _14819_/A _14758_/B _14758_/C vssd1 vssd1 vccd1 vccd1 _14760_/A sky130_fd_sc_hd__or3_4
XFILLER_232_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13709_ _18761_/Q _13707_/Y _13708_/Y _13707_/A vssd1 vssd1 vccd1 vccd1 _18761_/D
+ sky130_fd_sc_hd__o22a_1
X_17477_ _17486_/A0 _09934_/Y _17543_/S vssd1 vssd1 vccd1 vccd1 _17477_/X sky130_fd_sc_hd__mux2_1
XANTENNA__19956__RESET_B repeater245/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14689_ _18229_/Q _14682_/X _14580_/X _14684_/X vssd1 vssd1 vccd1 vccd1 _18229_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_60_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11280__A _18997_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19216_ _19221_/CLK _19216_/D hold365/X vssd1 vssd1 vccd1 vccd1 _19216_/Q sky130_fd_sc_hd__dfrtp_1
X_16428_ _17984_/Q vssd1 vssd1 vccd1 vccd1 _16428_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14376__A2 _14368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19147_ _19597_/CLK _19147_/D repeater281/X vssd1 vssd1 vccd1 vccd1 _19147_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__17378__S _17564_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16359_ _17959_/Q vssd1 vssd1 vccd1 vccd1 _16359_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19078_ _19115_/CLK _19078_/D hold355/X vssd1 vssd1 vccd1 vccd1 _19078_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_8_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16522__B1 _17301_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18029_ _18145_/CLK _18029_/D vssd1 vssd1 vccd1 vccd1 _18029_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_246_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15089__B1 _14791_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09802_ _09790_/A _09790_/B _09800_/Y _09767_/X vssd1 vssd1 vccd1 vccd1 _19978_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_113_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09733_ _09735_/B vssd1 vssd1 vccd1 vccd1 _09734_/A sky130_fd_sc_hd__buf_2
XFILLER_101_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_227_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09664_ _19996_/Q vssd1 vssd1 vccd1 vccd1 _09752_/A sky130_fd_sc_hd__inv_2
XFILLER_82_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_215_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09595_ _09595_/A vssd1 vssd1 vccd1 vccd1 _09595_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12075__B1 _12074_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15013__B1 _14992_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_7_0_HCLK clkbuf_3_7_0_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__17288__S _17534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10370_ _10370_/A vssd1 vssd1 vccd1 vccd1 _19858_/D sky130_fd_sc_hd__inv_2
XFILLER_164_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09029_ _09041_/A vssd1 vssd1 vccd1 vccd1 _09029_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_164_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16920__S _17547_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12040_ _19340_/Q _12034_/X _11909_/X _12036_/X vssd1 vssd1 vccd1 vccd1 _19340_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17069__A1 _19390_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold270 hold270/A vssd1 vssd1 vccd1 vccd1 hold270/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11889__B1 _09037_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold281 hold281/A vssd1 vssd1 vccd1 vccd1 hold281/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11353__A2 _18981_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold292 HWDATA[30] vssd1 vssd1 vccd1 vccd1 input61/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_120_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14827__B1 _14793_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13991_ _18683_/Q vssd1 vssd1 vccd1 vccd1 _14013_/A sky130_fd_sc_hd__inv_2
XFILLER_58_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15730_ _20041_/Q _10788_/Y _15729_/Y _19738_/Q _10791_/A vssd1 vssd1 vccd1 vccd1
+ _17622_/S sky130_fd_sc_hd__a221oi_2
XFILLER_45_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12942_ _19274_/Q vssd1 vssd1 vccd1 vccd1 _12942_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15661_ _15661_/A _15661_/B vssd1 vssd1 vccd1 vccd1 _15661_/Y sky130_fd_sc_hd__nor2_1
XPHY_4230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12873_ _12965_/C _12873_/B vssd1 vssd1 vccd1 vccd1 _12997_/A sky130_fd_sc_hd__or2_1
XFILLER_45_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17400_ _16176_/Y _16175_/Y _17564_/S vssd1 vssd1 vccd1 vccd1 _17400_/X sky130_fd_sc_hd__mux2_1
XPHY_4252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14612_ _18274_/Q _14601_/A hold320/X _14602_/A vssd1 vssd1 vccd1 vccd1 _18274_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18380_ _19515_/CLK _18380_/D vssd1 vssd1 vccd1 vccd1 _18380_/Q sky130_fd_sc_hd__dfxtp_1
X_11824_ _19444_/Q _11821_/X _10885_/X _11822_/X vssd1 vssd1 vccd1 vccd1 _19444_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15592_ _18592_/Q vssd1 vssd1 vccd1 vccd1 _15594_/A sky130_fd_sc_hd__inv_2
XPHY_4285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17331_ _17330_/X _12933_/Y _17487_/S vssd1 vssd1 vccd1 vccd1 _17331_/X sky130_fd_sc_hd__mux2_1
XFILLER_199_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14543_ _18314_/Q _14532_/A _14474_/X _14533_/A vssd1 vssd1 vccd1 vccd1 _18314_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11813__B1 _09067_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11755_ hold159/X _11750_/X _19487_/Q _11751_/X vssd1 vssd1 vccd1 vccd1 hold161/A
+ sky130_fd_sc_hd__o22a_1
XPHY_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10706_ _10706_/A vssd1 vssd1 vccd1 vccd1 _19776_/D sky130_fd_sc_hd__inv_2
XPHY_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17262_ _17261_/X _09686_/Y _17523_/S vssd1 vssd1 vccd1 vccd1 _17262_/X sky130_fd_sc_hd__mux2_1
XFILLER_186_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14474_ hold321/X vssd1 vssd1 vccd1 vccd1 _14474_/X sky130_fd_sc_hd__buf_2
X_11686_ _19531_/Q _11668_/A _10527_/A _11669_/X vssd1 vssd1 vccd1 vccd1 _19531_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19001_ _19585_/CLK _19001_/D hold363/X vssd1 vssd1 vccd1 vccd1 _19001_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__17198__S _17493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12369__B2 _12335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16213_ _16669_/A vssd1 vssd1 vccd1 vccd1 _16616_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_13425_ _13354_/A _13354_/B _13355_/Y _13489_/C vssd1 vssd1 vccd1 vccd1 _18867_/D
+ sky130_fd_sc_hd__a211oi_2
X_10637_ _19798_/Q _10609_/A _10942_/A _10606_/X vssd1 vssd1 vccd1 vccd1 _19798_/D
+ sky130_fd_sc_hd__o22a_1
X_17193_ _17192_/X _11452_/Y _17548_/S vssd1 vssd1 vccd1 vccd1 _17193_/X sky130_fd_sc_hd__mux2_1
XFILLER_155_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11041__A1 _19648_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16144_ _17438_/X _15900_/A _17406_/X _15908_/A vssd1 vssd1 vccd1 vccd1 _16144_/X
+ sky130_fd_sc_hd__o22a_2
X_10568_ _10595_/A _19812_/Q _10582_/A _19811_/Q vssd1 vssd1 vccd1 vccd1 _10569_/A
+ sky130_fd_sc_hd__or4b_4
X_13356_ _18868_/Q vssd1 vssd1 vccd1 vccd1 _13356_/Y sky130_fd_sc_hd__inv_2
XFILLER_143_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12307_ _19194_/Q _12276_/A _12238_/X _12277_/A vssd1 vssd1 vccd1 vccd1 _19194_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_115_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16075_ _17442_/X _16002_/X _17451_/X _16003_/X vssd1 vssd1 vccd1 vccd1 _16075_/X
+ sky130_fd_sc_hd__o22a_1
X_10499_ _10519_/D _19534_/Q vssd1 vssd1 vccd1 vccd1 _10502_/B sky130_fd_sc_hd__nand2_1
XANTENNA__16830__S _17459_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13287_ _13750_/A vssd1 vssd1 vccd1 vccd1 _13287_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_216_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15026_ _18041_/Q _15023_/X _14992_/X _15025_/X vssd1 vssd1 vccd1 vccd1 _18041_/D
+ sky130_fd_sc_hd__a22o_1
X_19903_ _20123_/CLK _19903_/D repeater195/X vssd1 vssd1 vccd1 vccd1 _19903_/Q sky130_fd_sc_hd__dfrtp_1
X_12238_ _12238_/A vssd1 vssd1 vccd1 vccd1 _12238_/X sky130_fd_sc_hd__buf_6
XFILLER_123_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19834_ _20058_/CLK _19834_/D repeater194/X vssd1 vssd1 vccd1 vccd1 _19834_/Q sky130_fd_sc_hd__dfrtp_4
X_12169_ _19270_/Q _12164_/X _11911_/X _12165_/X vssd1 vssd1 vccd1 vccd1 _19270_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_111_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19765_ _19771_/CLK _19765_/D repeater189/X vssd1 vssd1 vccd1 vccd1 _19765_/Q sky130_fd_sc_hd__dfstp_1
X_16977_ _16615_/Y _18980_/Q _17493_/S vssd1 vssd1 vccd1 vccd1 _16977_/X sky130_fd_sc_hd__mux2_1
XFILLER_209_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput5 input5/A vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_1
X_15928_ _18011_/Q vssd1 vssd1 vccd1 vccd1 _15928_/Y sky130_fd_sc_hd__inv_2
X_18716_ _18718_/CLK _18716_/D repeater253/X vssd1 vssd1 vccd1 vccd1 _18716_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_237_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_209_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19696_ _19720_/CLK _19696_/D repeater201/X vssd1 vssd1 vccd1 vccd1 _19696_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_224_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18647_ _20050_/CLK _18647_/D repeater197/X vssd1 vssd1 vccd1 vccd1 _18647_/Q sky130_fd_sc_hd__dfrtp_1
X_15859_ _15859_/A vssd1 vssd1 vccd1 vccd1 _15859_/X sky130_fd_sc_hd__buf_4
XFILLER_240_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09380_ _19909_/Q vssd1 vssd1 vccd1 vccd1 _10011_/A sky130_fd_sc_hd__inv_4
X_18578_ _19437_/CLK _18578_/D repeater269/X vssd1 vssd1 vccd1 vccd1 _18578_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_240_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_233_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17529_ _17528_/X _09430_/Y _17529_/S vssd1 vssd1 vccd1 vccd1 _17529_/X sky130_fd_sc_hd__mux2_1
XANTENNA__19790__RESET_B repeater203/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11804__B1 hold317/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17918__S0 _17918_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19990__CLK _19992_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16025__B _16096_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14809__B1 _14808_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18672__RESET_B repeater252/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17471__A1 _11093_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17571__S _17584_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11185__A _11192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09716_ _09807_/C _19402_/Q _19977_/Q _09714_/Y _09715_/X vssd1 vssd1 vccd1 vccd1
+ _09716_/X sky130_fd_sc_hd__a221o_1
XFILLER_216_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09647_ _09788_/A _09787_/C _09647_/C _09647_/D vssd1 vssd1 vccd1 vccd1 _09739_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_27_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14037__B2 _18681_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12048__B1 _11920_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09578_ _20029_/Q _09577_/Y _09567_/X _09490_/B vssd1 vssd1 vccd1 vccd1 _20029_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_203_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11540_ _11461_/A _11540_/A2 _11523_/X _11538_/Y vssd1 vssd1 vccd1 vccd1 _19580_/D
+ sky130_fd_sc_hd__a211oi_2
XPHY_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19460__RESET_B repeater272/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11471_ _11471_/A _11520_/A vssd1 vssd1 vccd1 vccd1 _11472_/B sky130_fd_sc_hd__or2_2
XPHY_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17909__S0 _18760_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10422_ _19845_/Q _10417_/X _10421_/X _10419_/Y vssd1 vssd1 vccd1 vccd1 _19845_/D
+ sky130_fd_sc_hd__a22o_1
X_13210_ _13210_/A vssd1 vssd1 vccd1 vccd1 _13210_/Y sky130_fd_sc_hd__inv_2
X_14190_ _19116_/Q _18695_/Q _14189_/Y _14025_/A vssd1 vssd1 vccd1 vccd1 _14193_/C
+ sky130_fd_sc_hd__o22a_1
XFILLER_109_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10353_ _19862_/Q _10353_/B vssd1 vssd1 vccd1 vccd1 _10353_/Y sky130_fd_sc_hd__nor2_1
X_13141_ _19180_/Q vssd1 vssd1 vccd1 vccd1 _16645_/A sky130_fd_sc_hd__inv_2
XANTENNA__10264__A _19646_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11079__B _15858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13072_ _13072_/A _13193_/A vssd1 vssd1 vccd1 vccd1 _13073_/B sky130_fd_sc_hd__or2_2
Xclkbuf_leaf_120_HCLK clkbuf_4_4_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19595_/CLK sky130_fd_sc_hd__clkbuf_16
X_10284_ _10758_/B vssd1 vssd1 vccd1 vccd1 _10286_/A sky130_fd_sc_hd__inv_2
XANTENNA__18668__SET_B repeater222/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16900_ _17473_/A0 _16709_/Y _17512_/S vssd1 vssd1 vccd1 vccd1 _16900_/X sky130_fd_sc_hd__mux2_1
X_12023_ _12043_/A vssd1 vssd1 vccd1 vccd1 _12023_/X sky130_fd_sc_hd__clkbuf_2
X_17880_ _16078_/Y _16079_/Y _16080_/Y _16081_/Y _17913_/S0 _19632_/Q vssd1 vssd1
+ vccd1 vccd1 _17880_/X sky130_fd_sc_hd__mux4_2
XFILLER_104_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16831_ _16830_/X _19968_/Q _17488_/S vssd1 vssd1 vccd1 vccd1 _16831_/X sky130_fd_sc_hd__mux2_1
XFILLER_66_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17481__S _17529_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19550_ _19561_/CLK _19550_/D repeater269/X vssd1 vssd1 vccd1 vccd1 _19550_/Q sky130_fd_sc_hd__dfrtp_1
X_16762_ vssd1 vssd1 vccd1 vccd1 _16762_/HI _16762_/LO sky130_fd_sc_hd__conb_1
XFILLER_219_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12287__B1 _12028_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13974_ _18700_/Q vssd1 vssd1 vccd1 vccd1 _14030_/A sky130_fd_sc_hd__inv_2
XFILLER_18_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_108_HCLK_A clkbuf_4_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_234_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18501_ _19795_/CLK _18501_/D repeater219/X vssd1 vssd1 vccd1 vccd1 _18501_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_219_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15713_ _15713_/A _15713_/B vssd1 vssd1 vccd1 vccd1 _18648_/D sky130_fd_sc_hd__nor2_1
XFILLER_18_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19481_ _19506_/CLK hold170/X repeater256/X vssd1 vssd1 vccd1 vccd1 _19481_/Q sky130_fd_sc_hd__dfrtp_1
X_12925_ _19288_/Q vssd1 vssd1 vccd1 vccd1 _12925_/Y sky130_fd_sc_hd__inv_2
X_16693_ _19051_/Q vssd1 vssd1 vccd1 vccd1 _16693_/Y sky130_fd_sc_hd__inv_2
XFILLER_234_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18432_ _18435_/CLK _18432_/D vssd1 vssd1 vccd1 vccd1 _18432_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15644_ _15641_/Y _15642_/Y _15643_/X vssd1 vssd1 vccd1 vccd1 _15644_/X sky130_fd_sc_hd__o21a_1
XANTENNA__12039__B1 _12038_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19548__RESET_B hold346/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12856_ _18922_/Q vssd1 vssd1 vccd1 vccd1 _12859_/A sky130_fd_sc_hd__inv_2
XFILLER_222_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18363_ _18795_/CLK _18363_/D vssd1 vssd1 vccd1 vccd1 _18363_/Q sky130_fd_sc_hd__dfxtp_1
X_11807_ _11821_/A vssd1 vssd1 vccd1 vccd1 _11807_/X sky130_fd_sc_hd__clkbuf_2
X_15575_ _19437_/Q vssd1 vssd1 vccd1 vccd1 _15702_/A sky130_fd_sc_hd__inv_2
X_12787_ _18819_/Q vssd1 vssd1 vccd1 vccd1 _13542_/A sky130_fd_sc_hd__inv_2
XPHY_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16825__S _17522_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17314_ _16416_/Y _17844_/X _17568_/S vssd1 vssd1 vccd1 vccd1 _17314_/X sky130_fd_sc_hd__mux2_1
XFILLER_187_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14526_ _18324_/Q _14519_/A _14513_/X _14520_/A vssd1 vssd1 vccd1 vccd1 _18324_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09012__B _11996_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_230_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11738_ _11738_/A vssd1 vssd1 vccd1 vccd1 _11738_/X sky130_fd_sc_hd__clkbuf_4
X_18294_ _19847_/CLK _18294_/D vssd1 vssd1 vccd1 vccd1 _18294_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17245_ _17244_/X _18821_/Q _17386_/S vssd1 vssd1 vccd1 vccd1 _17245_/X sky130_fd_sc_hd__mux2_2
X_14457_ _18366_/Q _14451_/X _14415_/X _14453_/X vssd1 vssd1 vccd1 vccd1 _18366_/D
+ sky130_fd_sc_hd__a22o_1
X_11669_ _11669_/A vssd1 vssd1 vccd1 vccd1 _11669_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__16126__A _19717_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13408_ _20092_/Q _13483_/C _13406_/Y _18842_/Q _13407_/X vssd1 vssd1 vccd1 vccd1
+ _13417_/B sky130_fd_sc_hd__o221a_1
XANTENNA__12211__B1 _12104_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17176_ _17486_/A0 _13111_/Y _17543_/S vssd1 vssd1 vccd1 vccd1 _17176_/X sky130_fd_sc_hd__mux2_1
X_14388_ _18404_/Q _14381_/A _12729_/X _14382_/A vssd1 vssd1 vccd1 vccd1 _18404_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_6_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16127_ _19696_/Q vssd1 vssd1 vccd1 vccd1 _16127_/Y sky130_fd_sc_hd__inv_2
X_13339_ _13430_/A _13456_/A vssd1 vssd1 vccd1 vccd1 _13340_/B sky130_fd_sc_hd__or2_2
XANTENNA__17150__A0 _15963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_227_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16058_ _15335_/Y _16049_/X _16050_/Y _15836_/A _16057_/X vssd1 vssd1 vccd1 vccd1
+ _16058_/X sky130_fd_sc_hd__o221a_2
XFILLER_143_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15009_ _15058_/A _15094_/B _15009_/C vssd1 vssd1 vccd1 vccd1 _15011_/A sky130_fd_sc_hd__or3_4
XFILLER_97_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17453__A1 _12922_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19817_ _19822_/CLK _19817_/D repeater228/X vssd1 vssd1 vccd1 vccd1 _19817_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_57_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17391__S _17459_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16661__C1 _16660_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12278__B1 _12095_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19748_ _20070_/CLK _19748_/D repeater205/X vssd1 vssd1 vccd1 vccd1 _19748_/Q sky130_fd_sc_hd__dfrtp_1
X_09501_ _19313_/Q vssd1 vssd1 vccd1 vccd1 _09501_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19971__RESET_B repeater241/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19679_ _19772_/CLK _19679_/D repeater218/X vssd1 vssd1 vccd1 vccd1 _19679_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_37_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09432_ _19933_/Q vssd1 vssd1 vccd1 vccd1 _10009_/B sky130_fd_sc_hd__inv_2
XFILLER_52_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19900__RESET_B repeater195/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09363_ _20014_/Q vssd1 vssd1 vccd1 vccd1 _09474_/A sky130_fd_sc_hd__inv_2
XFILLER_178_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_240_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09294_ _09294_/A vssd1 vssd1 vccd1 vccd1 _09294_/X sky130_fd_sc_hd__buf_1
XFILLER_21_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_177_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_193_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12202__B1 _12088_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_143_HCLK clkbuf_4_1_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _18412_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_21_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17566__S _17566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17141__A0 _15768_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18853__RESET_B repeater231/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16495__A2 _16687_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_236_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10971_ _10243_/Y _10955_/Y _10968_/Y _19668_/Q _10970_/X vssd1 vssd1 vccd1 vccd1
+ _19668_/D sky130_fd_sc_hd__a32o_1
XFILLER_16_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_204_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12710_ _12710_/A vssd1 vssd1 vccd1 vccd1 _12711_/A sky130_fd_sc_hd__inv_2
XFILLER_244_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19641__RESET_B repeater261/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13690_ _18768_/Q _13685_/X _13680_/X _13686_/Y vssd1 vssd1 vccd1 vccd1 _18768_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_243_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12641_ _19005_/Q _12636_/X _12030_/A _12637_/X vssd1 vssd1 vccd1 vccd1 _19005_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15360_ _15364_/A _17589_/X vssd1 vssd1 vccd1 vccd1 _18501_/D sky130_fd_sc_hd__and2_1
XPHY_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12572_ _19050_/Q _12569_/X _12392_/X _12570_/X vssd1 vssd1 vccd1 vccd1 _19050_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18140__CLK _19851_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14311_ _18444_/Q _14304_/A _13678_/X _14305_/A vssd1 vssd1 vccd1 vccd1 _18444_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11523_ _11523_/A vssd1 vssd1 vccd1 vccd1 _11523_/X sky130_fd_sc_hd__clkbuf_4
XPHY_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15291_ _15389_/B _15285_/A _18630_/Q _15290_/Y vssd1 vssd1 vccd1 vccd1 _18630_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_178_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17030_ _17029_/X _19217_/Q _17545_/S vssd1 vssd1 vccd1 vccd1 _17030_/X sky130_fd_sc_hd__mux2_1
X_14242_ _18665_/Q _14236_/A _18505_/Q _14235_/A vssd1 vssd1 vccd1 vccd1 _18665_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11454_ _19561_/Q _11452_/Y _11453_/Y _19157_/Q vssd1 vssd1 vccd1 vccd1 _11454_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_194_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10405_ _19849_/Q _10404_/Y _10396_/A vssd1 vssd1 vccd1 vccd1 _19849_/D sky130_fd_sc_hd__o21a_1
XANTENNA__17476__S _17518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14173_ _19111_/Q vssd1 vssd1 vccd1 vccd1 _14173_/Y sky130_fd_sc_hd__inv_2
X_11385_ _19568_/Q vssd1 vssd1 vccd1 vccd1 _11581_/A sky130_fd_sc_hd__inv_2
XFILLER_180_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13124_ _19178_/Q vssd1 vssd1 vccd1 vccd1 _16618_/A sky130_fd_sc_hd__inv_2
XFILLER_124_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10336_ _10354_/A _10336_/B vssd1 vssd1 vccd1 vccd1 _10336_/X sky130_fd_sc_hd__and2_1
X_18981_ _19597_/CLK _18981_/D hold273/X vssd1 vssd1 vccd1 vccd1 _18981_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_3_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10267_ _19648_/Q vssd1 vssd1 vccd1 vccd1 _10267_/Y sky130_fd_sc_hd__inv_2
X_13055_ _18891_/Q vssd1 vssd1 vccd1 vccd1 _13064_/A sky130_fd_sc_hd__inv_2
X_17932_ _20036_/CLK _17932_/D vssd1 vssd1 vccd1 vccd1 _17932_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_repeater208_A repeater210/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12006_ _19360_/Q _12000_/X hold288/X _12003_/X vssd1 vssd1 vccd1 vccd1 _19360_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_79_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17863_ _16264_/Y _16265_/Y _16266_/Y _16267_/Y _17913_/S0 _19632_/Q vssd1 vssd1
+ vccd1 vccd1 _17863_/X sky130_fd_sc_hd__mux4_2
X_10198_ _19835_/Q vssd1 vssd1 vccd1 vccd1 _10198_/Y sky130_fd_sc_hd__inv_2
XFILLER_238_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19602_ _19610_/CLK _19602_/D hold343/X vssd1 vssd1 vccd1 vccd1 _19602_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_213_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16814_ _16813_/X _14039_/Y _17490_/S vssd1 vssd1 vccd1 vccd1 _16814_/X sky130_fd_sc_hd__mux2_2
XANTENNA__19729__RESET_B repeater207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17794_ _17790_/X _17791_/X _17792_/X _17793_/X _19647_/Q _19648_/Q vssd1 vssd1 vccd1
+ vccd1 _17794_/X sky130_fd_sc_hd__mux4_2
XFILLER_47_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19533_ _19540_/CLK _19533_/D repeater221/X vssd1 vssd1 vccd1 vccd1 _19533_/Q sky130_fd_sc_hd__dfrtp_4
Xclkbuf_leaf_24_HCLK clkbuf_4_9_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20051_/CLK sky130_fd_sc_hd__clkbuf_16
X_16745_ _16023_/Y _19640_/Q _15935_/Y _19627_/Q vssd1 vssd1 vccd1 vccd1 _16745_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_35_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13957_ _13957_/A vssd1 vssd1 vccd1 vccd1 _13957_/Y sky130_fd_sc_hd__inv_2
XFILLER_234_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19464_ _19470_/CLK _19464_/D repeater273/X vssd1 vssd1 vccd1 vccd1 _19464_/Q sky130_fd_sc_hd__dfrtp_1
X_12908_ _12908_/A _12908_/B _12908_/C _12908_/D vssd1 vssd1 vccd1 vccd1 _12956_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__19382__RESET_B repeater230/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09140__A3 hold344/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12680__B1 hold301/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16676_ _17072_/X _16594_/X _17030_/X _16595_/X vssd1 vssd1 vccd1 vccd1 _16678_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13209__C1 _13202_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13888_ _19211_/Q vssd1 vssd1 vccd1 vccd1 _13888_/Y sky130_fd_sc_hd__inv_2
XFILLER_234_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09023__A hold289/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15627_ _15666_/A _15627_/B vssd1 vssd1 vccd1 vccd1 _15627_/Y sky130_fd_sc_hd__nor2_1
X_18415_ _19849_/CLK _18415_/D vssd1 vssd1 vccd1 vccd1 _18415_/Q sky130_fd_sc_hd__dfxtp_1
X_19395_ _19933_/CLK _19395_/D repeater236/X vssd1 vssd1 vccd1 vccd1 _19395_/Q sky130_fd_sc_hd__dfrtp_4
X_12839_ _18946_/Q vssd1 vssd1 vccd1 vccd1 _12888_/B sky130_fd_sc_hd__inv_2
XANTENNA__09428__B2 _09424_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_222_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18346_ _19630_/CLK _18346_/D vssd1 vssd1 vccd1 vccd1 _18346_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11235__B2 _19021_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15558_ _15556_/Y _15557_/Y _15542_/X vssd1 vssd1 vccd1 vccd1 _15558_/X sky130_fd_sc_hd__o21a_1
XANTENNA__12432__B1 _12234_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14509_ hold325/X vssd1 vssd1 vccd1 vccd1 _14509_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_174_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18277_ _18435_/CLK _18277_/D vssd1 vssd1 vccd1 vccd1 _18277_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12384__A hold279/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15489_ _18567_/Q vssd1 vssd1 vccd1 vccd1 _15491_/A sky130_fd_sc_hd__inv_2
XFILLER_174_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17228_ _17486_/A0 _16485_/Y _17517_/S vssd1 vssd1 vccd1 vccd1 _17228_/X sky130_fd_sc_hd__mux2_1
Xinput30 input30/A vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__buf_1
Xinput41 input41/A vssd1 vssd1 vccd1 vccd1 input41/X sky130_fd_sc_hd__buf_1
Xinput52 input52/A vssd1 vssd1 vccd1 vccd1 input52/X sky130_fd_sc_hd__clkbuf_4
Xinput63 input63/A vssd1 vssd1 vccd1 vccd1 input63/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17386__S _17386_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput74 RsRx_S1 vssd1 vssd1 vccd1 vccd1 input74/X sky130_fd_sc_hd__clkbuf_4
X_17159_ _15963_/X _09547_/Y _17534_/S vssd1 vssd1 vccd1 vccd1 _17159_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10746__B1 _10451_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09981_ _09981_/A vssd1 vssd1 vccd1 vccd1 _09981_/Y sky130_fd_sc_hd__inv_2
XFILLER_170_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15845__D _15845_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08932_ _08927_/Y _18787_/Q _19867_/Q _08928_/Y _08931_/X vssd1 vssd1 vccd1 vccd1
+ _08970_/B sky130_fd_sc_hd__o221a_1
XFILLER_69_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_218_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12559__A _12598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_154_HCLK_A clkbuf_4_1_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09415_ _10040_/A _19384_/Q _19924_/Q _09414_/Y vssd1 vssd1 vccd1 vccd1 _09416_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_13_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10079__A _10079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09346_ _20031_/Q vssd1 vssd1 vccd1 vccd1 _09491_/A sky130_fd_sc_hd__inv_2
XFILLER_40_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12423__B1 _12356_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09277_ _20052_/Q _09270_/A _09101_/X _09271_/A vssd1 vssd1 vccd1 vccd1 _20052_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_138_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold203_A HADDR[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17296__S _17542_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11170_ _19625_/Q _11170_/B vssd1 vssd1 vccd1 vccd1 _11170_/X sky130_fd_sc_hd__or2_2
XFILLER_106_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10121_ _18571_/Q _18570_/Q _15498_/A vssd1 vssd1 vccd1 vccd1 _15509_/B sky130_fd_sc_hd__or3_4
XFILLER_164_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10052_ _19933_/Q _19932_/Q _10052_/C vssd1 vssd1 vccd1 vccd1 _10052_/X sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_47_HCLK clkbuf_opt_2_HCLK/A vssd1 vssd1 vccd1 vccd1 _18633_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_102_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19893__RESET_B repeater205/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14860_ _14860_/A vssd1 vssd1 vccd1 vccd1 _14860_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_235_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13811_ _18714_/Q vssd1 vssd1 vccd1 vccd1 _13951_/A sky130_fd_sc_hd__inv_2
XFILLER_17_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18506__CLK _18506_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input19_A HADDR[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14791_ _14791_/A vssd1 vssd1 vccd1 vccd1 _14791_/X sky130_fd_sc_hd__buf_2
XFILLER_180_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16530_ _16530_/A vssd1 vssd1 vccd1 vccd1 _16684_/A sky130_fd_sc_hd__buf_2
XFILLER_56_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13742_ _13737_/A _13259_/B _13259_/A vssd1 vssd1 vccd1 vccd1 _13742_/X sky130_fd_sc_hd__o21a_1
X_10954_ _10954_/A _10954_/B vssd1 vssd1 vccd1 vccd1 _10978_/A sky130_fd_sc_hd__or2_2
XFILLER_113_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16461_ _17051_/X _16494_/A _17311_/X _15999_/A vssd1 vssd1 vccd1 vccd1 _16461_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_188_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13673_ _18777_/Q _13671_/X _12602_/X _13672_/X vssd1 vssd1 vccd1 vccd1 _18777_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_13_HCLK_A clkbuf_4_2_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10885_ _14279_/A vssd1 vssd1 vccd1 vccd1 _10885_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_204_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18200_ _18216_/CLK _18200_/D vssd1 vssd1 vccd1 vccd1 _18200_/Q sky130_fd_sc_hd__dfxtp_1
X_15412_ _18538_/Q _13225_/B _13226_/B vssd1 vssd1 vccd1 vccd1 _15412_/X sky130_fd_sc_hd__a21bo_1
XFILLER_188_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_76_HCLK_A clkbuf_opt_4_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12624_ _19018_/Q _12622_/X _12389_/X _12623_/X vssd1 vssd1 vccd1 vccd1 _19018_/D
+ sky130_fd_sc_hd__a22o_1
X_19180_ _19293_/CLK _19180_/D repeater187/X vssd1 vssd1 vccd1 vccd1 _19180_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16392_ _17338_/X _16494_/A _17341_/X _15999_/A vssd1 vssd1 vccd1 vccd1 _16392_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_1_HCLK_A clkbuf_4_0_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19901__CLK _20123_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18131_ _18198_/CLK _18131_/D vssd1 vssd1 vccd1 vccd1 _18131_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15343_ _15347_/A _17597_/X vssd1 vssd1 vccd1 vccd1 _18493_/D sky130_fd_sc_hd__and2_1
XPHY_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12555_ _19058_/Q _12553_/Y _12556_/B _12554_/X vssd1 vssd1 vccd1 vccd1 _19058_/D
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10717__A _10842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_repeater158_A _17544_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11506_ _11523_/A vssd1 vssd1 vccd1 vccd1 _11506_/X sky130_fd_sc_hd__clkbuf_4
X_18062_ _18465_/CLK _18062_/D vssd1 vssd1 vccd1 vccd1 _18062_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15274_ _18640_/Q _18637_/Q _18636_/Q _15323_/A vssd1 vssd1 vccd1 vccd1 _15275_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_184_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12486_ _19093_/Q _12457_/A _12241_/X _12458_/A vssd1 vssd1 vccd1 vccd1 _19093_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18704__RESET_B repeater253/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17013_ _17012_/X _09724_/Y _17523_/S vssd1 vssd1 vccd1 vccd1 _17013_/X sky130_fd_sc_hd__mux2_1
XFILLER_184_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14225_ _18495_/Q _14225_/B vssd1 vssd1 vccd1 vccd1 _14226_/B sky130_fd_sc_hd__or2_1
XFILLER_208_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11437_ _11549_/A _19126_/Q _19560_/Q _11429_/Y _11436_/X vssd1 vssd1 vccd1 vccd1
+ _11437_/X sky130_fd_sc_hd__a221o_1
XFILLER_125_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10728__B1 _10423_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output87_A _16600_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14156_ _19109_/Q vssd1 vssd1 vccd1 vccd1 _14156_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11368_ _19550_/Q vssd1 vssd1 vccd1 vccd1 _11620_/A sky130_fd_sc_hd__inv_2
XFILLER_113_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13107_ _16718_/A _18916_/Q _19165_/Q _13067_/A vssd1 vssd1 vccd1 vccd1 _13107_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_140_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10319_ _10319_/A _13285_/A vssd1 vssd1 vccd1 vccd1 _10368_/A sky130_fd_sc_hd__or2_2
XANTENNA__18036__CLK _19851_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14087_ _19077_/Q vssd1 vssd1 vccd1 vccd1 _14087_/Y sky130_fd_sc_hd__inv_2
X_18964_ _19208_/CLK _18964_/D hold370/X vssd1 vssd1 vccd1 vccd1 _18964_/Q sky130_fd_sc_hd__dfrtp_4
X_11299_ _11261_/X _11299_/B _11299_/C _11299_/D vssd1 vssd1 vccd1 vccd1 _11299_/X
+ sky130_fd_sc_hd__and4b_1
XFILLER_224_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17915_ _18337_/Q _18217_/Q _18209_/Q _18201_/Q _17918_/S0 _18750_/Q vssd1 vssd1
+ vccd1 vccd1 _17915_/X sky130_fd_sc_hd__mux4_1
X_13038_ _18908_/Q vssd1 vssd1 vccd1 vccd1 _13080_/A sky130_fd_sc_hd__inv_2
X_18895_ _19352_/CLK _18895_/D hold372/X vssd1 vssd1 vccd1 vccd1 _18895_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_94_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17846_ _16351_/Y _16352_/Y _16353_/Y _16354_/Y _17908_/S0 _18759_/Q vssd1 vssd1
+ vccd1 vccd1 _17846_/X sky130_fd_sc_hd__mux4_2
XANTENNA__10900__B1 _10863_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19873__SET_B repeater261/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17777_ _18324_/Q _18004_/Q _18308_/Q _18300_/Q _17923_/S0 _19646_/Q vssd1 vssd1
+ vccd1 vccd1 _17777_/X sky130_fd_sc_hd__mux4_2
X_14989_ _18058_/Q _14978_/A _14782_/X _14979_/A vssd1 vssd1 vccd1 vccd1 _18058_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11283__A _19018_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19516_ _19867_/CLK hold215/X repeater262/X vssd1 vssd1 vccd1 vccd1 _19516_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__12653__B1 _12602_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16728_ _16728_/A _16728_/B _16728_/C _16728_/D vssd1 vssd1 vccd1 vccd1 _16728_/X
+ sky130_fd_sc_hd__or4_4
XFILLER_81_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16659_ _19048_/Q vssd1 vssd1 vccd1 vccd1 _16659_/Y sky130_fd_sc_hd__inv_2
X_19447_ _20058_/CLK _19447_/D repeater194/X vssd1 vssd1 vccd1 vccd1 _19447_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_23_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16395__B2 _16394_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09200_ _13283_/B _09198_/A _09205_/B vssd1 vssd1 vccd1 vccd1 _09200_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__12405__B1 _12404_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19378_ _19937_/CLK _19378_/D repeater230/X vssd1 vssd1 vccd1 vccd1 _19378_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_176_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09131_ _09131_/A _09136_/B vssd1 vssd1 vccd1 vccd1 _09131_/X sky130_fd_sc_hd__or2_1
X_18329_ _19637_/CLK _18329_/D vssd1 vssd1 vccd1 vccd1 _18329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09062_ _20105_/Q _09053_/X _09061_/X _09055_/X vssd1 vssd1 vccd1 vccd1 _20105_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_191_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16314__A _19770_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09964_ _09968_/A vssd1 vssd1 vccd1 vccd1 _09964_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_134_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14330__B1 _14329_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08915_ _20124_/Q vssd1 vssd1 vccd1 vccd1 _10132_/B sky130_fd_sc_hd__inv_2
X_20084_ _20085_/CLK _20084_/D repeater204/X vssd1 vssd1 vccd1 vccd1 _20084_/Q sky130_fd_sc_hd__dfrtp_1
X_09895_ _09895_/A _09895_/B _09895_/C _09895_/D vssd1 vssd1 vccd1 vccd1 _09948_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_100_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14397__B1 _14351_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_213_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10670_ _10677_/A vssd1 vssd1 vccd1 vccd1 _10670_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_213_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_179_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16208__B _16212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09329_ _09329_/A _09329_/B vssd1 vssd1 vccd1 vccd1 _15724_/A sky130_fd_sc_hd__or2_1
XFILLER_139_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16923__S _17413_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12340_ _19175_/Q _12334_/X _12104_/X _12335_/X vssd1 vssd1 vccd1 vccd1 _19175_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_216_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12271_ _19219_/Q _12269_/X _12083_/X _12270_/X vssd1 vssd1 vccd1 vccd1 _19219_/D
+ sky130_fd_sc_hd__a22o_1
X_14010_ _14010_/A _14139_/A vssd1 vssd1 vccd1 vccd1 _14011_/B sky130_fd_sc_hd__or2_2
XFILLER_153_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11222_ _19599_/Q _11217_/Y _19578_/Q _11218_/Y _11221_/X vssd1 vssd1 vccd1 vccd1
+ _11223_/D sky130_fd_sc_hd__o221a_1
X_11153_ _19627_/Q vssd1 vssd1 vccd1 vccd1 _11153_/Y sky130_fd_sc_hd__inv_2
XFILLER_122_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10104_ _10104_/A vssd1 vssd1 vccd1 vccd1 _10107_/A sky130_fd_sc_hd__inv_2
XANTENNA__14321__B1 _14273_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11084_ _19059_/Q vssd1 vssd1 vccd1 vccd1 _11085_/C sky130_fd_sc_hd__inv_2
X_15961_ _15961_/A vssd1 vssd1 vccd1 vccd1 _16436_/B sky130_fd_sc_hd__buf_1
XFILLER_49_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17700_ _19818_/Q _19760_/Q _18548_/Q vssd1 vssd1 vccd1 vccd1 _17700_/X sky130_fd_sc_hd__mux2_1
X_10035_ _10035_/A _10077_/A vssd1 vssd1 vccd1 vccd1 _10036_/B sky130_fd_sc_hd__or2_2
X_14912_ _18104_/Q _14908_/X _14703_/X _14910_/X vssd1 vssd1 vccd1 vccd1 _18104_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_248_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18680_ _18686_/CLK _18680_/D hold359/X vssd1 vssd1 vccd1 vccd1 _18680_/Q sky130_fd_sc_hd__dfrtp_1
X_15892_ _17550_/X vssd1 vssd1 vccd1 vccd1 _15892_/Y sky130_fd_sc_hd__inv_2
XFILLER_209_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14843_ _18146_/Q _14833_/A _14842_/X _14834_/A vssd1 vssd1 vccd1 vccd1 _18146_/D
+ sky130_fd_sc_hd__a22o_1
X_17631_ _19878_/Q _15717_/Y _17631_/S vssd1 vssd1 vccd1 vccd1 _17631_/X sky130_fd_sc_hd__mux2_1
XFILLER_48_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output125_A _15777_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17562_ _17561_/X _13289_/Y _17567_/S vssd1 vssd1 vccd1 vccd1 _17562_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12635__B1 _12410_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14774_ _18185_/Q _14771_/X _14745_/X _14773_/X vssd1 vssd1 vccd1 vccd1 _18185_/D
+ sky130_fd_sc_hd__a22o_1
X_11986_ _19367_/Q _11955_/A _11924_/X _11956_/A vssd1 vssd1 vccd1 vccd1 _19367_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_44_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16513_ _16513_/A vssd1 vssd1 vccd1 vccd1 _16513_/X sky130_fd_sc_hd__buf_2
X_19301_ _19952_/CLK _19301_/D repeater242/X vssd1 vssd1 vccd1 vccd1 _19301_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_216_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13725_ _13725_/A vssd1 vssd1 vccd1 vccd1 _13733_/A sky130_fd_sc_hd__buf_1
X_10937_ _10937_/A vssd1 vssd1 vccd1 vccd1 _19672_/D sky130_fd_sc_hd__inv_2
X_17493_ _17492_/X _11351_/Y _17493_/S vssd1 vssd1 vccd1 vccd1 _17493_/X sky130_fd_sc_hd__mux2_1
XANTENNA__18956__RESET_B repeater257/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_231_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16444_ _18478_/Q vssd1 vssd1 vccd1 vccd1 _16444_/Y sky130_fd_sc_hd__inv_2
X_19232_ _19314_/CLK _19232_/D repeater214/X vssd1 vssd1 vccd1 vccd1 _19232_/Q sky130_fd_sc_hd__dfrtp_4
X_13656_ _13671_/A vssd1 vssd1 vccd1 vccd1 _13656_/X sky130_fd_sc_hd__clkbuf_2
X_10868_ _12238_/A vssd1 vssd1 vccd1 vccd1 _10868_/X sky130_fd_sc_hd__buf_2
XFILLER_231_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12607_ _19026_/Q _12576_/A _12541_/X _12577_/A vssd1 vssd1 vccd1 vccd1 _19026_/D
+ sky130_fd_sc_hd__a22o_1
X_19163_ _19214_/CLK _19163_/D hold367/X vssd1 vssd1 vccd1 vccd1 _19163_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16375_ _19715_/Q vssd1 vssd1 vccd1 vccd1 _16375_/Y sky130_fd_sc_hd__inv_2
XPHY_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13587_ _18819_/Q _13586_/Y _13574_/X _13543_/B vssd1 vssd1 vccd1 vccd1 _18819_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_185_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16833__S _17385_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10799_ _19738_/Q _10794_/B _18653_/Q vssd1 vssd1 vccd1 vccd1 _10800_/B sky130_fd_sc_hd__o21ai_1
XFILLER_219_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18114_ _19435_/CLK _18114_/D vssd1 vssd1 vccd1 vccd1 _18114_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15326_ _15326_/A vssd1 vssd1 vccd1 vccd1 _15326_/Y sky130_fd_sc_hd__inv_2
XFILLER_185_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19094_ _19609_/CLK _19094_/D hold359/X vssd1 vssd1 vccd1 vccd1 _19094_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_8_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12538_ _13678_/A vssd1 vssd1 vccd1 vccd1 _12538_/X sky130_fd_sc_hd__buf_4
XFILLER_157_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18045_ _18959_/CLK _18045_/D vssd1 vssd1 vccd1 vccd1 _18045_/Q sky130_fd_sc_hd__dfxtp_1
X_15257_ _15268_/C vssd1 vssd1 vccd1 vccd1 _15257_/Y sky130_fd_sc_hd__inv_2
XFILLER_184_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12469_ _19106_/Q _12464_/X hold256/X _12465_/X vssd1 vssd1 vccd1 vccd1 _19106_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12662__A _12698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14208_ _19119_/Q _14028_/A _19098_/Q _14008_/A vssd1 vssd1 vccd1 vccd1 _14208_/X
+ sky130_fd_sc_hd__o22a_1
X_15188_ _17931_/Q _14251_/A _10715_/X _14252_/A vssd1 vssd1 vccd1 vccd1 _17931_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_125_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14139_ _14139_/A vssd1 vssd1 vccd1 vccd1 _14139_/Y sky130_fd_sc_hd__clkinv_1
XFILLER_113_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19744__RESET_B repeater207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19996_ _19997_/CLK _19996_/D repeater192/X vssd1 vssd1 vccd1 vccd1 _19996_/Q sky130_fd_sc_hd__dfrtp_1
X_18947_ _18947_/CLK _18947_/D repeater211/X vssd1 vssd1 vccd1 vccd1 _18947_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_79_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09680_ _19401_/Q vssd1 vssd1 vccd1 vccd1 _09680_/Y sky130_fd_sc_hd__inv_2
X_18878_ _20048_/CLK _18878_/D repeater208/X vssd1 vssd1 vccd1 vccd1 _18878_/Q sky130_fd_sc_hd__dfrtp_1
X_17829_ _17825_/X _17826_/X _17827_/X _17828_/X _18751_/Q _18752_/Q vssd1 vssd1 vccd1
+ vccd1 _17829_/X sky130_fd_sc_hd__mux4_2
XFILLER_94_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12626__B1 _12394_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18697__RESET_B hold351/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17317__A0 _17473_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09114_ _20086_/Q vssd1 vssd1 vccd1 vccd1 _09138_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__15867__B _15867_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09045_ hold301/X vssd1 vssd1 vccd1 vccd1 hold300/A sky130_fd_sc_hd__buf_4
XANTENNA__16540__A1 _17152_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11365__B1 _19610_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17574__S _17584_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15883__A _15883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19485__RESET_B repeater260/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16698__B _16698_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09947_ _09947_/A _09947_/B _09947_/C _09947_/D vssd1 vssd1 vccd1 vccd1 _09948_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_131_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19414__RESET_B repeater210/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_219_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20067_ _20124_/CLK _20067_/D repeater207/X vssd1 vssd1 vccd1 vccd1 _20067_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_218_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09878_ _09878_/A vssd1 vssd1 vccd1 vccd1 _09878_/Y sky130_fd_sc_hd__inv_2
XANTENNA__10820__A _12257_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16918__S _17529_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater280 hold358/A vssd1 vssd1 vccd1 vccd1 hold360/A sky130_fd_sc_hd__buf_8
XFILLER_72_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11840_ _10147_/X _15643_/A _11840_/S vssd1 vssd1 vccd1 vccd1 _19437_/D sky130_fd_sc_hd__mux2_1
XPHY_4434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12617__B1 _12375_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11771_ _11771_/A vssd1 vssd1 vccd1 vccd1 _11771_/X sky130_fd_sc_hd__clkbuf_2
XPHY_4489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13510_ _18762_/Q vssd1 vssd1 vccd1 vccd1 _14628_/B sky130_fd_sc_hd__clkbuf_2
XPHY_3766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10722_ _10722_/A vssd1 vssd1 vccd1 vccd1 _10722_/X sky130_fd_sc_hd__buf_1
XFILLER_54_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11840__A1 _15643_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14490_ _14490_/A _14963_/B _15094_/C vssd1 vssd1 vccd1 vccd1 _14492_/A sky130_fd_sc_hd__or3_4
XFILLER_213_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13441_ _13433_/B _13348_/B _13439_/Y _13489_/C vssd1 vssd1 vccd1 vccd1 _18861_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_201_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10653_ _19793_/Q _10653_/B vssd1 vssd1 vccd1 vccd1 _10654_/B sky130_fd_sc_hd__or2_1
XFILLER_13_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10267__A _19648_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16160_ _18166_/Q vssd1 vssd1 vccd1 vccd1 _16160_/Y sky130_fd_sc_hd__inv_2
X_13372_ _13360_/X _13372_/B _13372_/C _13372_/D vssd1 vssd1 vccd1 vccd1 _13418_/A
+ sky130_fd_sc_hd__and4b_1
XANTENNA__14790__B1 _14751_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10584_ _10614_/A _15297_/B _10584_/C _10584_/D vssd1 vssd1 vccd1 vccd1 _10584_/X
+ sky130_fd_sc_hd__and4bb_1
XFILLER_154_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15111_ _15111_/A vssd1 vssd1 vccd1 vccd1 _15112_/A sky130_fd_sc_hd__inv_2
X_12323_ _19188_/Q _12318_/X _12074_/X _12321_/X vssd1 vssd1 vccd1 vccd1 _19188_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_186_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16091_ _18405_/Q vssd1 vssd1 vccd1 vccd1 _16091_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15042_ _18029_/Q _15035_/X _15002_/X _15037_/X vssd1 vssd1 vccd1 vccd1 _18029_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14542__B1 hold334/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12254_ _10954_/B _12253_/X _12252_/S vssd1 vssd1 vccd1 vccd1 _12254_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_123_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17484__S _17535_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11205_ _19022_/Q vssd1 vssd1 vccd1 vccd1 _11205_/Y sky130_fd_sc_hd__inv_2
X_19850_ _19851_/CLK _19850_/D repeater258/X vssd1 vssd1 vccd1 vccd1 _19850_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_123_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12185_ _12187_/A _12372_/A vssd1 vssd1 vccd1 vccd1 _12186_/S sky130_fd_sc_hd__or2_1
XANTENNA__18844__CLK _18866_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18801_ _19900_/CLK _18801_/D repeater199/X vssd1 vssd1 vccd1 vccd1 _18801_/Q sky130_fd_sc_hd__dfrtp_2
X_11136_ _19225_/Q vssd1 vssd1 vccd1 vccd1 _12708_/B sky130_fd_sc_hd__inv_2
X_19781_ _20057_/CLK _19781_/D repeater202/X vssd1 vssd1 vccd1 vccd1 _19781_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_205_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16993_ _15768_/Y _14189_/Y _17546_/S vssd1 vssd1 vccd1 vccd1 _16993_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18732_ _19224_/CLK _18732_/D repeater186/X vssd1 vssd1 vccd1 vccd1 _18732_/Q sky130_fd_sc_hd__dfrtp_1
X_11067_ _11061_/X _11066_/B _15058_/A _19851_/Q _11123_/B vssd1 vssd1 vccd1 vccd1
+ _11067_/X sky130_fd_sc_hd__a32o_1
XFILLER_95_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15944_ _18267_/Q vssd1 vssd1 vccd1 vccd1 _15944_/Y sky130_fd_sc_hd__inv_2
XFILLER_237_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10018_ _10040_/A _10039_/A _10041_/A _10038_/A vssd1 vssd1 vccd1 vccd1 _10019_/D
+ sky130_fd_sc_hd__or4_4
XFILLER_237_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18663_ _20064_/CLK _18663_/D repeater198/X vssd1 vssd1 vccd1 vccd1 _18663_/Q sky130_fd_sc_hd__dfrtp_1
X_15875_ _19365_/Q _15878_/B vssd1 vssd1 vccd1 vccd1 _15875_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__16828__S _17385_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17614_ _15201_/X _15201_/B _17614_/S vssd1 vssd1 vccd1 vccd1 _17614_/X sky130_fd_sc_hd__mux2_1
X_14826_ _18158_/Q _14820_/X _14791_/X _14822_/X vssd1 vssd1 vccd1 vccd1 _18158_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_224_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17890__S0 _17913_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12608__B1 _12543_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18594_ _19855_/CLK _18594_/D repeater265/X vssd1 vssd1 vccd1 vccd1 _18594_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_224_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14757_ _18194_/Q _14746_/A _14693_/X _14747_/A vssd1 vssd1 vccd1 vccd1 _18194_/D
+ sky130_fd_sc_hd__a22o_1
X_17545_ _17544_/X _13863_/Y _17545_/S vssd1 vssd1 vccd1 vccd1 _17545_/X sky130_fd_sc_hd__mux2_2
X_11969_ _11977_/A vssd1 vssd1 vccd1 vccd1 _11969_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_44_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18790__RESET_B repeater261/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10095__B1 _10026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13708_ _18761_/Q vssd1 vssd1 vccd1 vccd1 _13708_/Y sky130_fd_sc_hd__inv_2
X_17476_ _17475_/X _15450_/A _17518_/S vssd1 vssd1 vccd1 vccd1 _17476_/X sky130_fd_sc_hd__mux2_1
X_14688_ _18230_/Q _14682_/X _14578_/X _14684_/X vssd1 vssd1 vccd1 vccd1 _18230_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_60_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19215_ _19221_/CLK _19215_/D hold365/X vssd1 vssd1 vccd1 vccd1 _19215_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__15968__A _19686_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13639_ _18797_/Q _13637_/Y _13637_/B _13638_/X vssd1 vssd1 vccd1 vccd1 _18797_/D
+ sky130_fd_sc_hd__o22a_1
X_16427_ _18265_/Q vssd1 vssd1 vccd1 vccd1 _16427_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13584__A1 _18821_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19146_ _19597_/CLK _19146_/D repeater281/X vssd1 vssd1 vccd1 vccd1 _19146_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__14781__B1 _14780_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16358_ _17983_/Q vssd1 vssd1 vccd1 vccd1 _16358_/Y sky130_fd_sc_hd__inv_2
XFILLER_173_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19996__RESET_B repeater192/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15309_ _18628_/Q vssd1 vssd1 vccd1 vccd1 _15309_/Y sky130_fd_sc_hd__inv_2
XFILLER_145_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12392__A hold308/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19077_ _19609_/CLK _19077_/D hold343/X vssd1 vssd1 vccd1 vccd1 _19077_/Q sky130_fd_sc_hd__dfrtp_1
X_16289_ _18103_/Q vssd1 vssd1 vccd1 vccd1 _16289_/Y sky130_fd_sc_hd__inv_2
X_18028_ _19510_/CLK _18028_/D vssd1 vssd1 vccd1 vccd1 _18028_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17394__S _19498_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09801_ _19979_/Q _09800_/Y _09731_/A _09792_/B vssd1 vssd1 vccd1 vccd1 _19979_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_141_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19979_ _19992_/CLK _19979_/D repeater192/X vssd1 vssd1 vccd1 vccd1 _19979_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_115_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09732_ _20003_/Q _09738_/A _09670_/Y _09669_/A _09731_/X vssd1 vssd1 vccd1 vccd1
+ _20003_/D sky130_fd_sc_hd__o221a_1
X_09663_ _19997_/Q vssd1 vssd1 vccd1 vccd1 _09753_/A sky130_fd_sc_hd__inv_2
XFILLER_83_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18878__RESET_B repeater208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_227_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09594_ _09480_/A _09480_/B _09592_/Y _09587_/X vssd1 vssd1 vccd1 vccd1 _20020_/D
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__17881__S0 _17913_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18807__RESET_B repeater231/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_opt_4_HCLK_A clkbuf_opt_4_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09028_ _20118_/Q _09015_/X _09027_/X _09019_/X vssd1 vssd1 vccd1 vccd1 _20118_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14524__B1 _14509_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold260 input68/X vssd1 vssd1 vccd1 vccd1 hold260/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold271 input41/X vssd1 vssd1 vccd1 vccd1 hold271/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 input43/X vssd1 vssd1 vccd1 vccd1 hold282/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold293 hold358/X vssd1 vssd1 vccd1 vccd1 hold357/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20119_ _20120_/CLK _20119_/D repeater234/X vssd1 vssd1 vccd1 vccd1 _20119_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_172_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13990_ _18684_/Q vssd1 vssd1 vccd1 vccd1 _14014_/A sky130_fd_sc_hd__inv_2
XFILLER_219_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12941_ _12941_/A _12941_/B _12941_/C _12941_/D vssd1 vssd1 vccd1 vccd1 _12956_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_46_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15660_ _15661_/A vssd1 vssd1 vccd1 vccd1 _15660_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17872__S0 _17913_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12872_ _13000_/A _12967_/A vssd1 vssd1 vccd1 vccd1 _12873_/B sky130_fd_sc_hd__or2_2
XPHY_4220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14611_ _18275_/Q _14601_/A _14567_/X _14602_/A vssd1 vssd1 vccd1 vccd1 _18275_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11823_ _19445_/Q _11821_/X _10882_/X _11822_/X vssd1 vssd1 vccd1 vccd1 _19445_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15591_ _15594_/B _15589_/X _15590_/X vssd1 vssd1 vccd1 vccd1 _15591_/X sky130_fd_sc_hd__o21a_1
XFILLER_45_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17330_ _17486_/A0 _13152_/Y _17543_/S vssd1 vssd1 vccd1 vccd1 _17330_/X sky130_fd_sc_hd__mux2_1
XPHY_4297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14542_ _18315_/Q _14532_/A hold334/X _14533_/A vssd1 vssd1 vccd1 vccd1 _18315_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_60_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11754_ hold153/X _11750_/X _19488_/Q _11751_/X vssd1 vssd1 vccd1 vccd1 hold155/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_230_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10705_ _15404_/A _10704_/B _10701_/Y _10702_/Y _10716_/S vssd1 vssd1 vccd1 vccd1
+ _10706_/A sky130_fd_sc_hd__o32a_1
X_17261_ _17486_/A0 _09942_/Y _17543_/S vssd1 vssd1 vccd1 vccd1 _17261_/X sky130_fd_sc_hd__mux2_1
XANTENNA__17479__S _17518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14473_ _18355_/Q _14464_/A hold334/X _14465_/A vssd1 vssd1 vccd1 vccd1 _18355_/D
+ sky130_fd_sc_hd__a22o_1
X_11685_ _19532_/Q _11669_/A _15270_/B _11666_/X vssd1 vssd1 vccd1 vccd1 _19532_/D
+ sky130_fd_sc_hd__o22a_1
XPHY_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16212_ _16212_/A _16212_/B vssd1 vssd1 vccd1 vccd1 _16212_/Y sky130_fd_sc_hd__nor2_1
X_19000_ _19585_/CLK _19000_/D hold363/X vssd1 vssd1 vccd1 vccd1 _19000_/Q sky130_fd_sc_hd__dfrtp_1
X_13424_ _13445_/A vssd1 vssd1 vccd1 vccd1 _13489_/C sky130_fd_sc_hd__buf_2
XANTENNA__12369__A2 _12334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10636_ _19799_/Q _10606_/A _10614_/B _10609_/X vssd1 vssd1 vccd1 vccd1 _19799_/D
+ sky130_fd_sc_hd__a22o_1
X_17192_ _17191_/X _11334_/Y _17493_/S vssd1 vssd1 vccd1 vccd1 _17192_/X sky130_fd_sc_hd__mux2_1
XANTENNA__14763__B1 _14749_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16143_ _16141_/Y _15884_/X _16142_/Y _15915_/X vssd1 vssd1 vccd1 vccd1 _16143_/X
+ sky130_fd_sc_hd__o22a_1
X_13355_ _13355_/A vssd1 vssd1 vccd1 vccd1 _13355_/Y sky130_fd_sc_hd__inv_2
X_10567_ _10583_/A _10939_/C _10567_/C _10567_/D vssd1 vssd1 vccd1 vccd1 _10613_/A
+ sky130_fd_sc_hd__nor4_2
XANTENNA_repeater238_A repeater239/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14515__B1 hold334/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12306_ _19195_/Q _12298_/X _12236_/X _12300_/X vssd1 vssd1 vccd1 vccd1 _19195_/D
+ sky130_fd_sc_hd__a22o_1
X_16074_ _17454_/X _15997_/X _17457_/X _15998_/X _16073_/X vssd1 vssd1 vccd1 vccd1
+ _16074_/X sky130_fd_sc_hd__o221a_2
XFILLER_182_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13286_ _13746_/A _15192_/B vssd1 vssd1 vccd1 vccd1 _13750_/A sky130_fd_sc_hd__nand2_1
X_10498_ _10732_/C _19542_/Q _10732_/B _10519_/D vssd1 vssd1 vccd1 vccd1 _11651_/A
+ sky130_fd_sc_hd__and4b_1
XFILLER_143_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15025_ _15025_/A vssd1 vssd1 vccd1 vccd1 _15025_/X sky130_fd_sc_hd__clkbuf_2
X_19902_ _20123_/CLK _19902_/D repeater195/X vssd1 vssd1 vccd1 vccd1 _19902_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_216_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12237_ _19229_/Q _12228_/X _12236_/X _12229_/X vssd1 vssd1 vccd1 vccd1 _19229_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_69_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19833_ _20058_/CLK _19833_/D repeater194/X vssd1 vssd1 vccd1 vccd1 _19833_/Q sky130_fd_sc_hd__dfrtp_4
X_12168_ _19271_/Q _12164_/X _11909_/X _12165_/X vssd1 vssd1 vccd1 vccd1 _19271_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_229_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11119_ _19635_/Q _11119_/B vssd1 vssd1 vccd1 vccd1 _11119_/X sky130_fd_sc_hd__or2_1
X_19764_ _19814_/CLK _19764_/D repeater223/X vssd1 vssd1 vccd1 vccd1 _19764_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_96_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12099_ _19314_/Q _12094_/X _12098_/X _12096_/X vssd1 vssd1 vccd1 vccd1 _19314_/D
+ sky130_fd_sc_hd__a22o_1
X_16976_ _16975_/X _19213_/Q _17545_/S vssd1 vssd1 vccd1 vccd1 _16976_/X sky130_fd_sc_hd__mux2_1
XFILLER_232_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18715_ _18718_/CLK _18715_/D repeater252/X vssd1 vssd1 vccd1 vccd1 _18715_/Q sky130_fd_sc_hd__dfrtp_1
Xinput6 input6/A vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_1
X_15927_ _18163_/Q vssd1 vssd1 vccd1 vccd1 _15927_/Y sky130_fd_sc_hd__inv_2
X_19695_ _20051_/CLK _19695_/D repeater208/X vssd1 vssd1 vccd1 vccd1 _19695_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_37_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17863__S0 _17913_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18646_ _20059_/CLK _18646_/D repeater197/X vssd1 vssd1 vccd1 vccd1 _18646_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_209_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15858_ _15858_/A _15858_/B _15858_/C _15858_/D vssd1 vssd1 vccd1 vccd1 _15859_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14809_ _18167_/Q _14801_/X _14808_/X _14804_/X vssd1 vssd1 vccd1 vccd1 _18167_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_91_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18577_ _19437_/CLK _18577_/D repeater273/X vssd1 vssd1 vccd1 vccd1 _18577_/Q sky130_fd_sc_hd__dfrtp_1
X_15789_ _18050_/Q vssd1 vssd1 vccd1 vccd1 _15789_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16991__A1 _19423_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_205_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17528_ _17527_/X _09521_/Y _17534_/S vssd1 vssd1 vccd1 vccd1 _17528_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17389__S _17544_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17459_ _17458_/X _11316_/Y _17459_/S vssd1 vssd1 vccd1 vccd1 _17459_/X sky130_fd_sc_hd__mux2_1
XFILLER_177_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17918__S1 _18750_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19129_ _19470_/CLK _19129_/D repeater274/X vssd1 vssd1 vccd1 vccd1 _19129_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_146_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14506__B1 _14437_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19006__RESET_B hold346/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11740__B1 _16931_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09715_ _09745_/A _19418_/Q _09789_/A _19406_/Q vssd1 vssd1 vccd1 vccd1 _09715_/X
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_80_HCLK clkbuf_4_13_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19325_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_28_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09646_ _09793_/A _09792_/A _09646_/C _09794_/A vssd1 vssd1 vccd1 vccd1 _09647_/D
+ sky130_fd_sc_hd__or4_4
XFILLER_216_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17854__S0 _19633_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09577_ _09577_/A vssd1 vssd1 vccd1 vccd1 _09577_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13245__B1 _12599_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17299__S _17534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11470_ _11470_/A _11470_/B vssd1 vssd1 vccd1 vccd1 _11520_/A sky130_fd_sc_hd__or2_1
XPHY_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16216__B _17517_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17909__S1 _18761_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10421_ _12234_/A vssd1 vssd1 vccd1 vccd1 _10421_/X sky130_fd_sc_hd__buf_4
XANTENNA__16931__S _16950_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13140_ _19162_/Q vssd1 vssd1 vccd1 vccd1 _16210_/A sky130_fd_sc_hd__inv_2
XFILLER_124_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10352_ _10352_/A vssd1 vssd1 vccd1 vccd1 _10353_/B sky130_fd_sc_hd__inv_2
XFILLER_125_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13071_ _13071_/A _13071_/B vssd1 vssd1 vccd1 vccd1 _13193_/A sky130_fd_sc_hd__or2_1
XANTENNA__12760__A _19229_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11079__C _15190_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10283_ _18643_/Q vssd1 vssd1 vccd1 vccd1 _10758_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_151_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12022_ _19348_/Q _12016_/X _09051_/X _12017_/X vssd1 vssd1 vccd1 vccd1 _19348_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__20022__CLK _20091_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16830_ _16721_/Y _19430_/Q _17459_/S vssd1 vssd1 vccd1 vccd1 _16830_/X sky130_fd_sc_hd__mux2_1
XFILLER_238_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18729__RESET_B repeater253/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16761_ vssd1 vssd1 vccd1 vccd1 _16761_/HI _16761_/LO sky130_fd_sc_hd__conb_1
X_13973_ _18701_/Q vssd1 vssd1 vccd1 vccd1 _14031_/A sky130_fd_sc_hd__inv_2
X_18500_ _19795_/CLK _18500_/D repeater219/X vssd1 vssd1 vccd1 vccd1 _18500_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_18_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15712_ _15712_/A _15713_/B vssd1 vssd1 vccd1 vccd1 _18647_/D sky130_fd_sc_hd__nor2_1
X_12924_ _12916_/X _12924_/B _12924_/C _12924_/D vssd1 vssd1 vccd1 vccd1 _12956_/B
+ sky130_fd_sc_hd__and4b_1
XFILLER_234_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17845__S0 _17908_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19480_ _19506_/CLK hold179/X repeater256/X vssd1 vssd1 vccd1 vccd1 _19480_/Q sky130_fd_sc_hd__dfrtp_1
X_16692_ _19465_/Q vssd1 vssd1 vccd1 vccd1 _16692_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18431_ _18431_/CLK _18431_/D vssd1 vssd1 vccd1 vccd1 _18431_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15643_ _15643_/A vssd1 vssd1 vccd1 vccd1 _15643_/X sky130_fd_sc_hd__clkbuf_2
X_12855_ _18923_/Q vssd1 vssd1 vccd1 vccd1 _13002_/A sky130_fd_sc_hd__inv_2
XPHY_4050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11806_ _19456_/Q _11800_/X _09051_/X _11801_/X vssd1 vssd1 vccd1 vccd1 _19456_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_33_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18362_ _19515_/CLK _18362_/D vssd1 vssd1 vccd1 vccd1 _18362_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14984__B1 hold244/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15574_ _10130_/B _15573_/X _15542_/X vssd1 vssd1 vccd1 vccd1 _15574_/X sky130_fd_sc_hd__o21a_1
XPHY_4094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12786_ _19242_/Q vssd1 vssd1 vccd1 vccd1 _12786_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12000__A _12016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11798__B1 _09037_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_230_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14525_ _18325_/Q _14518_/X hold330/X _14520_/X vssd1 vssd1 vccd1 vccd1 _18325_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17313_ _16433_/X _17968_/Q _17564_/S vssd1 vssd1 vccd1 vccd1 _17313_/X sky130_fd_sc_hd__mux2_1
XPHY_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11737_ _11737_/A vssd1 vssd1 vccd1 vccd1 _11737_/X sky130_fd_sc_hd__clkbuf_4
X_18293_ _18435_/CLK _18293_/D vssd1 vssd1 vccd1 vccd1 _18293_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_230_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17002__S _17548_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17244_ _16586_/Y _20108_/Q _17385_/S vssd1 vssd1 vccd1 vccd1 _17244_/X sky130_fd_sc_hd__mux2_1
X_14456_ _18367_/Q _14451_/X _14443_/X _14453_/X vssd1 vssd1 vccd1 vccd1 _18367_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14736__B1 _14604_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11668_ _11668_/A vssd1 vssd1 vccd1 vccd1 _11668_/X sky130_fd_sc_hd__clkbuf_2
XPHY_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13407_ _20108_/Q _13429_/B _20096_/Q _13465_/A vssd1 vssd1 vccd1 vccd1 _13407_/X
+ sky130_fd_sc_hd__o22a_1
X_10619_ _10612_/Y _10598_/A _10617_/X _10567_/C _10618_/X vssd1 vssd1 vccd1 vccd1
+ _10620_/A sky130_fd_sc_hd__o32a_1
XPHY_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17175_ _17174_/X _13074_/A _17542_/S vssd1 vssd1 vccd1 vccd1 _17175_/X sky130_fd_sc_hd__mux2_1
XANTENNA__16841__S _17474_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14387_ _18405_/Q _14380_/X _12726_/X _14382_/X vssd1 vssd1 vccd1 vccd1 _18405_/D
+ sky130_fd_sc_hd__a22o_1
X_11599_ _11583_/A _11583_/B _11569_/A _11597_/Y vssd1 vssd1 vccd1 vccd1 _19570_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_227_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16126_ _19717_/Q vssd1 vssd1 vccd1 vccd1 _16126_/Y sky130_fd_sc_hd__inv_2
X_13338_ _13430_/B _13338_/B vssd1 vssd1 vccd1 vccd1 _13456_/A sky130_fd_sc_hd__or2_1
XFILLER_155_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19170__RESET_B hold370/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16057_ _16051_/Y _15866_/A _10829_/Y _15840_/A _16056_/X vssd1 vssd1 vccd1 vccd1
+ _16057_/X sky130_fd_sc_hd__o221a_1
X_13269_ _14286_/B _13259_/B _14270_/B _17918_/S0 _13268_/Y vssd1 vssd1 vccd1 vccd1
+ _13278_/B sky130_fd_sc_hd__a221o_1
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15008_ _18050_/Q _14993_/A _14842_/X _14994_/A vssd1 vssd1 vccd1 vccd1 _18050_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__20075__RESET_B repeater196/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17672__S _17683_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19816_ _19822_/CLK _19816_/D repeater227/X vssd1 vssd1 vccd1 vccd1 _19816_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__15981__A _19757_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14267__A2 _14259_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19747_ _20070_/CLK _19747_/D repeater205/X vssd1 vssd1 vccd1 vccd1 _19747_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_38_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16959_ _16958_/X _18907_/Q _17542_/S vssd1 vssd1 vccd1 vccd1 _16959_/X sky130_fd_sc_hd__mux2_1
X_09500_ _19312_/Q vssd1 vssd1 vccd1 vccd1 _09500_/Y sky130_fd_sc_hd__inv_2
XFILLER_225_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17836__S0 _17908_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19678_ _19772_/CLK _19678_/D repeater218/X vssd1 vssd1 vccd1 vccd1 _19678_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_53_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09431_ _19387_/Q vssd1 vssd1 vccd1 vccd1 _09431_/Y sky130_fd_sc_hd__inv_2
X_18629_ _19780_/CLK _18629_/D repeater227/X vssd1 vssd1 vccd1 vccd1 _18629_/Q sky130_fd_sc_hd__dfstp_1
X_09362_ _20015_/Q vssd1 vssd1 vccd1 vccd1 _09475_/A sky130_fd_sc_hd__inv_2
XFILLER_212_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11789__B1 _09021_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09293_ _09293_/A vssd1 vssd1 vccd1 vccd1 _09293_/X sky130_fd_sc_hd__buf_1
XANTENNA__19940__RESET_B hold371/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15875__B _15878_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11961__B1 _09051_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_114_HCLK_A clkbuf_opt_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13676__A hold331/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput140 _19672_/Q vssd1 vssd1 vccd1 vccd1 scl_oen_o_S4 sky130_fd_sc_hd__clkbuf_2
XFILLER_217_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17582__S _17584_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15891__A _16633_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18822__RESET_B repeater217/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16652__B1 _17018_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10970_ _10989_/A _17614_/S _10968_/A _10954_/A vssd1 vssd1 vccd1 vccd1 _10970_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__17827__S0 _17918_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14300__A _14300_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09629_ _09629_/A _09629_/B vssd1 vssd1 vccd1 vccd1 _09754_/A sky130_fd_sc_hd__or2_1
XFILLER_15_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12640_ _19006_/Q _12636_/X _12028_/A _12637_/X vssd1 vssd1 vccd1 vccd1 _19006_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_243_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_246_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12571_ _19051_/Q _12569_/X _12389_/X _12570_/X vssd1 vssd1 vccd1 vccd1 _19051_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19681__RESET_B repeater219/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14310_ _18445_/Q _14303_/X _13676_/X _14305_/X vssd1 vssd1 vccd1 vccd1 _18445_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11522_ _19591_/Q _11520_/Y _11521_/X _11522_/C1 vssd1 vssd1 vccd1 vccd1 _19591_/D
+ sky130_fd_sc_hd__o211a_1
X_15290_ _15290_/A vssd1 vssd1 vccd1 vccd1 _15290_/Y sky130_fd_sc_hd__inv_2
XPHY_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14241_ _18666_/Q _14236_/X _18665_/Q _14235_/A vssd1 vssd1 vccd1 vccd1 _18666_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_7_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11453_ _19577_/Q vssd1 vssd1 vccd1 vccd1 _11453_/Y sky130_fd_sc_hd__inv_2
XPHY_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10404_ _10404_/A _14378_/B vssd1 vssd1 vccd1 vccd1 _10404_/Y sky130_fd_sc_hd__nor2_1
X_14172_ _19121_/Q vssd1 vssd1 vccd1 vccd1 _14172_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08948__B2 _08947_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11384_ _19558_/Q vssd1 vssd1 vccd1 vccd1 _11571_/A sky130_fd_sc_hd__inv_2
XFILLER_194_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11952__B1 hold305/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13123_ _19168_/Q vssd1 vssd1 vccd1 vccd1 _13123_/Y sky130_fd_sc_hd__inv_2
XFILLER_194_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10335_ _10335_/A _10335_/B vssd1 vssd1 vccd1 vccd1 _10336_/B sky130_fd_sc_hd__nand2_1
XANTENNA__15143__B1 _09339_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12490__A _12528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18980_ _19597_/CLK _18980_/D repeater281/X vssd1 vssd1 vccd1 vccd1 _18980_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_3_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16891__A0 _16890_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17931_ _19842_/CLK _17931_/D vssd1 vssd1 vccd1 vccd1 _17931_/Q sky130_fd_sc_hd__dfxtp_1
X_13054_ _18892_/Q vssd1 vssd1 vccd1 vccd1 _13065_/A sky130_fd_sc_hd__inv_2
X_10266_ _10266_/A _10266_/B vssd1 vssd1 vccd1 vccd1 _10268_/B sky130_fd_sc_hd__nor2_4
XFILLER_97_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_36_HCLK_A _18641_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17492__S _17546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12005_ _19361_/Q _12000_/X _09021_/X _12003_/X vssd1 vssd1 vccd1 vccd1 _19361_/D
+ sky130_fd_sc_hd__a22o_1
X_17862_ _16260_/Y _16261_/Y _16262_/Y _16263_/Y _17913_/S0 _19632_/Q vssd1 vssd1
+ vccd1 vccd1 _17862_/X sky130_fd_sc_hd__mux4_1
XFILLER_78_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_99_HCLK_A clkbuf_4_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10197_ _19662_/Q vssd1 vssd1 vccd1 vccd1 _10962_/A sky130_fd_sc_hd__inv_2
XFILLER_66_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_238_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19601_ _19608_/CLK _19601_/D hold355/X vssd1 vssd1 vccd1 vccd1 _19601_/Q sky130_fd_sc_hd__dfrtp_4
X_16813_ _15768_/Y _14196_/Y _17546_/S vssd1 vssd1 vccd1 vccd1 _16813_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17793_ _18295_/Q _18287_/Q _18279_/Q _18447_/Q _17923_/S0 _19646_/Q vssd1 vssd1
+ vccd1 vccd1 _17793_/X sky130_fd_sc_hd__mux4_2
XFILLER_213_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19532_ _19544_/CLK _19532_/D repeater221/X vssd1 vssd1 vccd1 vccd1 _19532_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_35_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16744_ hold368/A _17929_/Q vssd1 vssd1 vccd1 vccd1 hold230/A sky130_fd_sc_hd__or2_1
XFILLER_47_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17818__S0 _17918_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13956_ _13949_/A _13949_/B _13954_/Y _13919_/X vssd1 vssd1 vccd1 vccd1 _18712_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_35_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19980__CLK _19992_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19463_ _19470_/CLK _19463_/D repeater273/X vssd1 vssd1 vccd1 vccd1 _19463_/Q sky130_fd_sc_hd__dfrtp_1
X_12907_ _19288_/Q _12887_/C _19272_/Q _13008_/A _12906_/X vssd1 vssd1 vccd1 vccd1
+ _12908_/D sky130_fd_sc_hd__o221a_1
XANTENNA__12680__A1 _18980_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13887_ _19196_/Q vssd1 vssd1 vccd1 vccd1 _13887_/Y sky130_fd_sc_hd__inv_2
X_16675_ _17070_/X _16555_/X _16968_/X _16556_/X vssd1 vssd1 vccd1 vccd1 _16678_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_222_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16836__S _17487_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18414_ _18416_/CLK _18414_/D vssd1 vssd1 vccd1 vccd1 _18414_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_234_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15626_ _18600_/Q _15621_/A _15624_/Y _15621_/Y vssd1 vssd1 vccd1 vccd1 _15627_/B
+ sky130_fd_sc_hd__o22a_1
X_12838_ _18947_/Q vssd1 vssd1 vccd1 vccd1 _12888_/A sky130_fd_sc_hd__inv_2
X_19394_ _19933_/CLK _19394_/D repeater236/X vssd1 vssd1 vccd1 vccd1 _19394_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__12432__A1 _19129_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18345_ _18473_/CLK _18345_/D vssd1 vssd1 vccd1 vccd1 _18345_/Q sky130_fd_sc_hd__dfxtp_1
X_12769_ _12767_/Y _18830_/Q _19238_/Q _13538_/A vssd1 vssd1 vccd1 vccd1 _12769_/X
+ sky130_fd_sc_hd__o22a_1
X_15557_ _15557_/A _15557_/B vssd1 vssd1 vccd1 vccd1 _15557_/Y sky130_fd_sc_hd__nor2_1
XPHY_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10443__B1 _09075_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_230_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_202_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14508_ _18335_/Q _14503_/X _14443_/X _14505_/X vssd1 vssd1 vccd1 vccd1 _18335_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_2_1_0_HCLK_A clkbuf_2_1_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18276_ _19873_/CLK _18276_/D vssd1 vssd1 vccd1 vccd1 _18276_/Q sky130_fd_sc_hd__dfxtp_1
X_15488_ _15491_/B _15487_/Y _15483_/X vssd1 vssd1 vccd1 vccd1 _15488_/X sky130_fd_sc_hd__o21a_1
XANTENNA__19351__RESET_B repeater245/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15906__C1 _15905_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17371__A1 _08937_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15976__A _16055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17227_ _17226_/X _15611_/Y _17318_/S vssd1 vssd1 vccd1 vccd1 _17227_/X sky130_fd_sc_hd__mux2_2
Xinput20 HADDR[27] vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__buf_1
XANTENNA__17667__S _17683_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14439_ _14439_/A vssd1 vssd1 vccd1 vccd1 _14439_/X sky130_fd_sc_hd__clkbuf_2
Xinput31 input31/A vssd1 vssd1 vccd1 vccd1 input31/X sky130_fd_sc_hd__clkbuf_1
XFILLER_174_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12196__B1 _12078_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput42 input42/A vssd1 vssd1 vccd1 vccd1 input42/X sky130_fd_sc_hd__buf_1
Xinput53 input53/A vssd1 vssd1 vccd1 vccd1 input53/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__08939__B2 _18779_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput64 input64/A vssd1 vssd1 vccd1 vccd1 input64/X sky130_fd_sc_hd__buf_2
Xinput75 input75/A vssd1 vssd1 vccd1 vccd1 input75/X sky130_fd_sc_hd__buf_1
X_17158_ _17157_/X _13542_/A _17536_/S vssd1 vssd1 vccd1 vccd1 _17158_/X sky130_fd_sc_hd__mux2_2
XFILLER_128_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11943__B1 _09016_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16109_ _17956_/Q vssd1 vssd1 vccd1 vccd1 _16109_/Y sky130_fd_sc_hd__inv_2
X_17089_ _17088_/X _11450_/Y _17548_/S vssd1 vssd1 vccd1 vccd1 _17089_/X sky130_fd_sc_hd__mux2_1
X_09980_ _09861_/A _09861_/B _09978_/Y _09970_/X vssd1 vssd1 vccd1 vccd1 _19953_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_89_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16882__A0 _17473_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08931_ _10332_/A _18786_/Q _19866_/Q _08930_/Y vssd1 vssd1 vccd1 vccd1 _08931_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_130_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17809__S0 _18751_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12120__B1 _11975_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_1_HCLK clkbuf_1_0_1_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_226_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09414_ _19384_/Q vssd1 vssd1 vccd1 vccd1 _09414_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_241_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19439__RESET_B repeater193/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_110_HCLK clkbuf_opt_0_HCLK/A vssd1 vssd1 vccd1 vccd1 _19109_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_40_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09345_ _20032_/Q vssd1 vssd1 vccd1 vccd1 _09492_/A sky130_fd_sc_hd__inv_2
XFILLER_52_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09276_ _20053_/Q _09269_/X _09098_/X _09271_/X vssd1 vssd1 vccd1 vccd1 _20053_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_166_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17577__S _17584_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09052__B1 _09051_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17114__A1 _08928_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16322__C1 _16321_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16873__A0 _17486_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10120_ _18569_/Q _18568_/Q _15490_/A vssd1 vssd1 vccd1 vccd1 _15498_/A sky130_fd_sc_hd__or3_4
XANTENNA__13687__B1 _13674_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10051_ _10051_/A _10051_/B vssd1 vssd1 vccd1 vccd1 _10052_/C sky130_fd_sc_hd__nor2_1
XFILLER_248_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16625__B1 _17038_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13810_ _18715_/Q vssd1 vssd1 vccd1 vccd1 _13812_/C sky130_fd_sc_hd__inv_2
XFILLER_180_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14790_ _18175_/Q _14785_/X _14751_/X _14787_/X vssd1 vssd1 vccd1 vccd1 _18175_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12111__B1 _12028_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13741_ _13741_/A _13741_/B vssd1 vssd1 vccd1 vccd1 _18751_/D sky130_fd_sc_hd__nor2_1
XFILLER_43_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10953_ _19847_/Q vssd1 vssd1 vccd1 vccd1 _10954_/A sky130_fd_sc_hd__inv_2
XANTENNA__16928__A1 hold202/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_216_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13672_ _13672_/A vssd1 vssd1 vccd1 vccd1 _13672_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_32_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16460_ _17101_/X _16069_/X _17098_/X _16070_/X _16459_/X vssd1 vssd1 vccd1 vccd1
+ _16460_/X sky130_fd_sc_hd__o221a_1
X_10884_ hold245/X vssd1 vssd1 vccd1 vccd1 _14279_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_188_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15411_ _15413_/A _17575_/X vssd1 vssd1 vccd1 vccd1 _18537_/D sky130_fd_sc_hd__and2_1
X_12623_ _12630_/A vssd1 vssd1 vccd1 vccd1 _12623_/X sky130_fd_sc_hd__buf_1
X_16391_ _17326_/X _16069_/X _17323_/X _16070_/X _16390_/X vssd1 vssd1 vccd1 vccd1
+ _16391_/X sky130_fd_sc_hd__o221a_1
XPHY_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15342_ _18493_/Q _14223_/B _14224_/B vssd1 vssd1 vccd1 vccd1 _15342_/X sky130_fd_sc_hd__a21bo_1
X_18130_ _18198_/CLK _18130_/D vssd1 vssd1 vccd1 vccd1 _18130_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12554_ _12551_/A _12553_/A _12249_/A vssd1 vssd1 vccd1 vccd1 _12554_/X sky130_fd_sc_hd__o21a_1
XFILLER_196_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09291__B1 _09086_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11505_ _19601_/Q _11503_/Y _11504_/X _11505_/C1 vssd1 vssd1 vccd1 vccd1 _19601_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__17487__S _17487_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15273_ _18639_/Q _18638_/Q vssd1 vssd1 vccd1 vccd1 _15323_/A sky130_fd_sc_hd__or2_1
X_18061_ _18460_/CLK _18061_/D vssd1 vssd1 vccd1 vccd1 _18061_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12485_ _19094_/Q _12457_/A _12238_/X _12458_/A vssd1 vssd1 vccd1 vccd1 _19094_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_156_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12178__B1 _11924_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14224_ _18494_/Q _14224_/B vssd1 vssd1 vccd1 vccd1 _14225_/B sky130_fd_sc_hd__or2_1
X_17012_ _17473_/A0 _09918_/Y _17522_/S vssd1 vssd1 vccd1 vccd1 _17012_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11436_ _19557_/Q _19137_/Q _11551_/C _11435_/Y vssd1 vssd1 vccd1 vccd1 _11436_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_153_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11925__B1 _11924_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14155_ _19100_/Q vssd1 vssd1 vccd1 vccd1 _14155_/Y sky130_fd_sc_hd__inv_2
X_11367_ _19574_/Q vssd1 vssd1 vccd1 vccd1 _11547_/A sky130_fd_sc_hd__inv_2
XFILLER_152_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14205__A _19110_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16864__A0 _17473_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13106_ _19187_/Q vssd1 vssd1 vccd1 vccd1 _16718_/A sky130_fd_sc_hd__inv_2
XFILLER_140_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10318_ _18766_/Q vssd1 vssd1 vccd1 vccd1 _10319_/A sky130_fd_sc_hd__inv_2
X_14086_ _14084_/Y _18693_/Q _14035_/Y _18681_/Q _14085_/X vssd1 vssd1 vccd1 vccd1
+ _14093_/B sky130_fd_sc_hd__o221a_1
X_18963_ _19137_/CLK _18963_/D repeater249/X vssd1 vssd1 vccd1 vccd1 _18963_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_152_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11298_ _11298_/A _11298_/B _11298_/C _11298_/D vssd1 vssd1 vccd1 vccd1 _11299_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_239_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_160_HCLK_A clkbuf_4_0_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_224_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17914_ _17910_/X _17911_/X _17912_/X _17913_/X _19633_/Q _19634_/Q vssd1 vssd1 vccd1
+ vccd1 _17914_/X sky130_fd_sc_hd__mux4_2
X_13037_ _18909_/Q vssd1 vssd1 vccd1 vccd1 _13081_/A sky130_fd_sc_hd__inv_6
X_10249_ _13642_/B _11863_/A _12053_/B vssd1 vssd1 vccd1 vccd1 _15296_/A sky130_fd_sc_hd__or3_4
XFILLER_67_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18894_ _19214_/CLK _18894_/D hold372/X vssd1 vssd1 vccd1 vccd1 _18894_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_67_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17845_ _16347_/Y _16348_/Y _16349_/Y _16350_/Y _17908_/S0 _18759_/Q vssd1 vssd1
+ vccd1 vccd1 _17845_/X sky130_fd_sc_hd__mux4_2
XFILLER_227_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17776_ _18388_/Q _18380_/Q _18372_/Q _18364_/Q _17923_/S0 _19646_/Q vssd1 vssd1
+ vccd1 vccd1 _17776_/X sky130_fd_sc_hd__mux4_2
XFILLER_240_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14988_ _18059_/Q _14978_/A _14780_/X _14979_/A vssd1 vssd1 vccd1 vccd1 _18059_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_208_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19515_ _19515_/CLK hold226/X repeater259/X vssd1 vssd1 vccd1 vccd1 _19515_/Q sky130_fd_sc_hd__dfrtp_2
Xclkbuf_leaf_133_HCLK clkbuf_4_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19470_/CLK sky130_fd_sc_hd__clkbuf_16
X_16727_ _16800_/X _16597_/X _16829_/X _16598_/X vssd1 vssd1 vccd1 vccd1 _16728_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12653__A1 _18997_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13939_ _18719_/Q _13938_/Y _13819_/B _13925_/X vssd1 vssd1 vccd1 vccd1 _18719_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_223_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19446_ _20058_/CLK _19446_/D repeater194/X vssd1 vssd1 vccd1 vccd1 _19446_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__19532__RESET_B repeater221/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16658_ _19462_/Q vssd1 vssd1 vccd1 vccd1 _16658_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16395__A2 _16148_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19726__CLK _20051_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15609_ _18596_/Q _15605_/A _15608_/Y _15605_/Y vssd1 vssd1 vccd1 vccd1 _15610_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12405__A1 _19146_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19377_ _19971_/CLK _19377_/D repeater191/X vssd1 vssd1 vccd1 vccd1 _19377_/Q sky130_fd_sc_hd__dfrtp_4
X_16589_ _19456_/Q _16622_/B vssd1 vssd1 vccd1 vccd1 _16589_/Y sky130_fd_sc_hd__nand2_1
XFILLER_50_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09130_ _09139_/A _09136_/B _20090_/Q _09129_/Y vssd1 vssd1 vccd1 vccd1 _20090_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_176_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18328_ _19637_/CLK _18328_/D vssd1 vssd1 vccd1 vccd1 _18328_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17344__A1 _17854_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17397__S _17566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09061_ _12028_/A vssd1 vssd1 vccd1 vccd1 _09061_/X sky130_fd_sc_hd__buf_4
X_18259_ _20076_/CLK _18259_/D vssd1 vssd1 vccd1 vccd1 _18259_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__18750__CLK _19900_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19876__CLK _19900_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12169__B1 _11911_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20090__RESET_B repeater204/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09034__B1 _09033_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11916__B1 _10882_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09963_ _09963_/A vssd1 vssd1 vccd1 vccd1 _09963_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13669__B1 _12596_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08914_ _20123_/Q vssd1 vssd1 vccd1 vccd1 _08982_/A sky130_fd_sc_hd__inv_2
XFILLER_134_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20083_ _20085_/CLK _20083_/D repeater204/X vssd1 vssd1 vccd1 vccd1 _20083_/Q sky130_fd_sc_hd__dfrtp_1
X_09894_ _09855_/A _19338_/Q _19944_/Q _09891_/Y _09893_/X vssd1 vssd1 vccd1 vccd1
+ _09895_/D sky130_fd_sc_hd__o221a_1
XFILLER_112_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_82_HCLK_A clkbuf_4_13_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18130__CLK _18198_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17280__A0 _15963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_245_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18280__CLK _19847_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold146_A HADDR[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_241_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09328_ _15721_/A _09317_/X _18656_/Q _18657_/Q vssd1 vssd1 vccd1 vccd1 _09329_/B
+ sky130_fd_sc_hd__a31oi_1
XFILLER_178_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_hold313_A MSI_S3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09273__B1 _09086_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09812__A2 _09807_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20107__RESET_B repeater233/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14149__A1 _18673_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09259_ _10148_/A _09259_/B _10250_/C vssd1 vssd1 vccd1 vccd1 _12256_/C sky130_fd_sc_hd__or3_4
XANTENNA__16505__A _16505_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17100__S _17413_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10256__C _15190_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12270_ _12277_/A vssd1 vssd1 vccd1 vccd1 _12270_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_14_HCLK clkbuf_4_2_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _18198_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_209_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17099__A0 _15963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11907__B1 _09071_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11221_ _11466_/A _18999_/Q _19585_/Q _11220_/Y vssd1 vssd1 vccd1 vccd1 _11221_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_181_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12580__B1 _12406_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11152_ _14335_/A _11151_/X _14335_/A _11151_/X vssd1 vssd1 vccd1 vccd1 _11152_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_161_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10103_ _10103_/A _10103_/B _10107_/C vssd1 vssd1 vccd1 vccd1 _19909_/D sky130_fd_sc_hd__nor3_1
XFILLER_122_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11083_ _19057_/Q vssd1 vssd1 vccd1 vccd1 _12553_/A sky130_fd_sc_hd__inv_2
X_15960_ _20060_/Q _16204_/A vssd1 vssd1 vccd1 vccd1 _15960_/X sky130_fd_sc_hd__and2_1
XANTENNA__16240__A _16637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12332__B1 _12090_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_237_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10034_ _10034_/A _10034_/B vssd1 vssd1 vccd1 vccd1 _10077_/A sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_156_HCLK clkbuf_4_1_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _18416_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_88_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14911_ _18105_/Q _14908_/X _14699_/X _14910_/X vssd1 vssd1 vccd1 vccd1 _18105_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_102_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15891_ _16633_/A vssd1 vssd1 vccd1 vccd1 _16493_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_236_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_236_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17630_ _19889_/Q _19742_/Q _17630_/S vssd1 vssd1 vccd1 vccd1 _17630_/X sky130_fd_sc_hd__mux2_1
X_14842_ _18952_/Q vssd1 vssd1 vccd1 vccd1 _14842_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_236_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19749__CLK _20070_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12635__A1 _19009_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17561_ _17560_/X _08945_/Y _17566_/S vssd1 vssd1 vccd1 vccd1 _17561_/X sky130_fd_sc_hd__mux2_1
X_11985_ _19368_/Q _11977_/X _11922_/X _11979_/X vssd1 vssd1 vccd1 vccd1 _19368_/D
+ sky130_fd_sc_hd__a22o_1
X_14773_ _14773_/A vssd1 vssd1 vccd1 vccd1 _14773_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_90_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19300_ _20013_/CLK _19300_/D repeater242/X vssd1 vssd1 vccd1 vccd1 _19300_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_44_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16512_ _16512_/A vssd1 vssd1 vccd1 vccd1 _16512_/X sky130_fd_sc_hd__buf_2
X_10936_ _10933_/X _10658_/A _10936_/S vssd1 vssd1 vccd1 vccd1 _10937_/A sky130_fd_sc_hd__mux2_1
XFILLER_205_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13724_ _17763_/X vssd1 vssd1 vccd1 vccd1 _13725_/A sky130_fd_sc_hd__inv_2
X_17492_ _15768_/Y _11236_/Y _17546_/S vssd1 vssd1 vccd1 vccd1 _17492_/X sky130_fd_sc_hd__mux2_1
XFILLER_72_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19231_ _19282_/CLK _19231_/D repeater214/X vssd1 vssd1 vccd1 vccd1 _19231_/Q sky130_fd_sc_hd__dfrtp_2
X_16443_ _19716_/Q vssd1 vssd1 vccd1 vccd1 _16443_/Y sky130_fd_sc_hd__inv_2
XFILLER_231_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_repeater170_A _17386_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10867_ _19703_/Q _10856_/A _10866_/X _10857_/A vssd1 vssd1 vccd1 vccd1 _19703_/D
+ sky130_fd_sc_hd__a22o_1
X_13655_ _15199_/A _15169_/A vssd1 vssd1 vccd1 vccd1 _13671_/A sky130_fd_sc_hd__or2_4
XANTENNA__19899__CLK _19900_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12399__B1 _12398_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater268_A repeater269/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12606_ _19027_/Q _12598_/X _12538_/X _12600_/X vssd1 vssd1 vccd1 vccd1 _19027_/D
+ sky130_fd_sc_hd__a22o_1
X_19162_ _19208_/CLK _19162_/D hold370/X vssd1 vssd1 vccd1 vccd1 _19162_/Q sky130_fd_sc_hd__dfrtp_4
X_13586_ _13586_/A vssd1 vssd1 vccd1 vccd1 _13586_/Y sky130_fd_sc_hd__inv_2
X_16374_ _16372_/Y _16303_/X _16373_/Y _15831_/A vssd1 vssd1 vccd1 vccd1 _16374_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10798_ _19736_/Q _10797_/Y _10793_/B vssd1 vssd1 vccd1 vccd1 _19736_/D sky130_fd_sc_hd__o21a_1
XPHY_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18113_ _18137_/CLK _18113_/D vssd1 vssd1 vccd1 vccd1 _18113_/Q sky130_fd_sc_hd__dfxtp_1
X_15325_ _15325_/A vssd1 vssd1 vccd1 vccd1 _18637_/D sky130_fd_sc_hd__inv_2
X_12537_ _19064_/Q _12528_/X _12536_/X _12529_/X vssd1 vssd1 vccd1 vccd1 _19064_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_219_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19093_ _19109_/CLK _19093_/D hold361/X vssd1 vssd1 vccd1 vccd1 _19093_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_173_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18003__CLK _19847_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17010__S _17493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18044_ _19630_/CLK _18044_/D vssd1 vssd1 vccd1 vccd1 _18044_/Q sky130_fd_sc_hd__dfxtp_1
X_15256_ _15256_/A _15286_/B vssd1 vssd1 vccd1 vccd1 _15268_/C sky130_fd_sc_hd__or2_2
XFILLER_8_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12468_ _19107_/Q _12464_/X hold281/X _12465_/X vssd1 vssd1 vccd1 vccd1 _19107_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_8_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11419_ _19136_/Q vssd1 vssd1 vccd1 vccd1 _11419_/Y sky130_fd_sc_hd__inv_2
X_14207_ _14203_/Y _18687_/Q _14204_/Y _18677_/Q _14206_/X vssd1 vssd1 vccd1 vccd1
+ _14218_/A sky130_fd_sc_hd__o221a_1
X_15187_ _17932_/Q _14251_/A _10698_/X _14252_/A vssd1 vssd1 vccd1 vccd1 _17932_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_125_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12399_ _19148_/Q _12388_/X _12398_/X _12390_/X vssd1 vssd1 vccd1 vccd1 _19148_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_235_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12571__B1 _12389_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14138_ _14011_/A _14138_/A2 _14136_/Y _14106_/X vssd1 vssd1 vccd1 vccd1 _18680_/D
+ sky130_fd_sc_hd__a211oi_2
X_19995_ _19997_/CLK _19995_/D repeater192/X vssd1 vssd1 vccd1 vccd1 _19995_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_98_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14069_ _19073_/Q vssd1 vssd1 vccd1 vccd1 _14069_/Y sky130_fd_sc_hd__inv_2
X_18946_ _18947_/CLK _18946_/D repeater211/X vssd1 vssd1 vccd1 vccd1 _18946_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_239_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12323__B1 _12074_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18877_ _20048_/CLK _18877_/D repeater208/X vssd1 vssd1 vccd1 vccd1 _18877_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__19784__RESET_B repeater203/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_227_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17680__S _17683_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17828_ _17933_/Q _18455_/Q _18463_/Q _18063_/Q _17918_/S0 _18750_/Q vssd1 vssd1
+ vccd1 vccd1 _17828_/X sky130_fd_sc_hd__mux4_2
XFILLER_94_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14076__B1 _14072_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17759_ _17762_/S _15194_/Y _17761_/S vssd1 vssd1 vccd1 vccd1 _17759_/X sky130_fd_sc_hd__mux2_1
XFILLER_23_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19429_ _19997_/CLK _19429_/D repeater185/X vssd1 vssd1 vccd1 vccd1 _19429_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_176_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09113_ _09113_/A _09131_/A vssd1 vssd1 vccd1 vccd1 _09133_/C sky130_fd_sc_hd__or2_2
XFILLER_109_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09044_ _20112_/Q _09041_/X hold314/X _09043_/X vssd1 vssd1 vccd1 vccd1 _20112_/D
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_2_0_0_HCLK clkbuf_2_1_0_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_1_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_135_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16044__B _16096_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09946_ _09849_/A _19332_/Q _19955_/Q _09942_/Y _09945_/X vssd1 vssd1 vccd1 vccd1
+ _09947_/D sky130_fd_sc_hd__o221a_1
XFILLER_58_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20066_ _20066_/CLK _20066_/D repeater200/X vssd1 vssd1 vccd1 vccd1 _20066_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_219_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09877_ _09877_/A _09877_/B vssd1 vssd1 vccd1 vccd1 _09878_/A sky130_fd_sc_hd__or2_1
XANTENNA__10820__B _15845_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17253__A0 _17473_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17590__S _17600_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_3_4_0_HCLK_A clkbuf_3_5_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19454__RESET_B repeater272/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater270 repeater272/X vssd1 vssd1 vccd1 vccd1 repeater270/X sky130_fd_sc_hd__buf_8
XFILLER_73_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater281 hold273/X vssd1 vssd1 vccd1 vccd1 repeater281/X sky130_fd_sc_hd__buf_4
XFILLER_39_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12617__A1 _19023_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17005__A0 _17473_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11770_ hold183/X _11764_/X _19476_/Q _11765_/X vssd1 vssd1 vccd1 vccd1 hold185/A
+ sky130_fd_sc_hd__o22a_1
XPHY_4468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10721_ _10721_/A vssd1 vssd1 vccd1 vccd1 _10722_/A sky130_fd_sc_hd__inv_2
XPHY_3767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16934__S _16946_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18026__CLK _19510_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13440_ _18862_/Q _13439_/Y _13426_/X _13350_/B vssd1 vssd1 vccd1 vccd1 _18862_/D
+ sky130_fd_sc_hd__o211a_1
X_10652_ _19792_/Q _10652_/B vssd1 vssd1 vccd1 vccd1 _10653_/B sky130_fd_sc_hd__or2_1
XFILLER_167_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13371_ _20117_/Q _13350_/A _20101_/Q _13470_/A _13370_/X vssd1 vssd1 vccd1 vccd1
+ _13372_/D sky130_fd_sc_hd__o221a_1
XFILLER_10_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10583_ _10583_/A _10583_/B vssd1 vssd1 vccd1 vccd1 _10584_/D sky130_fd_sc_hd__or2_1
XANTENNA__16516__C1 _16515_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16235__A _16688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12322_ _19189_/Q _12318_/X _12069_/X _12321_/X vssd1 vssd1 vccd1 vccd1 _19189_/D
+ sky130_fd_sc_hd__a22o_1
X_15110_ _15111_/A vssd1 vssd1 vccd1 vccd1 _15110_/X sky130_fd_sc_hd__clkbuf_2
X_16090_ _18341_/Q vssd1 vssd1 vccd1 vccd1 _16090_/Y sky130_fd_sc_hd__inv_2
XFILLER_154_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18176__CLK _18198_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16531__A2 _16684_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15041_ _18030_/Q _15035_/X _15000_/X _15037_/X vssd1 vssd1 vccd1 vccd1 _18030_/D
+ sky130_fd_sc_hd__a22o_1
X_12253_ _12253_/A _12253_/B _15232_/C vssd1 vssd1 vccd1 vccd1 _12253_/X sky130_fd_sc_hd__or3_1
XFILLER_181_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16819__A0 _17486_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11204_ _11472_/A _19006_/Q _19596_/Q _11200_/Y _11203_/X vssd1 vssd1 vccd1 vccd1
+ _11223_/A sky130_fd_sc_hd__o221a_1
XFILLER_107_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12184_ _12180_/X _19260_/Q _12184_/S vssd1 vssd1 vccd1 vccd1 _19260_/D sky130_fd_sc_hd__mux2_1
XANTENNA__17492__A0 _15768_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18800_ _19900_/CLK _18800_/D repeater199/X vssd1 vssd1 vccd1 vccd1 _18800_/Q sky130_fd_sc_hd__dfrtp_4
X_11135_ _19630_/Q _11133_/Y _12708_/C vssd1 vssd1 vccd1 vccd1 _11135_/X sky130_fd_sc_hd__a21o_1
X_19780_ _19780_/CLK _19780_/D repeater227/X vssd1 vssd1 vccd1 vccd1 _19780_/Q sky130_fd_sc_hd__dfrtp_4
X_16992_ _16991_/X _19961_/Q _17488_/S vssd1 vssd1 vccd1 vccd1 _16992_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12305__B1 _12234_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18731_ _19224_/CLK _18731_/D repeater186/X vssd1 vssd1 vccd1 vccd1 _18731_/Q sky130_fd_sc_hd__dfrtp_1
X_11066_ _19633_/Q _11066_/B vssd1 vssd1 vccd1 vccd1 _11123_/B sky130_fd_sc_hd__nand2_1
XFILLER_95_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15943_ _17970_/Q vssd1 vssd1 vccd1 vccd1 _15943_/Y sky130_fd_sc_hd__inv_2
X_10017_ _10043_/A _10042_/A _10035_/A _10034_/A vssd1 vssd1 vccd1 vccd1 _10019_/C
+ sky130_fd_sc_hd__or4_4
XFILLER_209_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10867__B1 _10866_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18662_ _20055_/CLK hold312/X repeater204/X vssd1 vssd1 vccd1 vccd1 _18662_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12003__A _12017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19195__RESET_B repeater188/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15874_ _19938_/Q vssd1 vssd1 vccd1 vccd1 _15874_/Y sky130_fd_sc_hd__inv_2
XFILLER_237_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17613_ _15223_/Y _12247_/A _17614_/S vssd1 vssd1 vccd1 vccd1 _17613_/X sky130_fd_sc_hd__mux2_1
X_14825_ _18159_/Q _14820_/X _14751_/X _14822_/X vssd1 vssd1 vccd1 vccd1 _18159_/D
+ sky130_fd_sc_hd__a22o_1
X_18593_ _19667_/CLK _18593_/D repeater264/X vssd1 vssd1 vccd1 vccd1 _18593_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_221_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17890__S1 _19632_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17005__S _17512_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17544_ _17543_/X _14072_/Y _17544_/S vssd1 vssd1 vccd1 vccd1 _17544_/X sky130_fd_sc_hd__mux2_1
X_14756_ _18195_/Q _14746_/A _14691_/X _14747_/A vssd1 vssd1 vccd1 vccd1 _18195_/D
+ sky130_fd_sc_hd__a22o_1
X_11968_ _19378_/Q _11962_/X _09067_/X _11963_/X vssd1 vssd1 vccd1 vccd1 _19378_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_32_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13707_ _13707_/A vssd1 vssd1 vccd1 vccd1 _13707_/Y sky130_fd_sc_hd__inv_2
XFILLER_220_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10919_ _19682_/Q _10918_/X _18510_/Q _10914_/Y vssd1 vssd1 vccd1 vccd1 _19682_/D
+ sky130_fd_sc_hd__a211o_1
X_17475_ _17486_/A0 _15965_/Y _17517_/S vssd1 vssd1 vccd1 vccd1 _17475_/X sky130_fd_sc_hd__mux2_1
XANTENNA__16844__S _17548_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14687_ _18231_/Q _14682_/X _14606_/X _14684_/X vssd1 vssd1 vccd1 vccd1 _18231_/D
+ sky130_fd_sc_hd__a22o_1
X_11899_ _11915_/A vssd1 vssd1 vccd1 vccd1 _11899_/X sky130_fd_sc_hd__clkbuf_2
X_19214_ _19214_/CLK _19214_/D hold367/X vssd1 vssd1 vccd1 vccd1 _19214_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_149_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16426_ _18081_/Q vssd1 vssd1 vccd1 vccd1 _16426_/Y sky130_fd_sc_hd__inv_2
X_13638_ _13635_/A _13637_/A _12058_/B vssd1 vssd1 vccd1 vccd1 _13638_/X sky130_fd_sc_hd__o21a_1
XFILLER_60_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19145_ _19566_/CLK _19145_/D repeater255/X vssd1 vssd1 vccd1 vccd1 _19145_/Q sky130_fd_sc_hd__dfrtp_1
X_16357_ _18264_/Q vssd1 vssd1 vccd1 vccd1 _16357_/Y sky130_fd_sc_hd__inv_2
XFILLER_201_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13569_ _13569_/A vssd1 vssd1 vccd1 vccd1 _13569_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15308_ _15302_/Y _15307_/X _15290_/A vssd1 vssd1 vccd1 vccd1 _18627_/D sky130_fd_sc_hd__o21ai_1
XFILLER_157_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19076_ _19610_/CLK _19076_/D hold343/X vssd1 vssd1 vccd1 vccd1 _19076_/Q sky130_fd_sc_hd__dfrtp_1
X_16288_ _18087_/Q vssd1 vssd1 vccd1 vccd1 _16288_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16522__A2 _15896_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18027_ _18142_/CLK _18027_/D vssd1 vssd1 vccd1 vccd1 _18027_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17675__S _17683_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15239_ _18519_/Q vssd1 vssd1 vccd1 vccd1 _15304_/A sky130_fd_sc_hd__inv_2
XFILLER_160_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12544__B1 _12543_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17483__A0 _15963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09800_ _09800_/A vssd1 vssd1 vccd1 vccd1 _09800_/Y sky130_fd_sc_hd__inv_2
X_19978_ _19992_/CLK _19978_/D repeater192/X vssd1 vssd1 vccd1 vccd1 _19978_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__14297__B1 _13680_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18929_ _19325_/CLK _18929_/D repeater213/X vssd1 vssd1 vccd1 vccd1 _18929_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_68_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09731_ _09731_/A vssd1 vssd1 vccd1 vccd1 _09731_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_140_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0_HCLK HCLK vssd1 vssd1 vccd1 vccd1 clkbuf_0_HCLK/X sky130_fd_sc_hd__clkbuf_16
XFILLER_67_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10858__B1 _10446_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09662_ _19994_/Q vssd1 vssd1 vccd1 vccd1 _09750_/A sky130_fd_sc_hd__inv_2
XFILLER_28_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_227_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09593_ _20021_/Q _09592_/Y _09482_/B _09581_/X vssd1 vssd1 vccd1 vccd1 _20021_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__17881__S1 _19632_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18847__RESET_B repeater232/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15878__B _15878_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12583__A _12598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16055__A _16055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09027_ hold286/X vssd1 vssd1 vccd1 vccd1 _09027_/X sky130_fd_sc_hd__buf_4
XFILLER_163_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold250 hold250/A vssd1 vssd1 vccd1 vccd1 hold250/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold261 HWDATA[8] vssd1 vssd1 vccd1 vccd1 input68/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold272 HWDATA[12] vssd1 vssd1 vccd1 vccd1 input41/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold283 HWDATA[14] vssd1 vssd1 vccd1 vccd1 input43/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 input46/X vssd1 vssd1 vccd1 vccd1 hold294/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19635__RESET_B repeater258/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20118_ _20120_/CLK _20118_/D repeater217/X vssd1 vssd1 vccd1 vccd1 _20118_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_131_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09929_ _19335_/Q vssd1 vssd1 vccd1 vccd1 _16215_/A sky130_fd_sc_hd__inv_2
XANTENNA__17226__A0 _17473_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16929__S _16950_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10849__B1 _10418_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20049_ _20049_/CLK _20049_/D repeater208/X vssd1 vssd1 vccd1 vccd1 _20049_/Q sky130_fd_sc_hd__dfrtp_1
X_12940_ _12936_/Y _18920_/Q _12937_/Y _18922_/Q _12939_/X vssd1 vssd1 vccd1 vccd1
+ _12941_/D sky130_fd_sc_hd__o221a_1
XFILLER_219_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_234_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12871_ _13002_/A _13001_/C _12871_/C _12871_/D vssd1 vssd1 vccd1 vccd1 _12967_/A
+ sky130_fd_sc_hd__or4_4
XPHY_4221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17872__S1 _19632_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14610_ _18276_/Q _14601_/A _14582_/X _14602_/A vssd1 vssd1 vccd1 vccd1 _18276_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_65_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11822_ _11822_/A vssd1 vssd1 vccd1 vccd1 _11822_/X sky130_fd_sc_hd__clkbuf_2
XPHY_4254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15590_ _15643_/A vssd1 vssd1 vccd1 vccd1 _15590_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_61_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14460__B1 _14403_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14541_ _18316_/Q _14532_/A _14513_/X _14533_/A vssd1 vssd1 vccd1 vccd1 _18316_/D
+ sky130_fd_sc_hd__a22o_1
X_11753_ hold133/X _11750_/X _19489_/Q _11751_/X vssd1 vssd1 vccd1 vccd1 hold135/A
+ sky130_fd_sc_hd__o22a_1
XPHY_4298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18588__RESET_B repeater269/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10704_ _15391_/A _10704_/B vssd1 vssd1 vccd1 vccd1 _10716_/S sky130_fd_sc_hd__or2_2
XPHY_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17260_ _17259_/X _19143_/Q _17548_/S vssd1 vssd1 vccd1 vccd1 _17260_/X sky130_fd_sc_hd__mux2_1
XPHY_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11684_ _10508_/A _11674_/X _10516_/A _11675_/X vssd1 vssd1 vccd1 vccd1 _19533_/D
+ sky130_fd_sc_hd__o22ai_1
XPHY_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14472_ hold335/X vssd1 vssd1 vccd1 vccd1 hold334/A sky130_fd_sc_hd__buf_2
XFILLER_42_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08971__A _13285_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16211_ _16211_/A _16212_/B vssd1 vssd1 vccd1 vccd1 _16211_/Y sky130_fd_sc_hd__nor2_1
XPHY_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10635_ _19800_/Q _10609_/A _10594_/C _10606_/X vssd1 vssd1 vccd1 vccd1 _19800_/D
+ sky130_fd_sc_hd__o22a_1
X_13423_ _13423_/A vssd1 vssd1 vccd1 vccd1 _13445_/A sky130_fd_sc_hd__clkbuf_2
XPHY_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17191_ _15768_/Y _11230_/Y _17546_/S vssd1 vssd1 vccd1 vccd1 _17191_/X sky130_fd_sc_hd__mux2_1
XFILLER_195_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13354_ _13354_/A _13354_/B vssd1 vssd1 vccd1 vccd1 _13355_/A sky130_fd_sc_hd__or2_1
X_16142_ _17427_/X vssd1 vssd1 vccd1 vccd1 _16142_/Y sky130_fd_sc_hd__inv_2
X_10566_ _19810_/Q vssd1 vssd1 vccd1 vccd1 _10567_/C sky130_fd_sc_hd__inv_2
XANTENNA__18811__CLK _20115_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12305_ _19196_/Q _12298_/X _12234_/X _12300_/X vssd1 vssd1 vccd1 vccd1 _19196_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17495__S _19498_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16073_ _17460_/X _15904_/A _17467_/X _15999_/X vssd1 vssd1 vccd1 vccd1 _16073_/X
+ sky130_fd_sc_hd__o22a_1
X_13285_ _13285_/A _13285_/B vssd1 vssd1 vccd1 vccd1 _15192_/B sky130_fd_sc_hd__nand2_1
X_10497_ _10734_/A vssd1 vssd1 vccd1 vccd1 _10519_/D sky130_fd_sc_hd__inv_2
XFILLER_114_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11329__B2 _18980_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12526__B1 hold259/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_9_0_HCLK clkbuf_4_9_0_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_9_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_15024_ _15024_/A vssd1 vssd1 vccd1 vccd1 _15025_/A sky130_fd_sc_hd__inv_2
X_19901_ _20123_/CLK _19901_/D repeater195/X vssd1 vssd1 vccd1 vccd1 _19901_/Q sky130_fd_sc_hd__dfrtp_1
X_12236_ _13678_/A vssd1 vssd1 vccd1 vccd1 _12236_/X sky130_fd_sc_hd__buf_4
XFILLER_170_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19832_ _20058_/CLK _19832_/D repeater194/X vssd1 vssd1 vccd1 vccd1 _19832_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__11837__A _15867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12167_ _19272_/Q _12164_/X _12038_/X _12165_/X vssd1 vssd1 vccd1 vccd1 _19272_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19376__RESET_B repeater241/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11118_ _11118_/A vssd1 vssd1 vccd1 vccd1 _19637_/D sky130_fd_sc_hd__inv_2
X_19763_ _19772_/CLK _19763_/D repeater218/X vssd1 vssd1 vccd1 vccd1 _19763_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16975_ _16617_/Y _19081_/Q _17544_/S vssd1 vssd1 vccd1 vccd1 _16975_/X sky130_fd_sc_hd__mux2_1
X_12098_ hold301/X vssd1 vssd1 vccd1 vccd1 _12098_/X sky130_fd_sc_hd__buf_2
XANTENNA__16839__S _17318_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18714_ _18718_/CLK _18714_/D repeater252/X vssd1 vssd1 vccd1 vccd1 _18714_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_232_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11049_ _11049_/A vssd1 vssd1 vccd1 vccd1 _11049_/Y sky130_fd_sc_hd__inv_2
X_15926_ _18051_/Q vssd1 vssd1 vccd1 vccd1 _15926_/Y sky130_fd_sc_hd__inv_2
X_19694_ _20051_/CLK _19694_/D repeater208/X vssd1 vssd1 vccd1 vccd1 _19694_/Q sky130_fd_sc_hd__dfrtp_1
Xinput7 input7/A vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_1
XFILLER_37_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18645_ _20059_/CLK _18645_/D repeater197/X vssd1 vssd1 vccd1 vccd1 _18645_/Q sky130_fd_sc_hd__dfrtp_1
X_15857_ _15852_/Y _15836_/X _15853_/Y _15838_/X _15856_/X vssd1 vssd1 vccd1 vccd1
+ _15857_/X sky130_fd_sc_hd__o221a_2
XFILLER_37_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17863__S1 _19632_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_224_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14808_ _14808_/A vssd1 vssd1 vccd1 vccd1 _14808_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_18_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18576_ _19437_/CLK _18576_/D repeater269/X vssd1 vssd1 vccd1 vccd1 _18576_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_224_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15788_ _18034_/Q vssd1 vssd1 vccd1 vccd1 _15788_/Y sky130_fd_sc_hd__inv_2
XFILLER_205_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09042__A hold315/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17527_ _17526_/X _15872_/Y _17539_/S vssd1 vssd1 vccd1 vccd1 _17527_/X sky130_fd_sc_hd__mux2_1
X_14739_ _18205_/Q _14732_/X _14725_/X _14734_/X vssd1 vssd1 vccd1 vccd1 _18205_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_189_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17458_ _15768_/Y _11292_/Y _17546_/S vssd1 vssd1 vccd1 vccd1 _17458_/X sky130_fd_sc_hd__mux2_1
X_16409_ _18353_/Q vssd1 vssd1 vccd1 vccd1 _16409_/Y sky130_fd_sc_hd__inv_2
X_17389_ _16209_/Y _19065_/Q _17544_/S vssd1 vssd1 vccd1 vccd1 _17389_/X sky130_fd_sc_hd__mux2_1
XFILLER_119_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19128_ _19970_/CLK _19128_/D repeater249/X vssd1 vssd1 vccd1 vccd1 _19128_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_173_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19059_ _19630_/CLK _19059_/D repeater257/X vssd1 vssd1 vccd1 vccd1 _19059_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_133_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12517__B1 hold256/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11740__B2 _11738_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09714_ _19406_/Q vssd1 vssd1 vccd1 vccd1 _09714_/Y sky130_fd_sc_hd__inv_2
XFILLER_142_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14690__B1 _14582_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09645_ _19982_/Q vssd1 vssd1 vccd1 vccd1 _09794_/A sky130_fd_sc_hd__inv_2
XFILLER_16_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17854__S1 _19634_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09576_ _09490_/A _09490_/B _09607_/A _09574_/Y vssd1 vssd1 vccd1 vccd1 _20030_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_71_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14442__B1 _14441_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_137_HCLK_A clkbuf_4_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_212_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15889__A _16637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14793__A _14793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18681__RESET_B hold359/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10420_ _19846_/Q _10417_/X _10418_/X _10419_/Y vssd1 vssd1 vccd1 vccd1 _19846_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_149_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16498__A1 _17208_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10351_ _10351_/A vssd1 vssd1 vccd1 vccd1 _19863_/D sky130_fd_sc_hd__inv_2
XANTENNA__16498__B2 _15889_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16513__A _16513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12508__B1 _12404_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17790__S0 _17923_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11151__A1_N _19648_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13070_ _13070_/A _13070_/B vssd1 vssd1 vccd1 vccd1 _13071_/B sky130_fd_sc_hd__or2_2
XFILLER_151_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10282_ _17746_/X _17753_/S _12058_/A _10281_/X vssd1 vssd1 vccd1 vccd1 _19873_/D
+ sky130_fd_sc_hd__a22oi_1
XFILLER_140_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12021_ _19349_/Q _12016_/X _09049_/X _12017_/X vssd1 vssd1 vccd1 vccd1 _19349_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_105_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16760_ vssd1 vssd1 vccd1 vccd1 _16760_/HI _16760_/LO sky130_fd_sc_hd__conb_1
XFILLER_76_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13972_ _18702_/Q vssd1 vssd1 vccd1 vccd1 _14032_/A sky130_fd_sc_hd__inv_2
XANTENNA__08966__A _18778_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15711_ _15711_/A _15713_/B vssd1 vssd1 vccd1 vccd1 _18646_/D sky130_fd_sc_hd__nor2_1
XFILLER_246_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12923_ _12922_/Y _12859_/B _19264_/Q _18921_/Q vssd1 vssd1 vccd1 vccd1 _12924_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16691_ _16682_/X _16691_/B _16691_/C vssd1 vssd1 vccd1 vccd1 _16691_/Y sky130_fd_sc_hd__nand3b_4
XANTENNA__17845__S1 _18759_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12488__A _12528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18430_ _18795_/CLK _18430_/D vssd1 vssd1 vccd1 vccd1 _18430_/Q sky130_fd_sc_hd__dfxtp_1
X_15642_ _15642_/A _15642_/B vssd1 vssd1 vccd1 vccd1 _15642_/Y sky130_fd_sc_hd__nor2_1
XFILLER_234_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12854_ _19191_/Q vssd1 vssd1 vccd1 vccd1 _13000_/A sky130_fd_sc_hd__inv_2
XPHY_4051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14433__B1 _14403_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18361_ _19849_/CLK _18361_/D vssd1 vssd1 vccd1 vccd1 _18361_/Q sky130_fd_sc_hd__dfxtp_1
X_11805_ _19457_/Q _11800_/X _09049_/X _11801_/X vssd1 vssd1 vccd1 vccd1 _19457_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output100_A _16728_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15573_ _18586_/Q _15566_/A _18587_/Q vssd1 vssd1 vccd1 vccd1 _15573_/X sky130_fd_sc_hd__o21a_1
XPHY_4095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12785_ _18821_/Q vssd1 vssd1 vccd1 vccd1 _13544_/A sky130_fd_sc_hd__inv_2
XPHY_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17312_ _16434_/X _18779_/Q _17566_/S vssd1 vssd1 vccd1 vccd1 _17312_/X sky130_fd_sc_hd__mux2_1
X_14524_ _18326_/Q _14518_/X _14509_/X _14520_/X vssd1 vssd1 vccd1 vccd1 _18326_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18292_ _18435_/CLK _18292_/D vssd1 vssd1 vccd1 vccd1 _18292_/Q sky130_fd_sc_hd__dfxtp_1
X_11736_ _19501_/Q _11730_/X _16933_/X _11731_/X vssd1 vssd1 vccd1 vccd1 hold231/A
+ sky130_fd_sc_hd__a22o_1
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_230_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_59_HCLK_A clkbuf_4_12_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17243_ _17242_/X _13888_/Y _17545_/S vssd1 vssd1 vccd1 vccd1 _17243_/X sky130_fd_sc_hd__mux2_1
XPHY_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14455_ _18368_/Q _14451_/X _14441_/X _14453_/X vssd1 vssd1 vccd1 vccd1 _18368_/D
+ sky130_fd_sc_hd__a22o_1
X_11667_ _19544_/Q _11669_/A _11651_/B _11666_/X vssd1 vssd1 vccd1 vccd1 _19544_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_202_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13406_ _20096_/Q vssd1 vssd1 vccd1 vccd1 _13406_/Y sky130_fd_sc_hd__clkinvlp_4
XPHY_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10618_ _10618_/A vssd1 vssd1 vccd1 vccd1 _10618_/X sky130_fd_sc_hd__clkbuf_2
XPHY_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17174_ _17173_/X _12948_/Y _17541_/S vssd1 vssd1 vccd1 vccd1 _17174_/X sky130_fd_sc_hd__mux2_1
X_11598_ _11584_/A _11597_/A _19571_/Q _11597_/Y _11588_/X vssd1 vssd1 vccd1 vccd1
+ _19571_/D sky130_fd_sc_hd__o221a_1
X_14386_ _18406_/Q _14380_/X _12723_/X _14382_/X vssd1 vssd1 vccd1 vccd1 _18406_/D
+ sky130_fd_sc_hd__a22o_1
X_16125_ _19688_/Q vssd1 vssd1 vccd1 vccd1 _16125_/Y sky130_fd_sc_hd__inv_2
XFILLER_227_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10549_ _19810_/Q _10567_/D vssd1 vssd1 vccd1 vccd1 _10582_/A sky130_fd_sc_hd__or2_1
X_13337_ _13428_/C _13459_/A vssd1 vssd1 vccd1 vccd1 _13338_/B sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_4_7_0_HCLK_A clkbuf_4_7_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19557__RESET_B hold348/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17781__S0 _17923_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16056_ _16052_/Y _16053_/X _16054_/Y _16055_/X vssd1 vssd1 vccd1 vccd1 _16056_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_142_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15161__B2 _15160_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13268_ _17745_/X vssd1 vssd1 vccd1 vccd1 _13268_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15007_ _18051_/Q _14993_/A _15006_/X _14994_/A vssd1 vssd1 vccd1 vccd1 _18051_/D
+ sky130_fd_sc_hd__a22o_1
X_12219_ _12228_/A vssd1 vssd1 vccd1 vccd1 _12219_/X sky130_fd_sc_hd__clkbuf_2
X_13199_ _13199_/A _13199_/B _13199_/C vssd1 vssd1 vccd1 vccd1 _18897_/D sky130_fd_sc_hd__nor3_1
XFILLER_243_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09037__A hold296/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19815_ _19825_/CLK _19815_/D repeater228/X vssd1 vssd1 vccd1 vccd1 _19815_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_229_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19746_ _20070_/CLK _19746_/D repeater205/X vssd1 vssd1 vccd1 vccd1 _19746_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_37_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16958_ _16618_/Y _19282_/Q _17541_/S vssd1 vssd1 vccd1 vccd1 _16958_/X sky130_fd_sc_hd__mux2_1
X_15909_ _15909_/A vssd1 vssd1 vccd1 vccd1 _15999_/A sky130_fd_sc_hd__clkbuf_2
X_19677_ _19772_/CLK _19677_/D repeater201/X vssd1 vssd1 vccd1 vccd1 _19677_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12398__A hold298/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16889_ _15768_/Y _14211_/Y _17546_/S vssd1 vssd1 vccd1 vccd1 _16889_/X sky130_fd_sc_hd__mux2_1
XANTENNA__17836__S1 _18759_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09430_ _19366_/Q vssd1 vssd1 vccd1 vccd1 _09430_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18628_ _19545_/CLK _18628_/D repeater221/X vssd1 vssd1 vccd1 vccd1 _18628_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_80_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18857__CLK _18866_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09361_ _20016_/Q vssd1 vssd1 vccd1 vccd1 _09476_/A sky130_fd_sc_hd__inv_2
XFILLER_52_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18559_ _19992_/CLK _18559_/D repeater193/X vssd1 vssd1 vccd1 vccd1 _18559_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_205_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09292_ _20045_/Q _09285_/X _09090_/X _09287_/X vssd1 vssd1 vccd1 vccd1 _20045_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_20_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19980__RESET_B repeater192/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11961__A1 _19383_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17772__S0 _17923_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15152__B2 _15148_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput130 _18641_/Q vssd1 vssd1 vccd1 vccd1 RsTx_S0 sky130_fd_sc_hd__clkbuf_2
XFILLER_161_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput141 _19814_/Q vssd1 vssd1 vccd1 vccd1 scl_oen_o_S5 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11713__A1 _12370_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11713__B2 _16950_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17827__S1 _18750_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18862__RESET_B repeater232/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09628_ _19999_/Q vssd1 vssd1 vccd1 vccd1 _09629_/B sky130_fd_sc_hd__inv_2
XFILLER_244_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09559_ _19310_/Q vssd1 vssd1 vccd1 vccd1 _09559_/Y sky130_fd_sc_hd__inv_2
XPHY_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16508__A _16638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11940__A _11977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17103__S _17548_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12570_ _12577_/A vssd1 vssd1 vccd1 vccd1 _12570_/X sky130_fd_sc_hd__buf_1
XFILLER_24_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16168__B1 _11023_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11521_ _11521_/A vssd1 vssd1 vccd1 vccd1 _11521_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_156_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16942__S _16946_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14240_ _18667_/Q _14236_/X _18666_/Q _14235_/A vssd1 vssd1 vccd1 vccd1 _18667_/D
+ sky130_fd_sc_hd__a22o_1
X_11452_ _19141_/Q vssd1 vssd1 vccd1 vccd1 _11452_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10403_ _10403_/A vssd1 vssd1 vccd1 vccd1 _14378_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__08948__A2 _08946_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14171_ _19094_/Q vssd1 vssd1 vccd1 vccd1 _14171_/Y sky130_fd_sc_hd__inv_2
XFILLER_137_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11383_ _11623_/A _19133_/Q _19553_/Q _11379_/Y _11382_/X vssd1 vssd1 vccd1 vccd1
+ _11389_/C sky130_fd_sc_hd__o221a_1
XFILLER_152_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11952__A1 _19390_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10334_ _10368_/A vssd1 vssd1 vccd1 vccd1 _10335_/B sky130_fd_sc_hd__inv_2
X_13122_ _19176_/Q vssd1 vssd1 vccd1 vccd1 _13122_/Y sky130_fd_sc_hd__inv_2
XFILLER_180_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17930_ _18869_/CLK _17930_/D vssd1 vssd1 vccd1 vccd1 _17930_/Q sky130_fd_sc_hd__dfxtp_1
X_13053_ _18893_/Q vssd1 vssd1 vccd1 vccd1 _13066_/A sky130_fd_sc_hd__inv_2
XFILLER_180_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10265_ _19645_/Q vssd1 vssd1 vccd1 vccd1 _10266_/B sky130_fd_sc_hd__inv_2
XFILLER_127_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12004_ _19362_/Q _12000_/X _09016_/X _12003_/X vssd1 vssd1 vccd1 vccd1 _19362_/D
+ sky130_fd_sc_hd__a22o_1
X_17861_ _16256_/Y _16257_/Y _16258_/Y _16259_/Y _17913_/S0 _19632_/Q vssd1 vssd1
+ vccd1 vccd1 _17861_/X sky130_fd_sc_hd__mux4_2
X_10196_ _10196_/A _10196_/B vssd1 vssd1 vccd1 vccd1 _11863_/A sky130_fd_sc_hd__or2_2
XANTENNA__14103__C1 _14135_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19600_ _19600_/CLK _19600_/D hold355/X vssd1 vssd1 vccd1 vccd1 _19600_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_66_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16812_ _16811_/X _13860_/Y _17545_/S vssd1 vssd1 vccd1 vccd1 _16812_/X sky130_fd_sc_hd__mux2_1
X_17792_ _18327_/Q _18007_/Q _18311_/Q _18303_/Q _17923_/S0 _19646_/Q vssd1 vssd1
+ vccd1 vccd1 _17792_/X sky130_fd_sc_hd__mux4_2
XFILLER_143_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19531_ _19544_/CLK _19531_/D repeater221/X vssd1 vssd1 vccd1 vccd1 _19531_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_207_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16743_ _16682_/A _16743_/B _16743_/C vssd1 vssd1 vccd1 vccd1 _16743_/Y sky130_fd_sc_hd__nand3b_4
X_13955_ _18713_/Q _13954_/Y _13951_/B _13925_/X vssd1 vssd1 vccd1 vccd1 _18713_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__17818__S1 _18750_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12906_ _19278_/Q _12877_/A _12905_/Y _18935_/Q vssd1 vssd1 vccd1 vccd1 _12906_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_35_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19462_ _19462_/CLK _19462_/D repeater273/X vssd1 vssd1 vccd1 vccd1 _19462_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_74_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16674_ _16965_/X _16563_/X _16996_/X _16591_/X vssd1 vssd1 vccd1 vccd1 _16678_/A
+ sky130_fd_sc_hd__o22ai_4
XANTENNA__14406__B1 _14405_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13886_ _19218_/Q vssd1 vssd1 vccd1 vccd1 _13886_/Y sky130_fd_sc_hd__inv_2
X_18413_ _18416_/CLK _18413_/D vssd1 vssd1 vccd1 vccd1 _18413_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_222_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15625_ _15702_/A vssd1 vssd1 vccd1 vccd1 _15666_/A sky130_fd_sc_hd__clkbuf_2
X_19393_ _19933_/CLK _19393_/D repeater236/X vssd1 vssd1 vccd1 vccd1 _19393_/Q sky130_fd_sc_hd__dfrtp_1
X_12837_ _18949_/Q vssd1 vssd1 vccd1 vccd1 _12891_/A sky130_fd_sc_hd__inv_2
XANTENNA__17013__S _17523_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_120_HCLK_A clkbuf_4_4_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18344_ _18473_/CLK _18344_/D vssd1 vssd1 vccd1 vccd1 _18344_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15556_ _15556_/A vssd1 vssd1 vccd1 vccd1 _15556_/Y sky130_fd_sc_hd__inv_2
X_12768_ _18815_/Q vssd1 vssd1 vccd1 vccd1 _13538_/A sky130_fd_sc_hd__inv_2
XPHY_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14507_ _18336_/Q _14503_/X _14441_/X _14505_/X vssd1 vssd1 vccd1 vccd1 _18336_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10443__A1 _19836_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18275_ _19873_/CLK _18275_/D vssd1 vssd1 vccd1 vccd1 _18275_/Q sky130_fd_sc_hd__dfxtp_1
X_11719_ _19514_/Q _11716_/X _16946_/X _11717_/X vssd1 vssd1 vccd1 vccd1 hold216/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16852__S _17535_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15487_ _15487_/A _15487_/B vssd1 vssd1 vccd1 vccd1 _15487_/Y sky130_fd_sc_hd__nor2_1
XFILLER_202_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12699_ _12699_/A vssd1 vssd1 vccd1 vccd1 _12699_/X sky130_fd_sc_hd__buf_1
XPHY_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_238_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17226_ _17473_/A0 _16486_/Y _17473_/S vssd1 vssd1 vccd1 vccd1 _17226_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14438_ _14438_/A vssd1 vssd1 vccd1 vccd1 _14439_/A sky130_fd_sc_hd__inv_2
Xinput10 input10/A vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__clkbuf_1
Xinput21 HADDR[28] vssd1 vssd1 vccd1 vccd1 input21/X sky130_fd_sc_hd__buf_1
Xclkbuf_leaf_70_HCLK clkbuf_opt_2_HCLK/X vssd1 vssd1 vccd1 vccd1 _19541_/CLK sky130_fd_sc_hd__clkbuf_16
Xinput32 input32/A vssd1 vssd1 vccd1 vccd1 input32/X sky130_fd_sc_hd__clkbuf_1
Xinput43 input43/A vssd1 vssd1 vccd1 vccd1 input43/X sky130_fd_sc_hd__buf_1
XANTENNA__13393__B1 _13391_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput54 input54/A vssd1 vssd1 vccd1 vccd1 input54/X sky130_fd_sc_hd__clkbuf_4
X_17157_ _17156_/X _13409_/Y _17535_/S vssd1 vssd1 vccd1 vccd1 _17157_/X sky130_fd_sc_hd__mux2_1
Xinput65 input65/A vssd1 vssd1 vccd1 vccd1 input65/X sky130_fd_sc_hd__buf_4
X_14369_ _14369_/A vssd1 vssd1 vccd1 vccd1 _14369_/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput76 input76/A vssd1 vssd1 vccd1 vccd1 input76/X sky130_fd_sc_hd__buf_1
X_16108_ _17980_/Q vssd1 vssd1 vccd1 vccd1 _16108_/Y sky130_fd_sc_hd__inv_2
XFILLER_171_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17088_ _17087_/X _11300_/Y _17493_/S vssd1 vssd1 vccd1 vccd1 _17088_/X sky130_fd_sc_hd__mux2_1
XFILLER_104_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19655__CLK _19847_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17683__S _17683_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08930_ _18786_/Q vssd1 vssd1 vccd1 vccd1 _08930_/Y sky130_fd_sc_hd__inv_2
X_16039_ _18084_/Q vssd1 vssd1 vccd1 vccd1 _16039_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16600__B _16600_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_238_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19729_ _20055_/CLK _19729_/D repeater207/X vssd1 vssd1 vccd1 vccd1 _19729_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17809__S1 _18752_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_226_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09413_ _19924_/Q vssd1 vssd1 vccd1 vccd1 _10040_/A sky130_fd_sc_hd__inv_2
XFILLER_241_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09344_ _20033_/Q vssd1 vssd1 vccd1 vccd1 _09493_/A sky130_fd_sc_hd__inv_2
XFILLER_178_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20012__CLK _20013_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09275_ _20054_/Q _09269_/X _09094_/X _09271_/X vssd1 vssd1 vccd1 vccd1 _20054_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_148_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_42_HCLK_A clkbuf_opt_2_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19408__RESET_B repeater193/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13384__B1 _20115_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09052__A1 _20108_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17593__S _17600_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10050_ _19935_/Q _10049_/Y _10022_/C _10049_/A _10026_/X vssd1 vssd1 vccd1 vccd1
+ _19935_/D sky130_fd_sc_hd__o221a_1
XANTENNA__11698__B1 _10866_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15407__A _15413_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_189_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16937__S _16946_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13740_ _17764_/X _13262_/B _13256_/X vssd1 vssd1 vccd1 vccd1 _13741_/B sky130_fd_sc_hd__a21oi_1
X_10952_ hold148/X _10948_/X _19669_/Q _10951_/X vssd1 vssd1 vccd1 vccd1 hold150/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_189_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13671_ _13671_/A vssd1 vssd1 vccd1 vccd1 _13671_/X sky130_fd_sc_hd__clkbuf_2
X_10883_ _19699_/Q _10875_/X _10882_/X _10879_/X vssd1 vssd1 vccd1 vccd1 _19699_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_32_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15410_ _18537_/Q _13224_/B _13225_/B vssd1 vssd1 vccd1 vccd1 _15410_/X sky130_fd_sc_hd__a21bo_1
XPHY_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_188_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12622_ _12629_/A vssd1 vssd1 vccd1 vccd1 _12622_/X sky130_fd_sc_hd__buf_1
XPHY_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16390_ _17344_/X _15900_/A _17318_/X _16234_/A vssd1 vssd1 vccd1 vccd1 _16390_/X
+ sky130_fd_sc_hd__o22a_2
XPHY_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_93_HCLK clkbuf_4_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19965_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_200_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15341_ _15347_/A _17598_/X vssd1 vssd1 vccd1 vccd1 _18492_/D sky130_fd_sc_hd__and2_1
XPHY_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12553_ _12553_/A _12556_/B vssd1 vssd1 vccd1 vccd1 _12553_/Y sky130_fd_sc_hd__nor2_1
XPHY_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14981__A hold237/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_196_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19831__RESET_B repeater271/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11504_ _11504_/A vssd1 vssd1 vccd1 vccd1 _11504_/X sky130_fd_sc_hd__clkbuf_2
X_18060_ _18460_/CLK _18060_/D vssd1 vssd1 vccd1 vccd1 _18060_/Q sky130_fd_sc_hd__dfxtp_1
X_15272_ _19722_/Q _19721_/Q vssd1 vssd1 vccd1 vccd1 _18479_/D sky130_fd_sc_hd__or2_1
XFILLER_156_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12484_ _19095_/Q _12478_/X _12236_/X _12479_/X vssd1 vssd1 vccd1 vccd1 _19095_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17011_ _17010_/X _11428_/Y _17548_/S vssd1 vssd1 vccd1 vccd1 _17011_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13597__A _13597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14223_ _18493_/Q _14223_/B vssd1 vssd1 vccd1 vccd1 _14224_/B sky130_fd_sc_hd__or2_1
X_11435_ _19137_/Q vssd1 vssd1 vccd1 vccd1 _11435_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11925__B2 _11892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11366_ _19129_/Q vssd1 vssd1 vccd1 vccd1 _11366_/Y sky130_fd_sc_hd__inv_2
X_14154_ _16717_/A _18701_/Q _19102_/Q _14012_/B _14153_/X vssd1 vssd1 vccd1 vccd1
+ _14166_/A sky130_fd_sc_hd__o221a_1
XFILLER_138_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13105_ _19165_/Q vssd1 vssd1 vccd1 vccd1 _13105_/Y sky130_fd_sc_hd__inv_2
X_10317_ _15716_/A _19868_/Q _19869_/Q vssd1 vssd1 vccd1 vccd1 _19868_/D sky130_fd_sc_hd__a21o_1
XFILLER_4_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14085_ _19062_/Q _14004_/A _19088_/Q _14029_/A vssd1 vssd1 vccd1 vccd1 _14085_/X
+ sky130_fd_sc_hd__o22a_1
X_11297_ _19580_/Q _11292_/Y _11468_/B _19001_/Q _11296_/X vssd1 vssd1 vccd1 vccd1
+ _11298_/D sky130_fd_sc_hd__o221a_1
X_18962_ _19208_/CLK _18962_/D repeater249/X vssd1 vssd1 vccd1 vccd1 _18962_/Q sky130_fd_sc_hd__dfrtp_4
X_10248_ _10954_/B vssd1 vssd1 vccd1 vccd1 _12053_/B sky130_fd_sc_hd__inv_2
X_17913_ _15794_/Y _15795_/Y _15796_/Y _15797_/Y _17913_/S0 _19632_/Q vssd1 vssd1
+ vccd1 vccd1 _17913_/X sky130_fd_sc_hd__mux4_2
X_13036_ _18910_/Q vssd1 vssd1 vccd1 vccd1 _13082_/A sky130_fd_sc_hd__inv_2
X_18893_ _18908_/CLK _18893_/D hold372/X vssd1 vssd1 vccd1 vccd1 _18893_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18784__RESET_B repeater267/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17008__S _17318_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11845__A _12372_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17844_ _17840_/X _17841_/X _17842_/X _17843_/X _19633_/Q _19634_/Q vssd1 vssd1 vccd1
+ vccd1 _17844_/X sky130_fd_sc_hd__mux4_2
XFILLER_227_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10179_ _19879_/Q _10174_/X _09105_/X _10175_/X vssd1 vssd1 vccd1 vccd1 _19879_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18713__RESET_B repeater252/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17775_ _18316_/Q _18436_/Q _18428_/Q _18420_/Q _17923_/S0 _19646_/Q vssd1 vssd1
+ vccd1 vccd1 _17775_/X sky130_fd_sc_hd__mux4_1
X_14987_ _18060_/Q _14978_/A hold263/X _14979_/A vssd1 vssd1 vccd1 vccd1 _18060_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16847__S _17488_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19514_ _19515_/CLK hold216/X repeater259/X vssd1 vssd1 vccd1 vccd1 _19514_/Q sky130_fd_sc_hd__dfrtp_1
X_16726_ _16790_/X _16594_/X _16795_/X _16595_/X vssd1 vssd1 vccd1 vccd1 _16728_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_208_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13938_ _13938_/A vssd1 vssd1 vccd1 vccd1 _13938_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19445_ _20058_/CLK _19445_/D repeater194/X vssd1 vssd1 vccd1 vccd1 _19445_/Q sky130_fd_sc_hd__dfrtp_1
X_16657_ _19084_/Q vssd1 vssd1 vccd1 vccd1 _16657_/Y sky130_fd_sc_hd__inv_2
X_13869_ _19197_/Q _13945_/A _19210_/Q _13910_/B vssd1 vssd1 vccd1 vccd1 _13869_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__19919__RESET_B repeater230/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15052__B1 _14998_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15608_ _18596_/Q vssd1 vssd1 vccd1 vccd1 _15608_/Y sky130_fd_sc_hd__inv_2
X_19376_ _19971_/CLK _19376_/D repeater241/X vssd1 vssd1 vccd1 vccd1 _19376_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_50_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16588_ _16588_/A _16615_/B vssd1 vssd1 vccd1 vccd1 _16588_/Y sky130_fd_sc_hd__nor2_1
XFILLER_222_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18327_ _19637_/CLK _18327_/D vssd1 vssd1 vccd1 vccd1 _18327_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17678__S _17696_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15539_ _18577_/Q _15530_/A _15530_/B _18578_/Q vssd1 vssd1 vccd1 vccd1 _15539_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_148_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09060_ hold282/X vssd1 vssd1 vccd1 vccd1 _12028_/A sky130_fd_sc_hd__buf_4
X_18258_ _18260_/CLK _18258_/D vssd1 vssd1 vccd1 vccd1 _18258_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17209_ _15768_/Y _11244_/Y _17546_/S vssd1 vssd1 vccd1 vccd1 _17209_/X sky130_fd_sc_hd__mux2_1
XFILLER_191_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18189_ _18216_/CLK _18189_/D vssd1 vssd1 vccd1 vccd1 _18189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09962_ _09871_/A _09871_/B _09960_/Y _09987_/B vssd1 vssd1 vccd1 vccd1 _19963_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_103_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13669__A1 _18779_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08913_ _20123_/Q vssd1 vssd1 vccd1 vccd1 _10133_/A sky130_fd_sc_hd__clkbuf_2
X_20082_ _20090_/CLK _20082_/D repeater204/X vssd1 vssd1 vccd1 vccd1 _20082_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_69_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09893_ _09876_/A _19360_/Q _19946_/Q _09892_/Y vssd1 vssd1 vccd1 vccd1 _09893_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_58_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_225_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15043__B1 _15004_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_241_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16791__A0 _15768_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17588__S _17600_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15897__A _15897_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09327_ _20043_/Q _15721_/A _09324_/Y _09325_/Y _09326_/Y vssd1 vssd1 vccd1 vccd1
+ _09327_/X sky130_fd_sc_hd__o221a_1
XFILLER_139_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09258_ _19516_/Q vssd1 vssd1 vccd1 vccd1 _10148_/A sky130_fd_sc_hd__inv_2
XFILLER_193_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19242__RESET_B repeater239/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09189_ _10133_/B _08983_/B _09188_/X vssd1 vssd1 vccd1 vccd1 _20073_/D sky130_fd_sc_hd__o21a_1
XFILLER_153_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11220_ _18999_/Q vssd1 vssd1 vccd1 vccd1 _11220_/Y sky130_fd_sc_hd__inv_2
XFILLER_153_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11151_ _19648_/Q _11053_/B _19648_/Q _11053_/B vssd1 vssd1 vccd1 vccd1 _11151_/X
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__16846__A1 _12929_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10102_ _10011_/B _10104_/A _10011_/A vssd1 vssd1 vccd1 vccd1 _10103_/B sky130_fd_sc_hd__o21a_1
X_11082_ _19058_/Q vssd1 vssd1 vccd1 vccd1 _12551_/A sky130_fd_sc_hd__inv_2
XFILLER_1_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10033_ _10081_/B _10033_/B vssd1 vssd1 vccd1 vccd1 _10034_/B sky130_fd_sc_hd__or2_2
X_14910_ _14910_/A vssd1 vssd1 vccd1 vccd1 _14910_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_209_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15890_ _15890_/A vssd1 vssd1 vccd1 vccd1 _16633_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_236_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_248_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input24_A HADDR[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14841_ _18147_/Q _14833_/A _14816_/X _14834_/A vssd1 vssd1 vccd1 vccd1 _18147_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_75_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17560_ _17559_/X _16750_/A _17565_/S vssd1 vssd1 vccd1 vccd1 _17560_/X sky130_fd_sc_hd__mux2_1
X_14772_ _14772_/A vssd1 vssd1 vccd1 vccd1 _14773_/A sky130_fd_sc_hd__inv_2
XFILLER_91_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11984_ _19369_/Q _11977_/X _11920_/X _11979_/X vssd1 vssd1 vccd1 vccd1 _19369_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_56_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16511_ _17298_/X _16508_/X _17284_/X _16235_/X _16510_/X vssd1 vssd1 vccd1 vccd1
+ _16511_/X sky130_fd_sc_hd__o221a_1
XANTENNA__17023__A1 _12952_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_205_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13723_ _13723_/A vssd1 vssd1 vccd1 vccd1 _14366_/A sky130_fd_sc_hd__clkbuf_2
X_10935_ _18508_/Q _15213_/A _10617_/B vssd1 vssd1 vccd1 vccd1 _10936_/S sky130_fd_sc_hd__o21ai_1
XFILLER_189_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17491_ _17490_/X _13846_/Y _17545_/S vssd1 vssd1 vccd1 vccd1 _17491_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_205_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_189_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19230_ _19282_/CLK _19230_/D repeater214/X vssd1 vssd1 vccd1 vccd1 _19230_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_204_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16442_ _16440_/Y _15828_/A _16441_/Y _16303_/X vssd1 vssd1 vccd1 vccd1 _16442_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_32_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13654_ _13654_/A vssd1 vssd1 vccd1 vccd1 _15169_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__16782__A0 _17473_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10866_ _13678_/A vssd1 vssd1 vccd1 vccd1 _10866_/X sky130_fd_sc_hd__buf_2
X_12605_ _19028_/Q _12598_/X _12536_/X _12600_/X vssd1 vssd1 vccd1 vccd1 _19028_/D
+ sky130_fd_sc_hd__a22o_1
X_19161_ _19968_/CLK _19161_/D hold370/X vssd1 vssd1 vccd1 vccd1 _19161_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16373_ _18483_/Q vssd1 vssd1 vccd1 vccd1 _16373_/Y sky130_fd_sc_hd__inv_2
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13585_ _13543_/A _13543_/B _13571_/X _13583_/Y vssd1 vssd1 vccd1 vccd1 _18820_/D
+ sky130_fd_sc_hd__a211oi_2
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10797_ _10797_/A vssd1 vssd1 vccd1 vccd1 _10797_/Y sky130_fd_sc_hd__inv_2
XFILLER_129_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18112_ _18137_/CLK _18112_/D vssd1 vssd1 vccd1 vccd1 _18112_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15324_ _15388_/A _15323_/Y _15216_/C _10907_/B _15204_/X vssd1 vssd1 vccd1 vccd1
+ _15325_/A sky130_fd_sc_hd__o32a_1
XPHY_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19092_ _19609_/CLK _19092_/D hold357/X vssd1 vssd1 vccd1 vccd1 _19092_/Q sky130_fd_sc_hd__dfrtp_4
X_12536_ hold331/X vssd1 vssd1 vccd1 vccd1 _12536_/X sky130_fd_sc_hd__buf_4
XFILLER_173_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18043_ _18954_/CLK _18043_/D vssd1 vssd1 vccd1 vccd1 _18043_/Q sky130_fd_sc_hd__dfxtp_1
X_15255_ _15250_/Y _15253_/Y _15254_/Y _18551_/Q vssd1 vssd1 vccd1 vccd1 _15286_/B
+ sky130_fd_sc_hd__a31o_1
X_12467_ _19108_/Q _12464_/X _12344_/X _12465_/X vssd1 vssd1 vccd1 vccd1 _19108_/D
+ sky130_fd_sc_hd__a22o_1
X_14206_ _19108_/Q _14017_/A _16583_/A _18689_/Q vssd1 vssd1 vccd1 vccd1 _14206_/X
+ sky130_fd_sc_hd__o22a_1
X_11418_ _19142_/Q vssd1 vssd1 vccd1 vccd1 _11418_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12020__B1 hold317/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15186_ _17933_/Q _14250_/X _10451_/A _14252_/X vssd1 vssd1 vccd1 vccd1 _17933_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_126_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12398_ hold298/X vssd1 vssd1 vccd1 vccd1 _12398_/X sky130_fd_sc_hd__buf_2
XANTENNA__18965__RESET_B hold370/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14137_ _14012_/B _14137_/A2 _18681_/Q _14136_/Y _14096_/X vssd1 vssd1 vccd1 vccd1
+ _18681_/D sky130_fd_sc_hd__o221a_1
XFILLER_126_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11349_ _11467_/A _18968_/Q _11483_/A _18985_/Q vssd1 vssd1 vccd1 vccd1 _11349_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_4_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19994_ _19997_/CLK _19994_/D repeater192/X vssd1 vssd1 vccd1 vccd1 _19994_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__14848__B1 _14802_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14068_ _19066_/Q vssd1 vssd1 vccd1 vccd1 _14068_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_100_HCLK clkbuf_4_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19222_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_101_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18945_ _18947_/CLK _18945_/D repeater211/X vssd1 vssd1 vccd1 vccd1 _18945_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_239_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13019_ _13019_/A vssd1 vssd1 vccd1 vccd1 _13023_/A sky130_fd_sc_hd__inv_2
XFILLER_239_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18876_ _20048_/CLK _18876_/D repeater208/X vssd1 vssd1 vccd1 vccd1 _18876_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_239_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09045__A hold301/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17827_ _18359_/Q _17999_/Q _18415_/Q _18399_/Q _17918_/S0 _18750_/Q vssd1 vssd1
+ vccd1 vccd1 _17827_/X sky130_fd_sc_hd__mux4_2
XFILLER_227_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12087__B1 _12086_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17758_ _17763_/S _13254_/Y _17764_/S vssd1 vssd1 vccd1 vccd1 _17758_/X sky130_fd_sc_hd__mux2_1
XFILLER_81_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11834__A0 _10147_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16709_ _19467_/Q vssd1 vssd1 vccd1 vccd1 _16709_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18508__D _18508_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17689_ _15476_/X _19446_/Q _17696_/S vssd1 vssd1 vccd1 vccd1 _18563_/D sky130_fd_sc_hd__mux2_1
XANTENNA__19753__RESET_B repeater196/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19428_ _19976_/CLK _19428_/D repeater185/X vssd1 vssd1 vccd1 vccd1 _19428_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_200_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19359_ _19970_/CLK _19359_/D repeater249/X vssd1 vssd1 vccd1 vccd1 _19359_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17201__S _17535_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09112_ _20088_/Q vssd1 vssd1 vccd1 vccd1 _09131_/A sky130_fd_sc_hd__inv_2
XFILLER_13_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09043_ _09043_/A vssd1 vssd1 vccd1 vccd1 _09043_/X sky130_fd_sc_hd__buf_1
XFILLER_163_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13030__A _18916_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12011__B1 _09030_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14839__B1 _14812_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13684__B _15169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09945_ _19970_/Q _09943_/Y _19963_/Q _16671_/A vssd1 vssd1 vccd1 vccd1 _09945_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_77_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20065_ _20066_/CLK _20065_/D repeater200/X vssd1 vssd1 vccd1 vccd1 _20065_/Q sky130_fd_sc_hd__dfrtp_1
X_09876_ _09876_/A _09954_/A vssd1 vssd1 vccd1 vccd1 _09877_/B sky130_fd_sc_hd__or2_1
XFILLER_161_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater260 repeater261/X vssd1 vssd1 vccd1 vccd1 repeater260/X sky130_fd_sc_hd__buf_8
Xrepeater271 repeater272/X vssd1 vssd1 vccd1 vccd1 repeater271/X sky130_fd_sc_hd__buf_8
XPHY_4403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater282 hold273/X vssd1 vssd1 vccd1 vccd1 repeater282/X sky130_fd_sc_hd__buf_6
XPHY_4414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11825__B1 _10861_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19494__RESET_B repeater260/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15016__B1 _15000_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13290__A2 _17918_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_199_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10720_ _10721_/A vssd1 vssd1 vccd1 vccd1 _10720_/X sky130_fd_sc_hd__buf_1
XPHY_3757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19423__RESET_B repeater274/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10651_ _19791_/Q _10651_/B vssd1 vssd1 vccd1 vccd1 _10652_/B sky130_fd_sc_hd__or2_1
XFILLER_13_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17111__S _17488_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10582_ _10582_/A _10939_/C vssd1 vssd1 vccd1 vccd1 _10583_/B sky130_fd_sc_hd__or2_1
X_13370_ _13369_/Y _18853_/Q _20107_/Q _13429_/D vssd1 vssd1 vccd1 vccd1 _13370_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_155_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12321_ _12335_/A vssd1 vssd1 vccd1 vccd1 _12321_/X sky130_fd_sc_hd__buf_1
XFILLER_5_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_186_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16950__S _16950_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15040_ _18031_/Q _15035_/X _14998_/X _15037_/X vssd1 vssd1 vccd1 vccd1 _18031_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_154_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12252_ _19225_/Q _15232_/A _12252_/S vssd1 vssd1 vccd1 vccd1 _19226_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_123_HCLK clkbuf_4_4_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19576_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_5_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11203_ _19605_/Q _11201_/Y _11459_/A _18992_/Q vssd1 vssd1 vccd1 vccd1 _11203_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_108_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12183_ _12187_/A _12183_/B vssd1 vssd1 vccd1 vccd1 _12184_/S sky130_fd_sc_hd__or2_1
XFILLER_123_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11134_ _12053_/B _15232_/C vssd1 vssd1 vccd1 vccd1 _12708_/C sky130_fd_sc_hd__or2_1
XFILLER_122_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16991_ _16649_/Y _19423_/Q _17487_/S vssd1 vssd1 vccd1 vccd1 _16991_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11065_ _11065_/A vssd1 vssd1 vccd1 vccd1 _15058_/A sky130_fd_sc_hd__clkbuf_2
X_18730_ _19224_/CLK _18730_/D repeater186/X vssd1 vssd1 vccd1 vccd1 _18730_/Q sky130_fd_sc_hd__dfrtp_4
X_15942_ _17946_/Q vssd1 vssd1 vccd1 vccd1 _15942_/Y sky130_fd_sc_hd__inv_2
XFILLER_135_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10016_ _10082_/A _10081_/C _10016_/C _10016_/D vssd1 vssd1 vccd1 vccd1 _10033_/B
+ sky130_fd_sc_hd__or4_4
XANTENNA__17244__A1 _20108_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18661_ _20048_/CLK _18661_/D repeater191/X vssd1 vssd1 vccd1 vccd1 _18661_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_48_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output130_A _18641_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15873_ _19328_/Q _15878_/B vssd1 vssd1 vccd1 vccd1 _15873_/Y sky130_fd_sc_hd__nor2_1
XFILLER_36_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17612_ _15232_/X _15222_/Y _17614_/S vssd1 vssd1 vccd1 vccd1 _17612_/X sky130_fd_sc_hd__mux2_1
XFILLER_76_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14824_ _18160_/Q _14820_/X _14749_/X _14822_/X vssd1 vssd1 vccd1 vccd1 _18160_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_224_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18592_ _19667_/CLK _18592_/D repeater264/X vssd1 vssd1 vccd1 vccd1 _18592_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_48_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17543_ _15863_/Y _14152_/Y _17543_/S vssd1 vssd1 vccd1 vccd1 _17543_/X sky130_fd_sc_hd__mux2_1
X_14755_ _18196_/Q _14746_/A _14727_/X _14747_/A vssd1 vssd1 vccd1 vccd1 _18196_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11816__B1 _09071_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11967_ _19379_/Q _11962_/X _09064_/X _11963_/X vssd1 vssd1 vccd1 vccd1 _19379_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__15007__B1 _15006_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13706_ _13706_/A _13706_/B vssd1 vssd1 vccd1 vccd1 _13707_/A sky130_fd_sc_hd__or2_1
X_10918_ _19681_/Q _10924_/A vssd1 vssd1 vccd1 vccd1 _10918_/X sky130_fd_sc_hd__or2_1
X_17474_ _17473_/X _15581_/A _17474_/S vssd1 vssd1 vccd1 vccd1 _17474_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14686_ _18232_/Q _14682_/X _14604_/X _14684_/X vssd1 vssd1 vccd1 vccd1 _18232_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_205_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11898_ _11914_/A vssd1 vssd1 vccd1 vccd1 _11898_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_220_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19213_ _19214_/CLK _19213_/D hold367/X vssd1 vssd1 vccd1 vccd1 _19213_/Q sky130_fd_sc_hd__dfrtp_4
X_16425_ _18137_/Q vssd1 vssd1 vccd1 vccd1 _16425_/Y sky130_fd_sc_hd__inv_2
X_13637_ _13637_/A _13637_/B vssd1 vssd1 vccd1 vccd1 _13637_/Y sky130_fd_sc_hd__nor2_1
XFILLER_220_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10849_ _19713_/Q _10843_/X _10418_/X _10845_/X vssd1 vssd1 vccd1 vccd1 _19713_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17021__S _17482_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19144_ _19566_/CLK _19144_/D repeater255/X vssd1 vssd1 vccd1 vccd1 _19144_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__20069__RESET_B repeater207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16356_ _18080_/Q vssd1 vssd1 vccd1 vccd1 _16356_/Y sky130_fd_sc_hd__inv_2
X_13568_ _13553_/A _13553_/B _13597_/A _13566_/Y vssd1 vssd1 vccd1 vccd1 _18830_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_118_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18120__CLK _18169_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15307_ _15289_/A _18519_/Q _15243_/Y _15306_/X vssd1 vssd1 vccd1 vccd1 _15307_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_200_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19075_ _19610_/CLK _19075_/D hold343/X vssd1 vssd1 vccd1 vccd1 _19075_/Q sky130_fd_sc_hd__dfrtp_4
X_12519_ _12528_/A vssd1 vssd1 vccd1 vccd1 _12519_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_200_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16287_ _17958_/Q vssd1 vssd1 vccd1 vccd1 _16287_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16860__S _17512_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13499_ _13620_/A vssd1 vssd1 vccd1 vccd1 _13499_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_246_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18026_ _19510_/CLK _18026_/D vssd1 vssd1 vccd1 vccd1 _18026_/Q sky130_fd_sc_hd__dfxtp_1
X_15238_ _18481_/Q _15237_/Y _18635_/Q _15229_/B _15334_/B vssd1 vssd1 vccd1 vccd1
+ _18635_/D sky130_fd_sc_hd__a221o_1
XFILLER_160_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15169_ _15169_/A _16115_/A vssd1 vssd1 vccd1 vccd1 _15171_/A sky130_fd_sc_hd__or2_2
XANTENNA__19396__CLK _20091_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19977_ _19984_/CLK _19977_/D repeater193/X vssd1 vssd1 vccd1 vccd1 _19977_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17691__S _17696_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09730_ _09848_/B vssd1 vssd1 vccd1 vccd1 _09731_/A sky130_fd_sc_hd__clkbuf_2
X_18928_ _19325_/CLK _18928_/D repeater213/X vssd1 vssd1 vccd1 vccd1 _18928_/Q sky130_fd_sc_hd__dfrtp_1
X_09661_ _19995_/Q vssd1 vssd1 vccd1 vccd1 _09751_/A sky130_fd_sc_hd__inv_2
X_18859_ _18866_/CLK _18859_/D repeater232/X vssd1 vssd1 vccd1 vccd1 _18859_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_95_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_228_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17988__CLK _19851_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09592_ _09592_/A vssd1 vssd1 vccd1 vccd1 _09592_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12480__B1 _12299_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_146_HCLK clkbuf_4_1_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19667_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_176_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18887__RESET_B repeater212/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16770__S _17493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18816__RESET_B repeater217/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09026_ _20119_/Q _09015_/X _09025_/X _09019_/X vssd1 vssd1 vccd1 vccd1 _20119_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_105_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold240 input40/X vssd1 vssd1 vccd1 vccd1 hold240/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold251 input39/X vssd1 vssd1 vccd1 vccd1 hold251/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 hold262/A vssd1 vssd1 vccd1 vccd1 hold262/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 hold273/A vssd1 vssd1 vccd1 vccd1 hold273/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold284 input62/X vssd1 vssd1 vccd1 vccd1 hold284/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 HWDATA[17] vssd1 vssd1 vccd1 vccd1 input46/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10831__B _10831_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18763__CLK _20123_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20117_ _20120_/CLK _20117_/D repeater217/X vssd1 vssd1 vccd1 vccd1 _20117_/Q sky130_fd_sc_hd__dfrtp_1
X_09928_ _09928_/A _09928_/B _09928_/C _09928_/D vssd1 vssd1 vccd1 vccd1 _09948_/C
+ sky130_fd_sc_hd__and4_1
XANTENNA__12104__A hold294/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20048_ _20048_/CLK _20048_/D repeater208/X vssd1 vssd1 vccd1 vccd1 _20048_/Q sky130_fd_sc_hd__dfrtp_1
X_09859_ _09859_/A _09859_/B vssd1 vssd1 vccd1 vccd1 _09981_/A sky130_fd_sc_hd__or2_1
XFILLER_246_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_234_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17106__S _17566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15415__A _15419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16985__A0 _17829_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12870_ _13007_/A _13006_/A _12870_/C _13008_/A vssd1 vssd1 vccd1 vccd1 _12871_/D
+ sky130_fd_sc_hd__or4_4
XFILLER_171_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11821_ _11821_/A vssd1 vssd1 vccd1 vccd1 _11821_/X sky130_fd_sc_hd__clkbuf_2
XPHY_4244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16945__S _16946_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14540_ _18317_/Q _14530_/X hold330/X _14533_/X vssd1 vssd1 vccd1 vccd1 _18317_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_242_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11752_ hold171/X _11750_/X _19490_/Q _11751_/X vssd1 vssd1 vccd1 vccd1 hold173/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_42_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_214_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10703_ _18879_/Q vssd1 vssd1 vccd1 vccd1 _15391_/A sky130_fd_sc_hd__inv_2
XPHY_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14471_ _18356_/Q _14464_/A _14419_/X _14465_/A vssd1 vssd1 vccd1 vccd1 _18356_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11683_ _11671_/X _11672_/Y _18627_/Q _19534_/Q _11666_/X vssd1 vssd1 vccd1 vccd1
+ _19534_/D sky130_fd_sc_hd__a32o_1
XPHY_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16210_ _16210_/A _16212_/B vssd1 vssd1 vccd1 vccd1 _16210_/Y sky130_fd_sc_hd__nor2_1
X_13422_ _18868_/Q _13355_/Y _13356_/Y _13355_/A _13421_/X vssd1 vssd1 vccd1 vccd1
+ _18868_/D sky130_fd_sc_hd__o221a_1
XPHY_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10634_ _19801_/Q _10606_/A _10594_/A _10609_/X vssd1 vssd1 vccd1 vccd1 _19801_/D
+ sky130_fd_sc_hd__a22o_1
X_17190_ _17189_/X _13879_/Y _17545_/S vssd1 vssd1 vccd1 vccd1 _17190_/X sky130_fd_sc_hd__mux2_1
XPHY_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16141_ _17428_/X vssd1 vssd1 vccd1 vccd1 _16141_/Y sky130_fd_sc_hd__inv_2
X_13353_ _18866_/Q _13435_/A vssd1 vssd1 vccd1 vccd1 _13354_/B sky130_fd_sc_hd__nand2_2
X_10565_ _10614_/C _10613_/C vssd1 vssd1 vccd1 vccd1 _15334_/C sky130_fd_sc_hd__nor2_1
XANTENNA__18557__RESET_B repeater193/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12304_ _19197_/Q _12298_/X _12232_/X _12300_/X vssd1 vssd1 vccd1 vccd1 _19197_/D
+ sky130_fd_sc_hd__a22o_1
X_16072_ _17448_/X _16069_/X _17445_/X _16070_/X _16071_/X vssd1 vssd1 vccd1 vccd1
+ _16072_/X sky130_fd_sc_hd__o221a_1
X_13284_ _13284_/A vssd1 vssd1 vccd1 vccd1 _13285_/B sky130_fd_sc_hd__buf_1
X_10496_ _19541_/Q vssd1 vssd1 vccd1 vccd1 _10732_/B sky130_fd_sc_hd__inv_2
XANTENNA__12526__A1 _19069_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15023_ _15024_/A vssd1 vssd1 vccd1 vccd1 _15023_/X sky130_fd_sc_hd__clkbuf_2
X_19900_ _19900_/CLK _19900_/D repeater195/X vssd1 vssd1 vccd1 vccd1 _19900_/Q sky130_fd_sc_hd__dfrtp_1
X_12235_ _19230_/Q _12228_/X _12234_/X _12229_/X vssd1 vssd1 vccd1 vccd1 _19230_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17465__A1 _08941_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19831_ _20058_/CLK _19831_/D repeater271/X vssd1 vssd1 vccd1 vccd1 _19831_/Q sky130_fd_sc_hd__dfrtp_4
X_12166_ _19273_/Q _12164_/X _12035_/X _12165_/X vssd1 vssd1 vccd1 vccd1 _19273_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11837__B _15839_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11117_ _11094_/Y _11113_/B _11116_/Y _17755_/X _11110_/Y vssd1 vssd1 vccd1 vccd1
+ _11118_/A sky130_fd_sc_hd__o32a_1
X_19762_ _19772_/CLK _19762_/D repeater218/X vssd1 vssd1 vccd1 vccd1 _19762_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_19_HCLK_A clkbuf_4_3_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16974_ _16973_/X _13550_/A _17536_/S vssd1 vssd1 vccd1 vccd1 _16974_/X sky130_fd_sc_hd__mux2_2
X_12097_ _19315_/Q _12094_/X _12095_/X _12096_/X vssd1 vssd1 vccd1 vccd1 _19315_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_1_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17217__A1 _12919_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_27_HCLK clkbuf_4_9_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20055_/CLK sky130_fd_sc_hd__clkbuf_16
X_18713_ _18718_/CLK _18713_/D repeater252/X vssd1 vssd1 vccd1 vccd1 _18713_/Q sky130_fd_sc_hd__dfrtp_1
X_11048_ _11056_/A _14301_/B vssd1 vssd1 vccd1 vccd1 _11049_/A sky130_fd_sc_hd__or2_1
X_15925_ _18035_/Q vssd1 vssd1 vccd1 vccd1 _15925_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19693_ _20049_/CLK _19693_/D repeater208/X vssd1 vssd1 vccd1 vccd1 _19693_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_7_HCLK_A clkbuf_4_2_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput8 input8/A vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__clkbuf_1
XFILLER_92_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17016__S _17490_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15856_ _15753_/A _15854_/X _15855_/Y _15842_/X vssd1 vssd1 vccd1 vccd1 _15856_/X
+ sky130_fd_sc_hd__o22a_1
X_18644_ _20059_/CLK _18644_/D repeater197/X vssd1 vssd1 vccd1 vccd1 _18644_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__19345__RESET_B repeater245/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14807_ _18168_/Q _14801_/X _14806_/X _14804_/X vssd1 vssd1 vccd1 vccd1 _18168_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_224_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15787_ _18066_/Q vssd1 vssd1 vccd1 vccd1 _15787_/Y sky130_fd_sc_hd__inv_2
X_18575_ _19462_/CLK _18575_/D repeater273/X vssd1 vssd1 vccd1 vccd1 _18575_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__16855__S _17523_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12999_ _12965_/C _12873_/B _12997_/Y _12986_/X vssd1 vssd1 vccd1 vccd1 _18931_/D
+ sky130_fd_sc_hd__a211oi_2
X_17526_ _17525_/X _09815_/Y _17548_/S vssd1 vssd1 vccd1 vccd1 _17526_/X sky130_fd_sc_hd__mux2_1
X_14738_ _18206_/Q _14732_/X _14723_/X _14734_/X vssd1 vssd1 vccd1 vccd1 _18206_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12462__B1 _12408_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17457_ _17456_/X _13858_/Y _17545_/S vssd1 vssd1 vccd1 vccd1 _17457_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14669_ _14670_/A vssd1 vssd1 vccd1 vccd1 _14669_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_189_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12684__A _12698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16408_ _18153_/Q vssd1 vssd1 vccd1 vccd1 _16408_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18636__CLK _19780_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12214__B1 _12107_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17388_ _17387_/X _18891_/Q _17488_/S vssd1 vssd1 vccd1 vccd1 _17388_/X sky130_fd_sc_hd__mux2_2
XFILLER_146_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17686__S _17696_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19127_ _19576_/CLK _19127_/D repeater255/X vssd1 vssd1 vccd1 vccd1 _19127_/Q sky130_fd_sc_hd__dfrtp_1
X_16339_ _18352_/Q vssd1 vssd1 vccd1 vccd1 _16339_/Y sky130_fd_sc_hd__inv_2
X_19058_ _19630_/CLK _19058_/D repeater257/X vssd1 vssd1 vccd1 vccd1 _19058_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__16900__A0 _17473_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18009_ _18416_/CLK _18009_/D vssd1 vssd1 vccd1 vccd1 _18009_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_160_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11740__A2 _11737_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09713_ _09705_/X _09713_/B _09713_/C _09713_/D vssd1 vssd1 vccd1 vccd1 _09728_/C
+ sky130_fd_sc_hd__and4b_1
XFILLER_228_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09644_ _19983_/Q vssd1 vssd1 vccd1 vccd1 _09646_/C sky130_fd_sc_hd__inv_2
XANTENNA__19086__RESET_B hold351/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18166__CLK _18169_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09575_ _20031_/Q _09574_/Y _09567_/X _09492_/B vssd1 vssd1 vccd1 vccd1 _20031_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__16765__S _17386_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19411__CLK _19984_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12453__B1 _12392_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17596__S _17600_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17144__A0 _15963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16498__A2 _15898_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10350_ _10344_/B _10320_/X _10349_/Y _10345_/X _10329_/A vssd1 vssd1 vccd1 vccd1
+ _10351_/A sky130_fd_sc_hd__o32a_1
XFILLER_191_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12508__A1 _19081_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17790__S1 _19646_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09009_ _19510_/Q _19509_/Q _19512_/Q _19511_/Q vssd1 vssd1 vccd1 vccd1 _09010_/D
+ sky130_fd_sc_hd__or4_4
XANTENNA__11938__A _11977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10281_ _10281_/A _10281_/B _10281_/C _11150_/C vssd1 vssd1 vccd1 vccd1 _10281_/X
+ sky130_fd_sc_hd__or4b_4
XFILLER_124_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10842__A _10842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14314__A _14405_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12020_ _19350_/Q _12016_/X hold317/X _12017_/X vssd1 vssd1 vccd1 vccd1 _19350_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_104_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13971_ _13964_/A _13964_/B _18704_/Q _13913_/X _13907_/X vssd1 vssd1 vccd1 vccd1
+ _18704_/D sky130_fd_sc_hd__o221a_1
XFILLER_74_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15710_ _15710_/A _15713_/B vssd1 vssd1 vccd1 vccd1 _18645_/D sky130_fd_sc_hd__nor2_1
XFILLER_76_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12922_ _19264_/Q vssd1 vssd1 vccd1 vccd1 _12922_/Y sky130_fd_sc_hd__inv_1
X_16690_ _17011_/X _16687_/X _17058_/X _16688_/X _16689_/X vssd1 vssd1 vccd1 vccd1
+ _16691_/C sky130_fd_sc_hd__o221a_1
XFILLER_58_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15641_ _15649_/C vssd1 vssd1 vccd1 vccd1 _15641_/Y sky130_fd_sc_hd__inv_2
X_12853_ _18931_/Q vssd1 vssd1 vccd1 vccd1 _12965_/C sky130_fd_sc_hd__inv_2
XPHY_4030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_234_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18360_ _19849_/CLK _18360_/D vssd1 vssd1 vccd1 vccd1 _18360_/Q sky130_fd_sc_hd__dfxtp_1
X_11804_ _19458_/Q _11800_/X hold317/X _11801_/X vssd1 vssd1 vccd1 vccd1 _19458_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11247__B2 _19009_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15572_ _18587_/Q vssd1 vssd1 vccd1 vccd1 _15572_/Y sky130_fd_sc_hd__inv_2
X_12784_ _18825_/Q vssd1 vssd1 vccd1 vccd1 _13548_/A sky130_fd_sc_hd__inv_2
XPHY_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_221_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17311_ _16435_/Y _17839_/X _17568_/S vssd1 vssd1 vccd1 vccd1 _17311_/X sky130_fd_sc_hd__mux2_2
XANTENNA__19904__CLK _20123_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14523_ _18327_/Q _14518_/X _14443_/X _14520_/X vssd1 vssd1 vccd1 vccd1 _18327_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18291_ _19873_/CLK _18291_/D vssd1 vssd1 vccd1 vccd1 _18291_/Q sky130_fd_sc_hd__dfxtp_1
X_11735_ _19502_/Q _11730_/X _16934_/X _11731_/X vssd1 vssd1 vccd1 vccd1 hold229/A
+ sky130_fd_sc_hd__a22o_1
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17242_ _17241_/X _14038_/Y _17490_/S vssd1 vssd1 vccd1 vccd1 _17242_/X sky130_fd_sc_hd__mux2_2
XFILLER_30_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14454_ _18369_/Q _14451_/X _14437_/X _14453_/X vssd1 vssd1 vccd1 vccd1 _18369_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11666_ _11668_/A vssd1 vssd1 vccd1 vccd1 _11666_/X sky130_fd_sc_hd__clkbuf_2
XPHY_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13405_ _13403_/Y _18849_/Q _20103_/Q _13428_/D _13404_/X vssd1 vssd1 vccd1 vccd1
+ _13405_/X sky130_fd_sc_hd__a221o_1
XPHY_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10617_ _10617_/A _10617_/B vssd1 vssd1 vccd1 vccd1 _10617_/X sky130_fd_sc_hd__or2_2
X_17173_ _17486_/A0 _13128_/Y _17543_/S vssd1 vssd1 vccd1 vccd1 _17173_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14385_ _18407_/Q _14380_/X _12720_/X _14382_/X vssd1 vssd1 vccd1 vccd1 _18407_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_repeater243_A repeater244/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11597_ _11597_/A vssd1 vssd1 vccd1 vccd1 _11597_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12009__A _12016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16124_ _19712_/Q vssd1 vssd1 vccd1 vccd1 _16124_/Y sky130_fd_sc_hd__inv_2
X_13336_ _13428_/D _13336_/B vssd1 vssd1 vccd1 vccd1 _13459_/A sky130_fd_sc_hd__or2_1
X_10548_ _19809_/Q _10939_/D vssd1 vssd1 vccd1 vccd1 _10567_/D sky130_fd_sc_hd__or2_1
XFILLER_227_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16055_ _16055_/A vssd1 vssd1 vccd1 vccd1 _16055_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__17781__S1 _19646_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15161__A2 _15158_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18039__CLK _19851_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13267_ _18753_/Q vssd1 vssd1 vccd1 vccd1 _14270_/B sky130_fd_sc_hd__clkbuf_2
X_10479_ _17703_/X _10471_/A _19816_/Q _10472_/A vssd1 vssd1 vccd1 vccd1 _19816_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_142_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17438__A1 _17884_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15006_ _18953_/Q vssd1 vssd1 vccd1 vccd1 _15006_/X sky130_fd_sc_hd__buf_2
X_12218_ _19239_/Q _12212_/X _12032_/X _12213_/X vssd1 vssd1 vccd1 vccd1 _19239_/D
+ sky130_fd_sc_hd__a22o_1
X_13198_ _13069_/B _13198_/A2 _13069_/A vssd1 vssd1 vccd1 vccd1 _13199_/C sky130_fd_sc_hd__o21a_1
XFILLER_243_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19814_ _19814_/CLK _19814_/D repeater220/X vssd1 vssd1 vccd1 vccd1 _19814_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA_clkbuf_leaf_143_HCLK_A clkbuf_4_1_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12149_ _19284_/Q _12143_/X _12092_/X _12144_/X vssd1 vssd1 vccd1 vccd1 _19284_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_111_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19745_ _20070_/CLK _19745_/D repeater205/X vssd1 vssd1 vccd1 vccd1 _19745_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_238_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16957_ _17799_/X _18795_/Q _16957_/S vssd1 vssd1 vccd1 vccd1 _16957_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15908_ _15908_/A vssd1 vssd1 vccd1 vccd1 _15908_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_110_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19676_ _19794_/CLK _19676_/D repeater201/X vssd1 vssd1 vccd1 vccd1 _19676_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12683__B1 hold294/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16888_ _16887_/X _15703_/Y _17474_/S vssd1 vssd1 vccd1 vccd1 _16888_/X sky130_fd_sc_hd__mux2_1
XFILLER_237_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09053__A _09084_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18627_ _19545_/CLK _18627_/D repeater221/X vssd1 vssd1 vccd1 vccd1 _18627_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_25_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15839_ _15839_/A vssd1 vssd1 vccd1 vccd1 _15840_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_53_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_206_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09360_ _20017_/Q vssd1 vssd1 vccd1 vccd1 _09477_/A sky130_fd_sc_hd__inv_2
XANTENNA__20084__RESET_B repeater204/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12435__B1 _12241_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18558_ _20064_/CLK _18558_/D repeater193/X vssd1 vssd1 vccd1 vccd1 _18558_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_178_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17509_ _15881_/Y _15610_/A _17537_/S vssd1 vssd1 vccd1 vccd1 _17509_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09291_ _20046_/Q _09285_/X _09086_/X _09287_/X vssd1 vssd1 vccd1 vccd1 _20046_/D
+ sky130_fd_sc_hd__a22o_1
X_18489_ _19545_/CLK _18489_/D repeater225/X vssd1 vssd1 vccd1 vccd1 _18489_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_20_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12738__B2 _18821_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10749__B1 _10423_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11758__A _11772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17772__S1 _19646_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10662__A _10676_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput120 _16751_/X vssd1 vssd1 vccd1 vccd1 IRQ[2] sky130_fd_sc_hd__clkbuf_2
XANTENNA__15152__A2 _15146_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput131 _18642_/Q vssd1 vssd1 vccd1 vccd1 RsTx_S1 sky130_fd_sc_hd__clkbuf_2
Xoutput142 _16761_/LO vssd1 vssd1 vccd1 vccd1 sda_o_S4 sky130_fd_sc_hd__clkbuf_2
XFILLER_161_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11174__B1 _18879_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13973__A _18701_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19267__RESET_B repeater212/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_233_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_65_HCLK_A clkbuf_opt_4_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12674__B1 hold306/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_243_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_hold169_A HADDR[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18801__CLK _19900_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20091__CLK _20091_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09627_ _20000_/Q vssd1 vssd1 vccd1 vccd1 _09629_/A sky130_fd_sc_hd__inv_2
XFILLER_243_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09558_ _09471_/A _19300_/Q _09480_/A _19310_/Q _09557_/X vssd1 vssd1 vccd1 vccd1
+ _09564_/C sky130_fd_sc_hd__o221a_1
XANTENNA__12426__B1 _12296_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09489_ _09489_/A _09577_/A vssd1 vssd1 vccd1 vccd1 _09490_/B sky130_fd_sc_hd__or2_2
XPHY_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14179__B1 _16617_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11520_ _11520_/A vssd1 vssd1 vccd1 vccd1 _11520_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11451_ _19556_/Q vssd1 vssd1 vccd1 vccd1 _11626_/A sky130_fd_sc_hd__inv_2
XPHY_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10402_ _14477_/B _10396_/Y _10400_/X vssd1 vssd1 vccd1 vccd1 _19850_/D sky130_fd_sc_hd__o21a_1
X_14170_ _19111_/Q _14020_/A _19121_/Q _14030_/A _14169_/X vssd1 vssd1 vccd1 vccd1
+ _14184_/A sky130_fd_sc_hd__o221a_1
X_11382_ _19558_/Q _11380_/Y _19551_/Q _11381_/Y vssd1 vssd1 vccd1 vccd1 _11382_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_164_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13121_ _19158_/Q _13060_/A _13118_/Y _18906_/Q _13120_/X vssd1 vssd1 vccd1 vccd1
+ _13127_/C sky130_fd_sc_hd__o221a_1
X_10333_ _18766_/Q vssd1 vssd1 vccd1 vccd1 _10354_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_194_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13154__A1 _19166_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13052_ _18894_/Q vssd1 vssd1 vccd1 vccd1 _13067_/A sky130_fd_sc_hd__inv_2
X_10264_ _19646_/Q vssd1 vssd1 vccd1 vccd1 _10266_/A sky130_fd_sc_hd__inv_2
X_12003_ _12017_/A vssd1 vssd1 vccd1 vccd1 _12003_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_78_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10195_ _13635_/A _13637_/A _10195_/C vssd1 vssd1 vccd1 vccd1 _10196_/B sky130_fd_sc_hd__or3_1
X_17860_ _16252_/Y _16253_/Y _16254_/Y _16255_/Y _17913_/S0 _19632_/Q vssd1 vssd1
+ vccd1 vccd1 _17860_/X sky130_fd_sc_hd__mux4_2
XFILLER_120_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16811_ _16810_/X _14084_/Y _17490_/S vssd1 vssd1 vccd1 vccd1 _16811_/X sky130_fd_sc_hd__mux2_2
XFILLER_93_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17791_ _18391_/Q _18383_/Q _18375_/Q _18367_/Q _17923_/S0 _19646_/Q vssd1 vssd1
+ vccd1 vccd1 _17791_/X sky130_fd_sc_hd__mux4_2
XFILLER_120_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19530_ _19544_/CLK _19530_/D repeater221/X vssd1 vssd1 vccd1 vccd1 _19530_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_235_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16742_ _17063_/X _15904_/X _16888_/X _16235_/X _16741_/X vssd1 vssd1 vccd1 vccd1
+ _16743_/C sky130_fd_sc_hd__o221a_1
X_13954_ _13954_/A vssd1 vssd1 vccd1 vccd1 _13954_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12665__B1 hold284/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12905_ _19278_/Q vssd1 vssd1 vccd1 vccd1 _12905_/Y sky130_fd_sc_hd__inv_2
XFILLER_246_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16673_ _19049_/Q _16673_/B vssd1 vssd1 vccd1 vccd1 _16673_/Y sky130_fd_sc_hd__nand2_1
X_19461_ _19470_/CLK _19461_/D repeater273/X vssd1 vssd1 vccd1 vccd1 _19461_/Q sky130_fd_sc_hd__dfrtp_1
X_13885_ _13863_/Y _18704_/Q _19207_/Q _13911_/B _13884_/X vssd1 vssd1 vccd1 vccd1
+ _13885_/X sky130_fd_sc_hd__a221o_1
XFILLER_234_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18412_ _18412_/CLK _18412_/D vssd1 vssd1 vccd1 vccd1 _18412_/Q sky130_fd_sc_hd__dfxtp_1
X_12836_ _18951_/Q _13597_/A _12733_/Y vssd1 vssd1 vccd1 vccd1 _18951_/D sky130_fd_sc_hd__o21a_1
X_15624_ _18600_/Q vssd1 vssd1 vccd1 vccd1 _15624_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12417__B1 hold281/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19392_ _19933_/CLK _19392_/D repeater235/X vssd1 vssd1 vccd1 vccd1 _19392_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_222_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15555_ _18582_/Q _15555_/B vssd1 vssd1 vccd1 vccd1 _15556_/A sky130_fd_sc_hd__or2_1
X_18343_ _18954_/CLK _18343_/D vssd1 vssd1 vccd1 vccd1 _18343_/Q sky130_fd_sc_hd__dfxtp_1
X_12767_ _19253_/Q vssd1 vssd1 vccd1 vccd1 _12767_/Y sky130_fd_sc_hd__inv_2
XPHY_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14506_ _18337_/Q _14503_/X _14437_/X _14505_/X vssd1 vssd1 vccd1 vccd1 _18337_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13123__A _19168_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18274_ _19873_/CLK _18274_/D vssd1 vssd1 vccd1 vccd1 _18274_/Q sky130_fd_sc_hd__dfxtp_1
X_11718_ _19515_/Q _11716_/X _16947_/X _11717_/X vssd1 vssd1 vccd1 vccd1 hold226/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_42_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15486_ _15486_/A vssd1 vssd1 vccd1 vccd1 _15491_/B sky130_fd_sc_hd__inv_2
X_12698_ _12698_/A vssd1 vssd1 vccd1 vccd1 _12698_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__15906__B2 _15898_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18501__RESET_B repeater219/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14437_ _14745_/A vssd1 vssd1 vccd1 vccd1 _14437_/X sky130_fd_sc_hd__clkbuf_2
X_17225_ _17224_/X _13852_/Y _17545_/S vssd1 vssd1 vccd1 vccd1 _17225_/X sky130_fd_sc_hd__mux2_1
XFILLER_238_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11649_ _11649_/A _11649_/B vssd1 vssd1 vccd1 vccd1 _15271_/C sky130_fd_sc_hd__or2_1
Xinput11 input11/A vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__clkbuf_1
XFILLER_156_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput22 HADDR[29] vssd1 vssd1 vccd1 vccd1 input22/X sky130_fd_sc_hd__buf_1
XPHY_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput33 HREADY vssd1 vssd1 vccd1 vccd1 input33/X sky130_fd_sc_hd__buf_1
X_17156_ _15963_/X _12786_/Y _17534_/S vssd1 vssd1 vccd1 vccd1 _17156_/X sky130_fd_sc_hd__mux2_1
Xinput44 input44/A vssd1 vssd1 vccd1 vccd1 input44/X sky130_fd_sc_hd__buf_1
Xinput55 input55/A vssd1 vssd1 vccd1 vccd1 input55/X sky130_fd_sc_hd__clkbuf_4
X_14368_ _14368_/A vssd1 vssd1 vccd1 vccd1 _14369_/A sky130_fd_sc_hd__inv_2
Xinput66 input66/A vssd1 vssd1 vccd1 vccd1 input66/X sky130_fd_sc_hd__buf_4
Xinput77 input77/A vssd1 vssd1 vccd1 vccd1 input77/X sky130_fd_sc_hd__clkbuf_1
XFILLER_143_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16107_ _18261_/Q vssd1 vssd1 vccd1 vccd1 _16107_/Y sky130_fd_sc_hd__inv_2
X_13319_ _18840_/Q vssd1 vssd1 vccd1 vccd1 _13322_/A sky130_fd_sc_hd__clkinv_1
XFILLER_182_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17087_ _15768_/Y _11201_/Y _17546_/S vssd1 vssd1 vccd1 vccd1 _17087_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14299_ _14598_/B vssd1 vssd1 vccd1 vccd1 _14450_/B sky130_fd_sc_hd__buf_1
XFILLER_170_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14342__B1 hold324/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16038_ _17955_/Q vssd1 vssd1 vccd1 vccd1 _16038_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10903__B1 _10870_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17989_ _18165_/CLK _17989_/D vssd1 vssd1 vccd1 vccd1 _17989_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_245_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19728_ _20055_/CLK _19728_/D repeater207/X vssd1 vssd1 vccd1 vccd1 _19728_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12656__B1 _12538_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_238_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19659_ _19846_/CLK _19659_/D repeater270/X vssd1 vssd1 vccd1 vccd1 _19659_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_65_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17204__S _17529_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09412_ _10011_/B _09411_/Y _19908_/Q _19368_/Q vssd1 vssd1 vccd1 vccd1 _09416_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_25_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09343_ _20034_/Q vssd1 vssd1 vccd1 vccd1 _09494_/A sky130_fd_sc_hd__inv_2
XFILLER_178_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17347__A0 _17473_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_221_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09274_ _20055_/Q _09269_/X _09090_/X _09271_/X vssd1 vssd1 vccd1 vccd1 _20055_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_139_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_178_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16322__A1 _17356_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09760__B1 _09759_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08989_ _10819_/A vssd1 vssd1 vccd1 vccd1 _11830_/A sky130_fd_sc_hd__inv_2
XFILLER_102_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12647__B1 hold267/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10951_ _11772_/A vssd1 vssd1 vccd1 vccd1 _10951_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_243_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17114__S _17566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13670_ _18778_/Q _13664_/X _12599_/X _13665_/X vssd1 vssd1 vccd1 vccd1 _18778_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_71_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10882_ _14277_/A vssd1 vssd1 vccd1 vccd1 _10882_/X sky130_fd_sc_hd__buf_4
XFILLER_243_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12621_ _19019_/Q _12613_/X _12386_/X _12616_/X vssd1 vssd1 vccd1 vccd1 _19019_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15340_ _18492_/Q _14222_/B _14223_/B vssd1 vssd1 vccd1 vccd1 _15340_/X sky130_fd_sc_hd__a21bo_1
XPHY_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12552_ _11085_/C _12551_/X _12548_/Y vssd1 vssd1 vccd1 vccd1 _19059_/D sky130_fd_sc_hd__a21oi_1
XPHY_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11503_ _11503_/A vssd1 vssd1 vccd1 vccd1 _11503_/Y sky130_fd_sc_hd__inv_2
XPHY_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15271_ _15271_/A _15271_/B _15271_/C _15271_/D vssd1 vssd1 vccd1 vccd1 _15271_/X
+ sky130_fd_sc_hd__or4_4
XPHY_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13878__A _19210_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12483_ _19096_/Q _12478_/X _12234_/X _12479_/X vssd1 vssd1 vccd1 vccd1 _19096_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17010_ _17009_/X _16679_/Y _17493_/S vssd1 vssd1 vccd1 vccd1 _17010_/X sky130_fd_sc_hd__mux2_1
X_14222_ _18492_/Q _14222_/B vssd1 vssd1 vccd1 vccd1 _14223_/B sky130_fd_sc_hd__or2_1
XPHY_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11434_ _19557_/Q vssd1 vssd1 vccd1 vccd1 _11551_/C sky130_fd_sc_hd__inv_2
XFILLER_171_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19871__RESET_B repeater207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11925__A2 _11891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14153_ _19099_/Q _14009_/A _14152_/Y _18672_/Q vssd1 vssd1 vccd1 vccd1 _14153_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_164_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11365_ _11223_/X _11248_/X _11299_/X _19610_/Q _11504_/A vssd1 vssd1 vccd1 vccd1
+ _19610_/D sky130_fd_sc_hd__a32o_1
XFILLER_98_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19800__RESET_B repeater222/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18847__CLK _18866_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13104_ _13101_/Y _18914_/Q _19172_/Q _13073_/A _13103_/X vssd1 vssd1 vccd1 vccd1
+ _13109_/C sky130_fd_sc_hd__o221a_1
X_10316_ _19869_/Q _10290_/B _10291_/X vssd1 vssd1 vccd1 vccd1 _19869_/D sky130_fd_sc_hd__o21a_1
X_18961_ _19600_/CLK _18961_/D hold273/X vssd1 vssd1 vccd1 vccd1 _18961_/Q sky130_fd_sc_hd__dfrtp_4
X_14084_ _19082_/Q vssd1 vssd1 vccd1 vccd1 _14084_/Y sky130_fd_sc_hd__inv_2
X_11296_ _19587_/Q _11294_/Y _19607_/Q _16716_/A vssd1 vssd1 vccd1 vccd1 _11296_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_4_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17912_ _15790_/Y _15791_/Y _15792_/Y _15793_/Y _17913_/S0 _19632_/Q vssd1 vssd1
+ vccd1 vccd1 _17912_/X sky130_fd_sc_hd__mux4_1
X_13035_ _18911_/Q vssd1 vssd1 vccd1 vccd1 _13083_/A sky130_fd_sc_hd__inv_2
X_10247_ _10209_/X _10247_/B _10247_/C _10247_/D vssd1 vssd1 vccd1 vccd1 _10954_/B
+ sky130_fd_sc_hd__and4b_4
X_18892_ _19968_/CLK _18892_/D hold372/X vssd1 vssd1 vccd1 vccd1 _18892_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_repeater206_A repeater207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_239_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17843_ _16410_/Y _16411_/Y _16412_/Y _16413_/Y _17913_/S0 _19632_/Q vssd1 vssd1
+ vccd1 vccd1 _17843_/X sky130_fd_sc_hd__mux4_2
XFILLER_66_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10178_ _19880_/Q _10174_/X _09101_/X _10175_/X vssd1 vssd1 vccd1 vccd1 _19880_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_227_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17774_ _17770_/X _17771_/X _17772_/X _17773_/X _19647_/Q _19648_/Q vssd1 vssd1 vccd1
+ vccd1 _17774_/X sky130_fd_sc_hd__mux4_2
XANTENNA__12638__B1 _12413_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14986_ _18061_/Q _14976_/X _14793_/X _14979_/X vssd1 vssd1 vccd1 vccd1 _18061_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_82_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19513_ _19513_/CLK hold224/X repeater259/X vssd1 vssd1 vccd1 vccd1 _19513_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_75_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16725_ _16781_/X _16555_/A _16831_/X _16556_/A vssd1 vssd1 vccd1 vccd1 _16728_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_235_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13937_ _13910_/D _13819_/B _13935_/Y _13927_/X vssd1 vssd1 vccd1 vccd1 _18720_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_34_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15333__A _15333_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18753__RESET_B repeater195/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17024__S _17542_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19444_ _20058_/CLK _19444_/D repeater198/X vssd1 vssd1 vccd1 vccd1 _19444_/Q sky130_fd_sc_hd__dfrtp_1
X_16656_ _16656_/A _16656_/B _16656_/C _16656_/D vssd1 vssd1 vccd1 vccd1 _16656_/X
+ sky130_fd_sc_hd__or4_4
X_13868_ _19221_/Q vssd1 vssd1 vccd1 vccd1 _13868_/Y sky130_fd_sc_hd__inv_2
XFILLER_223_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12819_ _19228_/Q _13529_/A _19254_/Q _13554_/A vssd1 vssd1 vccd1 vccd1 _12819_/X
+ sky130_fd_sc_hd__o22a_1
X_15607_ _15605_/Y _15606_/Y _15590_/X vssd1 vssd1 vccd1 vccd1 _15607_/X sky130_fd_sc_hd__o21a_1
X_19375_ _19971_/CLK _19375_/D repeater191/X vssd1 vssd1 vccd1 vccd1 _19375_/Q sky130_fd_sc_hd__dfrtp_1
X_16587_ _16587_/A _16615_/B vssd1 vssd1 vccd1 vccd1 _16587_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__16863__S _17318_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13799_ _18707_/Q vssd1 vssd1 vccd1 vccd1 _13802_/A sky130_fd_sc_hd__inv_2
XFILLER_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18326_ _19637_/CLK _18326_/D vssd1 vssd1 vccd1 vccd1 _18326_/Q sky130_fd_sc_hd__dfxtp_1
X_15538_ _15538_/A vssd1 vssd1 vccd1 vccd1 _15538_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19622__CLK _19920_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15469_ _18562_/Q vssd1 vssd1 vccd1 vccd1 _15471_/A sky130_fd_sc_hd__inv_2
X_18257_ _20077_/CLK _18257_/D vssd1 vssd1 vccd1 vccd1 _18257_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12692__A _12699_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17208_ _17207_/X _09474_/B _17414_/S vssd1 vssd1 vccd1 vccd1 _17208_/X sky130_fd_sc_hd__mux2_2
XFILLER_191_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18188_ _18216_/CLK _18188_/D vssd1 vssd1 vccd1 vccd1 _18188_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17694__S _17696_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17139_ _16542_/Y _18974_/Q _17493_/S vssd1 vssd1 vccd1 vccd1 _17139_/X sky130_fd_sc_hd__mux2_1
XANTENNA__19541__RESET_B repeater221/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14315__B1 _14314_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09961_ _19964_/Q _09960_/Y _09950_/X _09873_/B vssd1 vssd1 vccd1 vccd1 _19964_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_143_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20081_ _20081_/CLK _20081_/D repeater204/X vssd1 vssd1 vccd1 vccd1 _20081_/Q sky130_fd_sc_hd__dfrtp_1
X_09892_ _19338_/Q vssd1 vssd1 vccd1 vccd1 _09892_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18494__RESET_B repeater203/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11771__A _11771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16773__S _17385_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09326_ _20043_/Q _15721_/A vssd1 vssd1 vccd1 vccd1 _09326_/Y sky130_fd_sc_hd__nand2_1
XFILLER_166_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09257_ _10819_/A vssd1 vssd1 vccd1 vccd1 _12370_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_239_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19629__RESET_B repeater257/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14554__B1 _14513_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09188_ _20072_/Q _20071_/Q _10133_/A _08980_/Y _20073_/Q vssd1 vssd1 vccd1 vccd1
+ _09188_/X sky130_fd_sc_hd__a41o_1
XFILLER_193_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12107__A hold277/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14306__B1 _14273_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11150_ _11150_/A _11150_/B _11150_/C _17756_/X vssd1 vssd1 vccd1 vccd1 _11150_/X
+ sky130_fd_sc_hd__or4b_4
XFILLER_161_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10101_ _10101_/A _10101_/B _10101_/C vssd1 vssd1 vccd1 vccd1 _10104_/A sky130_fd_sc_hd__or3_4
XANTENNA__17109__S _17543_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11081_ _19060_/Q vssd1 vssd1 vccd1 vccd1 _11086_/A sky130_fd_sc_hd__inv_2
XFILLER_68_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10032_ _10032_/A _10032_/B _10032_/C vssd1 vssd1 vccd1 vccd1 _19936_/D sky130_fd_sc_hd__nor3_1
XFILLER_48_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_209_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16948__S _16950_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_248_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_236_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14840_ _18148_/Q _14833_/A _14814_/X _14834_/A vssd1 vssd1 vccd1 vccd1 _18148_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_75_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14085__A2 _14004_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_60_HCLK clkbuf_4_12_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20006_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_input17_A HADDR[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14771_ _14772_/A vssd1 vssd1 vccd1 vccd1 _14771_/X sky130_fd_sc_hd__clkbuf_2
X_11983_ _19370_/Q _11977_/X _11918_/X _11979_/X vssd1 vssd1 vccd1 vccd1 _19370_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_63_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16510_ _17211_/X _15904_/X _17307_/X _16509_/X vssd1 vssd1 vccd1 vccd1 _16510_/X
+ sky130_fd_sc_hd__o22a_1
X_13722_ _18757_/Q _13721_/Y _13715_/Y _13499_/X vssd1 vssd1 vccd1 vccd1 _18757_/D
+ sky130_fd_sc_hd__o22a_1
X_10934_ _15224_/A vssd1 vssd1 vccd1 vccd1 _15213_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_205_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17490_ _17489_/X _14090_/Y _17490_/S vssd1 vssd1 vccd1 vccd1 _17490_/X sky130_fd_sc_hd__mux2_2
XFILLER_17_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16441_ _19708_/Q vssd1 vssd1 vccd1 vccd1 _16441_/Y sky130_fd_sc_hd__inv_2
X_13653_ _18788_/Q _13644_/A _16951_/X _13646_/A vssd1 vssd1 vccd1 vccd1 _18788_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_32_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10865_ hold264/X vssd1 vssd1 vccd1 vccd1 _13678_/A sky130_fd_sc_hd__buf_2
XFILLER_31_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_220_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12604_ _19029_/Q _12598_/X _12533_/X _12600_/X vssd1 vssd1 vccd1 vccd1 _19029_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16372_ _19707_/Q vssd1 vssd1 vccd1 vccd1 _16372_/Y sky130_fd_sc_hd__inv_2
X_19160_ _19968_/CLK _19160_/D hold370/X vssd1 vssd1 vccd1 vccd1 _19160_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13584_ _18821_/Q _13583_/Y _13574_/X _13545_/B vssd1 vssd1 vccd1 vccd1 _18821_/D
+ sky130_fd_sc_hd__o211a_1
X_10796_ _10807_/A _10801_/A _19735_/Q vssd1 vssd1 vccd1 vccd1 _10797_/A sky130_fd_sc_hd__or3b_4
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15323_ _15323_/A vssd1 vssd1 vccd1 vccd1 _15323_/Y sky130_fd_sc_hd__inv_2
X_18111_ _18137_/CLK _18111_/D vssd1 vssd1 vccd1 vccd1 _18111_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12535_ hold332/X vssd1 vssd1 vccd1 vccd1 hold331/A sky130_fd_sc_hd__clkbuf_2
X_19091_ _19609_/CLK _19091_/D hold343/X vssd1 vssd1 vccd1 vccd1 _19091_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_12_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_repeater156_A _17523_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15254_ _19779_/Q vssd1 vssd1 vccd1 vccd1 _15254_/Y sky130_fd_sc_hd__inv_2
XFILLER_157_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18042_ _18954_/CLK _18042_/D vssd1 vssd1 vccd1 vccd1 _18042_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12466_ _19109_/Q _12464_/X _12413_/X _12465_/X vssd1 vssd1 vccd1 vccd1 _19109_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_173_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14205_ _19110_/Q vssd1 vssd1 vccd1 vccd1 _16583_/A sky130_fd_sc_hd__inv_2
XFILLER_172_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11417_ _11622_/A _19132_/Q _11579_/A _19146_/Q _11416_/X vssd1 vssd1 vccd1 vccd1
+ _11417_/X sky130_fd_sc_hd__a221o_1
X_15185_ _17934_/Q _14250_/X _10448_/A _14252_/X vssd1 vssd1 vccd1 vccd1 _17934_/D
+ sky130_fd_sc_hd__a22o_1
X_12397_ _19149_/Q _12388_/X _12396_/X _12390_/X vssd1 vssd1 vccd1 vccd1 _19149_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12017__A _12017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output85_A _16568_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14136_ _14136_/A vssd1 vssd1 vccd1 vccd1 _14136_/Y sky130_fd_sc_hd__clkinv_1
XFILLER_99_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11348_ _18976_/Q vssd1 vssd1 vccd1 vccd1 _11348_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19993_ _20003_/CLK _19993_/D repeater192/X vssd1 vssd1 vccd1 vccd1 _19993_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_235_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17019__S _17534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14067_ _14065_/Y _18682_/Q _19065_/Q _14007_/A _14066_/X vssd1 vssd1 vccd1 vccd1
+ _14067_/X sky130_fd_sc_hd__a221o_1
X_18944_ _18947_/CLK _18944_/D repeater211/X vssd1 vssd1 vccd1 vccd1 _18944_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_141_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11279_ _11482_/A _19016_/Q _11484_/A _19018_/Q _11278_/X vssd1 vssd1 vccd1 vccd1
+ _11298_/A sky130_fd_sc_hd__o221a_1
XFILLER_95_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13018_ _18924_/Q _13017_/Y _13004_/B _12958_/X vssd1 vssd1 vccd1 vccd1 _18924_/D
+ sky130_fd_sc_hd__o211a_1
X_18875_ _20048_/CLK _18875_/D repeater210/X vssd1 vssd1 vccd1 vccd1 _18875_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__16858__S _17529_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17826_ _18191_/Q _18183_/Q _18175_/Q _18159_/Q _17918_/S0 _18750_/Q vssd1 vssd1
+ vccd1 vccd1 _17826_/X sky130_fd_sc_hd__mux4_2
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17893__S0 _17913_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_239_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12087__A1 _19319_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17757_ _18520_/Q _15271_/X _18546_/Q vssd1 vssd1 vccd1 vccd1 _17757_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14969_ _18071_/Q _14964_/X _14808_/X _14966_/X vssd1 vssd1 vccd1 vccd1 _18071_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_207_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16708_ _19429_/Q vssd1 vssd1 vccd1 vccd1 _16708_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17688_ _15479_/Y _19447_/Q _17696_/S vssd1 vssd1 vccd1 vccd1 _18564_/D sky130_fd_sc_hd__mux2_1
XFILLER_35_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09061__A _12028_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19427_ _19997_/CLK _19427_/D repeater271/X vssd1 vssd1 vccd1 vccd1 _19427_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17689__S _17696_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16639_ _16912_/X _16637_/X _16916_/X _16638_/X vssd1 vssd1 vccd1 vccd1 _16639_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__16773__A1 _13399_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19358_ _19970_/CLK _19358_/D hold370/X vssd1 vssd1 vccd1 vccd1 _19358_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__19793__RESET_B repeater219/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09111_ _20089_/Q vssd1 vssd1 vccd1 vccd1 _09113_/A sky130_fd_sc_hd__inv_2
X_18309_ _18416_/CLK _18309_/D vssd1 vssd1 vccd1 vccd1 _18309_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19289_ _19290_/CLK _19289_/D repeater211/X vssd1 vssd1 vccd1 vccd1 _19289_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__19722__RESET_B repeater219/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09042_ hold315/X vssd1 vssd1 vccd1 vccd1 hold314/A sky130_fd_sc_hd__buf_4
XFILLER_136_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09944_ _19355_/Q vssd1 vssd1 vccd1 vccd1 _16671_/A sky130_fd_sc_hd__inv_2
XFILLER_89_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20064_ _20064_/CLK _20064_/D repeater200/X vssd1 vssd1 vccd1 vccd1 _20064_/Q sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_83_HCLK clkbuf_4_13_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19315_/CLK sky130_fd_sc_hd__clkbuf_16
X_09875_ _09875_/A _09875_/B vssd1 vssd1 vccd1 vccd1 _09954_/A sky130_fd_sc_hd__or2_1
XFILLER_131_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16768__S _17386_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18675__RESET_B repeater252/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17884__S0 _19633_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater250 hold367/A vssd1 vssd1 vccd1 vccd1 hold370/A sky130_fd_sc_hd__buf_8
XFILLER_234_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater261 repeater262/X vssd1 vssd1 vccd1 vccd1 repeater261/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__16461__B1 _17311_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater272 repeater273/X vssd1 vssd1 vccd1 vccd1 repeater272/X sky130_fd_sc_hd__buf_8
Xrepeater283 hold355/A vssd1 vssd1 vccd1 vccd1 hold273/A sky130_fd_sc_hd__buf_8
XPHY_4415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16069__A _16634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10089__B1 _10026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_hold249_A HWDATA[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17599__S _17600_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16764__A1 _13391_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10650_ _19790_/Q _10650_/B vssd1 vssd1 vccd1 vccd1 _10651_/B sky130_fd_sc_hd__or2_1
XANTENNA__14775__B1 _14749_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09309_ _18659_/Q _09303_/B _09304_/A vssd1 vssd1 vccd1 vccd1 _15726_/A sky130_fd_sc_hd__o21ai_1
XFILLER_22_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12250__A1 hold242/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10581_ _10581_/A _19805_/Q _10581_/C vssd1 vssd1 vccd1 vccd1 _10584_/C sky130_fd_sc_hd__or3_4
XFILLER_10_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12320_ _12362_/A vssd1 vssd1 vccd1 vccd1 _12335_/A sky130_fd_sc_hd__buf_2
XANTENNA__14527__B1 hold334/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_214_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12251_ _10954_/B _12245_/Y _15223_/A _12250_/Y vssd1 vssd1 vccd1 vccd1 _12252_/S
+ sky130_fd_sc_hd__o211ai_2
XFILLER_119_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11202_ _19578_/Q vssd1 vssd1 vccd1 vccd1 _11459_/A sky130_fd_sc_hd__inv_2
XFILLER_5_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12182_ _12180_/X _19261_/Q _12182_/S vssd1 vssd1 vccd1 vccd1 _19261_/D sky130_fd_sc_hd__mux2_1
XANTENNA__20025__CLK _20091_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11133_ _12253_/B vssd1 vssd1 vccd1 vccd1 _11133_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_3_2_0_HCLK clkbuf_3_3_0_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_5_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__18072__CLK _18169_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16990_ _16474_/Y _15608_/Y _17474_/S vssd1 vssd1 vccd1 vccd1 _16990_/X sky130_fd_sc_hd__mux2_2
X_11064_ _11064_/A _11064_/B vssd1 vssd1 vccd1 vccd1 _11066_/B sky130_fd_sc_hd__nor2_4
X_15941_ _18091_/Q vssd1 vssd1 vccd1 vccd1 _15941_/Y sky130_fd_sc_hd__inv_2
XFILLER_135_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10015_ _10087_/A _10086_/A _10015_/C _10088_/A vssd1 vssd1 vccd1 vccd1 _10016_/D
+ sky130_fd_sc_hd__or4_4
XFILLER_49_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_236_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18660_ _20048_/CLK _18660_/D repeater210/X vssd1 vssd1 vccd1 vccd1 _18660_/Q sky130_fd_sc_hd__dfrtp_1
X_15872_ _19971_/Q vssd1 vssd1 vccd1 vccd1 _15872_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17875__S0 _17908_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17611_ _15233_/Y _11861_/B _17614_/S vssd1 vssd1 vccd1 vccd1 _17611_/X sky130_fd_sc_hd__mux2_1
X_14823_ _18161_/Q _14820_/X _14745_/X _14822_/X vssd1 vssd1 vccd1 vccd1 _18161_/D
+ sky130_fd_sc_hd__a22o_1
X_18591_ _19437_/CLK _18591_/D repeater269/X vssd1 vssd1 vccd1 vccd1 _18591_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_63_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output123_A _15767_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17542_ _17541_/X _13060_/A _17542_/S vssd1 vssd1 vccd1 vccd1 _17542_/X sky130_fd_sc_hd__mux2_1
X_11966_ _19380_/Q _11962_/X _09061_/X _11963_/X vssd1 vssd1 vccd1 vccd1 _19380_/D
+ sky130_fd_sc_hd__a22o_1
X_14754_ _18197_/Q _14744_/X _14725_/X _14747_/X vssd1 vssd1 vccd1 vccd1 _18197_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_232_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10917_ _10923_/A vssd1 vssd1 vccd1 vccd1 _10924_/A sky130_fd_sc_hd__inv_2
XFILLER_189_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13705_ _18760_/Q _13710_/B vssd1 vssd1 vccd1 vccd1 _13706_/B sky130_fd_sc_hd__nand2_1
X_17473_ _17473_/A0 _15966_/Y _17473_/S vssd1 vssd1 vccd1 vccd1 _17473_/X sky130_fd_sc_hd__mux2_1
X_14685_ _18233_/Q _14682_/X _14600_/X _14684_/X vssd1 vssd1 vccd1 vccd1 _18233_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_205_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_repeater273_A repeater274/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11897_ _11897_/A1 _11891_/X _09051_/X _11892_/X vssd1 vssd1 vccd1 vccd1 _19418_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_177_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19212_ _19214_/CLK _19212_/D hold367/X vssd1 vssd1 vccd1 vccd1 _19212_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17302__S _17522_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13636_ _10195_/C _13635_/X _13632_/Y vssd1 vssd1 vccd1 vccd1 _18798_/D sky130_fd_sc_hd__a21oi_1
X_16424_ _18225_/Q vssd1 vssd1 vccd1 vccd1 _16424_/Y sky130_fd_sc_hd__inv_2
X_10848_ _19714_/Q _10843_/X _10451_/X _10845_/X vssd1 vssd1 vccd1 vccd1 _19714_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_220_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19143_ _19597_/CLK _19143_/D repeater281/X vssd1 vssd1 vccd1 vccd1 _19143_/Q sky130_fd_sc_hd__dfrtp_2
X_13567_ _18831_/Q _13566_/Y _13560_/X _13555_/B vssd1 vssd1 vccd1 vccd1 _18831_/D
+ sky130_fd_sc_hd__o211a_1
X_16355_ _18136_/Q vssd1 vssd1 vccd1 vccd1 _16355_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10779_ _17628_/X _10772_/X _19745_/Q _10774_/X vssd1 vssd1 vccd1 vccd1 _19745_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_12_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15306_ _15304_/Y _15305_/X _15287_/C _15289_/A vssd1 vssd1 vccd1 vccd1 _15306_/X
+ sky130_fd_sc_hd__a31o_1
X_12518_ _19073_/Q _12512_/X hold270/X _12513_/X vssd1 vssd1 vccd1 vccd1 _19073_/D
+ sky130_fd_sc_hd__a22o_1
X_19074_ _19610_/CLK _19074_/D hold343/X vssd1 vssd1 vccd1 vccd1 _19074_/Q sky130_fd_sc_hd__dfrtp_4
X_16286_ _17982_/Q vssd1 vssd1 vccd1 vccd1 _16286_/Y sky130_fd_sc_hd__inv_2
XFILLER_172_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13498_ _15195_/A _13618_/B vssd1 vssd1 vccd1 vccd1 _13620_/A sky130_fd_sc_hd__nand2_2
XFILLER_157_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18025_ _18145_/CLK _18025_/D vssd1 vssd1 vccd1 vccd1 _18025_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_246_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15237_ _15388_/B vssd1 vssd1 vccd1 vccd1 _15237_/Y sky130_fd_sc_hd__inv_2
X_12449_ _19120_/Q _12441_/X _12386_/X _12444_/X vssd1 vssd1 vccd1 vccd1 _19120_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_114_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15168_ _17945_/Q _15159_/A _20074_/Q _15160_/A vssd1 vssd1 vccd1 vccd1 _17945_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_99_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14119_ _14022_/A _14119_/A2 _14115_/Y _14118_/X vssd1 vssd1 vccd1 vccd1 _18692_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_125_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15099_ _17992_/Q _15095_/X _14806_/A _15097_/X vssd1 vssd1 vccd1 vccd1 _17992_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_99_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19976_ _19976_/CLK _19976_/D repeater244/X vssd1 vssd1 vccd1 vccd1 _19976_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_140_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18927_ _19325_/CLK _18927_/D repeater213/X vssd1 vssd1 vccd1 vccd1 _18927_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_140_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09660_ _09743_/A _09742_/A _09660_/C _09660_/D vssd1 vssd1 vccd1 vccd1 _09666_/B
+ sky130_fd_sc_hd__or4_4
X_18858_ _18866_/CLK _18858_/D repeater231/X vssd1 vssd1 vccd1 vccd1 _18858_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17866__S0 _17908_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_216_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17809_ _17805_/X _17806_/X _17807_/X _17808_/X _18751_/Q _18752_/Q vssd1 vssd1 vccd1
+ vccd1 _17809_/X sky130_fd_sc_hd__mux4_2
X_09591_ _09482_/A _09482_/B _09589_/Y _09587_/X vssd1 vssd1 vccd1 vccd1 _20022_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_27_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18789_ _19647_/CLK _18789_/D repeater260/X vssd1 vssd1 vccd1 vccd1 _18789_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_224_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19974__RESET_B repeater244/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16617__A _16617_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19903__RESET_B repeater195/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17212__S _17522_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14757__B1 _14693_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09025_ hold279/X vssd1 vssd1 vccd1 vccd1 _09025_/X sky130_fd_sc_hd__buf_4
XFILLER_156_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold230 hold230/A vssd1 vssd1 vccd1 vccd1 hold230/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold241 HWDATA[11] vssd1 vssd1 vccd1 vccd1 input40/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09400__A2 _19390_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold252 HWDATA[10] vssd1 vssd1 vccd1 vccd1 input39/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11743__B1 _16929_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18856__RESET_B repeater231/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold263 hold263/A vssd1 vssd1 vccd1 vccd1 hold263/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 input77/X vssd1 vssd1 vccd1 vccd1 hold274/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold285 HWDATA[31] vssd1 vssd1 vccd1 vccd1 input62/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold296 input53/X vssd1 vssd1 vccd1 vccd1 hold296/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20116_ _20120_/CLK _20116_/D repeater238/X vssd1 vssd1 vccd1 vccd1 _20116_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_131_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09927_ _19949_/Q _09924_/Y _09852_/A _19335_/Q _09926_/X vssd1 vssd1 vccd1 vccd1
+ _09928_/D sky130_fd_sc_hd__o221a_1
XFILLER_219_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09858_ _09858_/A _09858_/B vssd1 vssd1 vccd1 vccd1 _09859_/B sky130_fd_sc_hd__or2_2
XANTENNA__17857__S0 _17908_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20047_ _20048_/CLK _20047_/D repeater208/X vssd1 vssd1 vccd1 vccd1 _20047_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_85_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13248__B1 _12536_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09789_ _09789_/A _09803_/A vssd1 vssd1 vccd1 vccd1 _09790_/B sky130_fd_sc_hd__or2_2
XPHY_4201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11820_ _19446_/Q _11814_/X _10877_/X _11815_/X vssd1 vssd1 vccd1 vccd1 _19446_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11751_ _11772_/A vssd1 vssd1 vccd1 vccd1 _11751_/X sky130_fd_sc_hd__clkbuf_2
XPHY_4278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19644__RESET_B repeater261/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10702_ hold264/X vssd1 vssd1 vccd1 vccd1 _10702_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17122__S _17544_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14470_ _18357_/Q _14463_/X _14417_/X _14465_/X vssd1 vssd1 vccd1 vccd1 _18357_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14748__B1 _14745_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11682_ _19535_/Q _11668_/X _11649_/A _11669_/X vssd1 vssd1 vccd1 vccd1 _19535_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_202_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13421_ _13443_/A vssd1 vssd1 vccd1 vccd1 _13421_/X sky130_fd_sc_hd__clkbuf_2
XPHY_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10633_ _10633_/A vssd1 vssd1 vccd1 vccd1 _19802_/D sky130_fd_sc_hd__inv_2
XPHY_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16961__S _17535_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16140_ _16132_/Y _16049_/X _16133_/Y _15836_/X _16139_/X vssd1 vssd1 vccd1 vccd1
+ _16140_/X sky130_fd_sc_hd__o221a_2
XFILLER_139_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13352_ _18865_/Q _18864_/Q _13352_/C vssd1 vssd1 vccd1 vccd1 _13435_/A sky130_fd_sc_hd__and3_1
X_10564_ _15297_/A _17607_/X vssd1 vssd1 vccd1 vccd1 _10613_/C sky130_fd_sc_hd__or2b_1
XFILLER_154_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17162__A1 _19380_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11982__B1 _11981_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12303_ _19198_/Q _12298_/X _12302_/X _12300_/X vssd1 vssd1 vccd1 vccd1 _19198_/D
+ sky130_fd_sc_hd__a22o_1
X_16071_ _17472_/X _15901_/A _17440_/X _15908_/A vssd1 vssd1 vccd1 vccd1 _16071_/X
+ sky130_fd_sc_hd__o22a_2
XANTENNA__15173__B1 hold247/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13283_ _20070_/Q _13283_/B _13283_/C vssd1 vssd1 vccd1 vccd1 _13284_/A sky130_fd_sc_hd__and3_1
X_10495_ _10514_/C _10511_/A _10501_/C _11654_/B vssd1 vssd1 vccd1 vccd1 _10732_/C
+ sky130_fd_sc_hd__or4_4
XFILLER_155_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15022_ _15094_/A _15094_/B _15034_/C vssd1 vssd1 vccd1 vccd1 _15024_/A sky130_fd_sc_hd__or3_4
X_12234_ _12234_/A vssd1 vssd1 vccd1 vccd1 _12234_/X sky130_fd_sc_hd__buf_4
XFILLER_154_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18597__RESET_B repeater267/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19830_ _19846_/CLK _19830_/D repeater270/X vssd1 vssd1 vccd1 vccd1 _19830_/Q sky130_fd_sc_hd__dfrtp_4
X_12165_ _12172_/A vssd1 vssd1 vccd1 vccd1 _12165_/X sky130_fd_sc_hd__buf_1
XFILLER_122_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11116_ _11116_/A _11116_/B vssd1 vssd1 vccd1 vccd1 _11116_/Y sky130_fd_sc_hd__nor2_1
X_19761_ _19822_/CLK _19761_/D repeater228/X vssd1 vssd1 vccd1 vccd1 _19761_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_110_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16973_ _16972_/X _13414_/Y _17535_/S vssd1 vssd1 vccd1 vccd1 _16973_/X sky130_fd_sc_hd__mux2_1
X_12096_ _12096_/A vssd1 vssd1 vccd1 vccd1 _12096_/X sky130_fd_sc_hd__buf_1
X_18712_ _18718_/CLK _18712_/D repeater253/X vssd1 vssd1 vccd1 vccd1 _18712_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17848__S0 _17908_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11047_ _17753_/X vssd1 vssd1 vccd1 vccd1 _11056_/A sky130_fd_sc_hd__inv_2
X_15924_ _18067_/Q vssd1 vssd1 vccd1 vccd1 _15924_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19692_ _19720_/CLK _19692_/D repeater201/X vssd1 vssd1 vccd1 vccd1 _19692_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_65_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput9 input9/A vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__19983__CLK _19992_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18643_ _20050_/CLK _18643_/D repeater197/X vssd1 vssd1 vccd1 vccd1 _18643_/Q sky130_fd_sc_hd__dfrtp_4
X_15855_ _19815_/Q vssd1 vssd1 vccd1 vccd1 _15855_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14806_ _14806_/A vssd1 vssd1 vccd1 vccd1 _14806_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__12030__A _12030_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18574_ _19462_/CLK _18574_/D repeater272/X vssd1 vssd1 vccd1 vccd1 _18574_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__14987__B1 hold263/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15786_ _17986_/Q vssd1 vssd1 vccd1 vccd1 _15786_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_224_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12998_ _18932_/Q _12997_/Y _12980_/A _12875_/B vssd1 vssd1 vccd1 vccd1 _18932_/D
+ sky130_fd_sc_hd__o211a_1
X_17525_ _15873_/Y _10101_/B _17537_/S vssd1 vssd1 vccd1 vccd1 _17525_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12462__A1 _19111_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14737_ _18207_/Q _14732_/X _14606_/X _14734_/X vssd1 vssd1 vccd1 vccd1 _18207_/D
+ sky130_fd_sc_hd__a22o_1
X_11949_ _11956_/A vssd1 vssd1 vccd1 vccd1 _11949_/X sky130_fd_sc_hd__buf_1
XANTENNA__17032__S _17474_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17456_ _17455_/X _14053_/Y _17544_/S vssd1 vssd1 vccd1 vccd1 _17456_/X sky130_fd_sc_hd__mux2_1
XFILLER_220_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14668_ _15121_/A _14668_/B _15157_/C vssd1 vssd1 vccd1 vccd1 _14670_/A sky130_fd_sc_hd__or3_4
XFILLER_33_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_103_HCLK_A clkbuf_4_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16407_ _18017_/Q vssd1 vssd1 vccd1 vccd1 _16407_/Y sky130_fd_sc_hd__inv_2
X_13619_ _18757_/Q _15193_/A vssd1 vssd1 vccd1 vccd1 _13620_/B sky130_fd_sc_hd__or2_1
XFILLER_220_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16871__S _17535_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17387_ _16210_/Y _19266_/Q _17487_/S vssd1 vssd1 vccd1 vccd1 _17387_/X sky130_fd_sc_hd__mux2_1
X_14599_ _14601_/A vssd1 vssd1 vccd1 vccd1 _14599_/X sky130_fd_sc_hd__clkbuf_2
X_19126_ _19561_/CLK _19126_/D hold348/A vssd1 vssd1 vccd1 vccd1 _19126_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__19363__CLK _19984_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16338_ _18152_/Q vssd1 vssd1 vccd1 vccd1 _16338_/Y sky130_fd_sc_hd__inv_2
XANTENNA__09091__B1 _09090_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17153__A1 _19415_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11973__B1 _11909_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19057_ _19630_/CLK _19057_/D repeater257/X vssd1 vssd1 vccd1 vccd1 _19057_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_146_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16269_ _19637_/Q _16024_/Y _19636_/Q _15936_/Y _16268_/X vssd1 vssd1 vccd1 vccd1
+ _16269_/X sky130_fd_sc_hd__o221a_1
X_18008_ _18416_/CLK _18008_/D vssd1 vssd1 vccd1 vccd1 _18008_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13714__B2 _17908_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19959_ _19965_/CLK _19959_/D hold373/X vssd1 vssd1 vccd1 vccd1 _19959_/Q sky130_fd_sc_hd__dfrtp_4
X_09712_ _09635_/A _19404_/Q _09807_/C _19402_/Q _09711_/X vssd1 vssd1 vccd1 vccd1
+ _09713_/D sky130_fd_sc_hd__o221a_1
XANTENNA__17207__S _17413_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17839__S0 _18760_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09643_ _19980_/Q vssd1 vssd1 vccd1 vccd1 _09792_/A sky130_fd_sc_hd__inv_2
XFILLER_27_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09574_ _09574_/A vssd1 vssd1 vccd1 vccd1 _09574_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_231_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_113_HCLK clkbuf_opt_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _18623_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_224_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17392__A1 _19130_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16781__S _17414_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_25_HCLK_A clkbuf_4_9_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11964__B1 hold276/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_88_HCLK_A clkbuf_4_12_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09008_ _19506_/Q _19505_/Q vssd1 vssd1 vccd1 vccd1 _09010_/C sky130_fd_sc_hd__or2_1
XFILLER_164_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10280_ _19646_/Q _10279_/Y _19646_/Q _10279_/Y vssd1 vssd1 vccd1 vccd1 _11150_/C
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__10842__B _14245_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18690__RESET_B hold359/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16655__B1 _16914_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17117__S _17541_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13970_ _13970_/A _13970_/B _13970_/C vssd1 vssd1 vccd1 vccd1 _18705_/D sky130_fd_sc_hd__nor3_1
XFILLER_247_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12141__B1 _12078_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12921_ _12919_/Y _18928_/Q _19271_/Q _13007_/A _12920_/X vssd1 vssd1 vccd1 vccd1
+ _12924_/C sky130_fd_sc_hd__o221a_1
XFILLER_100_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17080__A0 _17486_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15640_ _18604_/Q _15640_/B vssd1 vssd1 vccd1 vccd1 _15649_/C sky130_fd_sc_hd__or2_2
XANTENNA__14969__B1 _14808_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12852_ _18932_/Q vssd1 vssd1 vccd1 vccd1 _12964_/D sky130_fd_sc_hd__inv_2
XPHY_4031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11803_ _19459_/Q _11800_/X hold300/X _11801_/X vssd1 vssd1 vccd1 vccd1 _19459_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_221_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12783_ _12764_/X _12783_/B _12783_/C _12783_/D vssd1 vssd1 vccd1 vccd1 _12834_/B
+ sky130_fd_sc_hd__and4b_1
X_15571_ _15571_/A _15571_/B vssd1 vssd1 vccd1 vccd1 _15571_/Y sky130_fd_sc_hd__nor2_1
XFILLER_92_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12785__A _18821_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10455__B1 _10421_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17310_ _16436_/Y _09222_/Y _19498_/Q vssd1 vssd1 vccd1 vccd1 _17310_/X sky130_fd_sc_hd__mux2_1
XFILLER_203_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11734_ _19503_/Q _11730_/X _16935_/X _11731_/X vssd1 vssd1 vccd1 vccd1 hold232/A
+ sky130_fd_sc_hd__a22o_1
X_14522_ _18328_/Q _14518_/X _14441_/X _14520_/X vssd1 vssd1 vccd1 vccd1 _18328_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_92_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_214_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18290_ _19873_/CLK _18290_/D vssd1 vssd1 vccd1 vccd1 _18290_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_186_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14197__A1 _19114_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17241_ _15768_/Y _14173_/Y _17546_/S vssd1 vssd1 vccd1 vccd1 _17241_/X sky130_fd_sc_hd__mux2_1
XPHY_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11665_ _11675_/A vssd1 vssd1 vccd1 vccd1 _11669_/A sky130_fd_sc_hd__inv_2
X_14453_ _14453_/A vssd1 vssd1 vccd1 vccd1 _14453_/X sky130_fd_sc_hd__clkbuf_2
XPHY_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10616_ _15297_/B _10616_/B _10616_/C _10616_/D vssd1 vssd1 vccd1 vccd1 _10617_/B
+ sky130_fd_sc_hd__or4_4
X_13404_ _20105_/Q _13430_/B _20105_/Q _13430_/B vssd1 vssd1 vccd1 vccd1 _13404_/X
+ sky130_fd_sc_hd__a2bb2o_1
XPHY_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17172_ _17171_/X _13539_/A _17536_/S vssd1 vssd1 vccd1 vccd1 _17172_/X sky130_fd_sc_hd__mux2_2
XANTENNA__09073__B1 _09071_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14384_ _18408_/Q _14380_/X _12717_/X _14382_/X vssd1 vssd1 vccd1 vccd1 _18408_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11596_ _19572_/Q _11591_/C _11592_/X _11594_/A vssd1 vssd1 vccd1 vccd1 _19572_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13335_ _13462_/A _13431_/A vssd1 vssd1 vccd1 vccd1 _13336_/B sky130_fd_sc_hd__or2_2
X_16123_ _19704_/Q vssd1 vssd1 vccd1 vccd1 _16123_/Y sky130_fd_sc_hd__inv_2
X_10547_ _19806_/Q _19805_/Q _10557_/C vssd1 vssd1 vccd1 vccd1 _10939_/D sky130_fd_sc_hd__or3_1
XFILLER_182_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17978__CLK _20123_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16054_ _19675_/Q vssd1 vssd1 vccd1 vccd1 _16054_/Y sky130_fd_sc_hd__inv_2
X_13266_ _13274_/B vssd1 vssd1 vccd1 vccd1 _14286_/B sky130_fd_sc_hd__clkbuf_2
X_10478_ _17702_/X _10471_/A _19817_/Q _10472_/A vssd1 vssd1 vccd1 vccd1 _19817_/D
+ sky130_fd_sc_hd__a22o_1
X_12217_ _19240_/Q _12212_/X _12030_/X _12213_/X vssd1 vssd1 vccd1 vccd1 _19240_/D
+ sky130_fd_sc_hd__a22o_1
X_15005_ _18052_/Q _14993_/A _15004_/X _14994_/A vssd1 vssd1 vccd1 vccd1 _18052_/D
+ sky130_fd_sc_hd__a22o_1
X_13197_ _18898_/Q _13199_/A _13180_/X _13197_/C1 vssd1 vssd1 vccd1 vccd1 _18898_/D
+ sky130_fd_sc_hd__o211a_1
X_19813_ _19813_/CLK _19813_/D repeater224/X vssd1 vssd1 vccd1 vccd1 _19813_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_111_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12148_ _19285_/Q _12143_/X _12090_/X _12144_/X vssd1 vssd1 vccd1 vccd1 _19285_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_243_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17027__S _17523_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19744_ _20070_/CLK _19744_/D repeater207/X vssd1 vssd1 vccd1 vccd1 _19744_/Q sky130_fd_sc_hd__dfrtp_1
X_12079_ _19322_/Q _12068_/X _12078_/X _12072_/X vssd1 vssd1 vccd1 vccd1 _19322_/D
+ sky130_fd_sc_hd__a22o_1
X_16956_ _17794_/X _18794_/Q _16957_/S vssd1 vssd1 vccd1 vccd1 _16956_/X sky130_fd_sc_hd__mux2_1
XFILLER_111_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_238_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_136_HCLK clkbuf_4_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20003_/CLK sky130_fd_sc_hd__clkbuf_16
X_15907_ _16234_/A vssd1 vssd1 vccd1 vccd1 _15908_/A sky130_fd_sc_hd__buf_1
X_19675_ _19822_/CLK _19675_/D repeater218/X vssd1 vssd1 vccd1 vccd1 _19675_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12683__A1 _18977_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16887_ _17473_/A0 _16738_/Y _17473_/S vssd1 vssd1 vccd1 vccd1 _16887_/X sky130_fd_sc_hd__mux2_1
XANTENNA__16866__S _17524_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_238_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18626_ _19814_/CLK _18626_/D repeater223/X vssd1 vssd1 vccd1 vccd1 _18626_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_92_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15838_ _15973_/A vssd1 vssd1 vccd1 vccd1 _15838_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_52_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18557_ _19992_/CLK _18557_/D repeater193/X vssd1 vssd1 vccd1 vccd1 _18557_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_17_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12435__B2 _12402_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15769_ _15769_/A vssd1 vssd1 vccd1 vccd1 _16669_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_206_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15071__A _15072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17508_ _17507_/X _17904_/X _17568_/S vssd1 vssd1 vccd1 vccd1 _17508_/X sky130_fd_sc_hd__mux2_1
X_09290_ _20047_/Q _09285_/X _09082_/X _09287_/X vssd1 vssd1 vccd1 vccd1 _20047_/D
+ sky130_fd_sc_hd__a22o_1
X_18488_ _19812_/CLK _18488_/D repeater225/X vssd1 vssd1 vccd1 vccd1 _18488_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_221_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17439_ _17473_/A0 _16048_/Y _17512_/S vssd1 vssd1 vccd1 vccd1 _17439_/X sky130_fd_sc_hd__mux2_1
XFILLER_165_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20053__RESET_B repeater205/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11946__B1 _09025_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16614__B _16614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19109_ _19109_/CLK _19109_/D hold361/X vssd1 vssd1 vccd1 vccd1 _19109_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__15137__B1 hold247/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14415__A hold325/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16885__A0 _17473_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput110 _16499_/Y vssd1 vssd1 vccd1 vccd1 HRDATA[9] sky130_fd_sc_hd__clkbuf_2
Xoutput121 _16752_/X vssd1 vssd1 vccd1 vccd1 IRQ[3] sky130_fd_sc_hd__clkbuf_2
Xoutput132 _19876_/Q vssd1 vssd1 vccd1 vccd1 SCLK_S2 sky130_fd_sc_hd__clkbuf_2
XFILLER_217_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput143 _16762_/LO vssd1 vssd1 vccd1 vccd1 sda_o_S5 sky130_fd_sc_hd__clkbuf_2
XFILLER_142_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_247_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12123__B1 _11978_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16776__S _17413_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09626_ _19998_/Q vssd1 vssd1 vccd1 vccd1 _09753_/C sky130_fd_sc_hd__inv_2
X_09557_ _20012_/Q _16471_/A _20029_/Q _09556_/Y vssd1 vssd1 vccd1 vccd1 _09557_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_43_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10437__B1 _09061_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_224_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09488_ _09488_/A _09488_/B vssd1 vssd1 vccd1 vccd1 _09577_/A sky130_fd_sc_hd__or2_1
XFILLER_23_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_hold329_A scl_i_S5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17400__S _17564_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11450_ _19153_/Q vssd1 vssd1 vccd1 vccd1 _11450_/Y sky130_fd_sc_hd__inv_2
XPHY_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_17_HCLK clkbuf_4_3_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _18460_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_127_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10401_ _14490_/A _14477_/B _10396_/Y _14990_/A _10400_/X vssd1 vssd1 vccd1 vccd1
+ _19851_/D sky130_fd_sc_hd__a32o_1
X_11381_ _19131_/Q vssd1 vssd1 vccd1 vccd1 _11381_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16876__A0 _15963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13120_ _19186_/Q _13087_/A _13119_/Y _18915_/Q vssd1 vssd1 vccd1 vccd1 _13120_/X
+ sky130_fd_sc_hd__o22a_1
X_10332_ _10332_/A _10332_/B vssd1 vssd1 vccd1 vccd1 _10335_/A sky130_fd_sc_hd__or2_1
XFILLER_164_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13051_ _18895_/Q vssd1 vssd1 vccd1 vccd1 _13068_/A sky130_fd_sc_hd__inv_2
XFILLER_127_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10263_ _19647_/Q vssd1 vssd1 vccd1 vccd1 _10263_/X sky130_fd_sc_hd__buf_1
X_12002_ _12044_/A vssd1 vssd1 vccd1 vccd1 _12017_/A sky130_fd_sc_hd__buf_2
XANTENNA__16628__B1 _17074_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_159_HCLK clkbuf_4_0_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _18441_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_78_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10194_ _18798_/Q vssd1 vssd1 vccd1 vccd1 _10195_/C sky130_fd_sc_hd__inv_2
XFILLER_239_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16810_ _15768_/Y _14167_/Y _17546_/S vssd1 vssd1 vccd1 vccd1 _16810_/X sky130_fd_sc_hd__mux2_1
X_17790_ _18319_/Q _18439_/Q _18431_/Q _18423_/Q _17923_/S0 _19646_/Q vssd1 vssd1
+ vccd1 vccd1 _17790_/X sky130_fd_sc_hd__mux4_1
X_16741_ _16884_/X _16513_/A _16886_/X _16002_/X vssd1 vssd1 vccd1 vccd1 _16741_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12665__A1 _18991_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13953_ _13951_/A _13951_/B _13951_/Y _13919_/X vssd1 vssd1 vccd1 vccd1 _18714_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_235_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19460_ _19462_/CLK _19460_/D repeater272/X vssd1 vssd1 vccd1 vccd1 _19460_/Q sky130_fd_sc_hd__dfrtp_4
X_12904_ _12901_/Y _18919_/Q _19262_/Q _12864_/A _12903_/X vssd1 vssd1 vccd1 vccd1
+ _12908_/C sky130_fd_sc_hd__o221a_1
XFILLER_235_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16672_ _19463_/Q _16673_/B vssd1 vssd1 vccd1 vccd1 _16672_/Y sky130_fd_sc_hd__nand2_1
XFILLER_47_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13884_ _19204_/Q _18715_/Q _13883_/Y _13812_/C vssd1 vssd1 vccd1 vccd1 _13884_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08993__A _19515_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_234_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14406__A2 _14395_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18411_ _18412_/CLK _18411_/D vssd1 vssd1 vccd1 vccd1 _18411_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_234_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15623_ _15621_/Y _15622_/Y _15614_/X vssd1 vssd1 vccd1 vccd1 _15623_/X sky130_fd_sc_hd__o21a_1
X_12835_ _13588_/A vssd1 vssd1 vccd1 vccd1 _13597_/A sky130_fd_sc_hd__clkbuf_4
X_19391_ _19933_/CLK _19391_/D repeater236/X vssd1 vssd1 vccd1 vccd1 _19391_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_62_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_repeater186_A repeater188/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10428__B1 _10427_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18342_ _18473_/CLK _18342_/D vssd1 vssd1 vccd1 vccd1 _18342_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_188_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15554_ _18582_/Q vssd1 vssd1 vccd1 vccd1 _15557_/A sky130_fd_sc_hd__inv_2
X_12766_ _18834_/Q vssd1 vssd1 vccd1 vccd1 _13557_/A sky130_fd_sc_hd__inv_2
XPHY_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14505_ _14505_/A vssd1 vssd1 vccd1 vccd1 _14505_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__18959__RESET_B repeater257/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11717_ _11731_/A vssd1 vssd1 vccd1 vccd1 _11717_/X sky130_fd_sc_hd__clkbuf_2
X_18273_ _20081_/CLK _18273_/D vssd1 vssd1 vccd1 vccd1 _18273_/Q sky130_fd_sc_hd__dfxtp_1
X_12697_ _18967_/Q _12691_/X _12596_/X _12692_/X vssd1 vssd1 vccd1 vccd1 _18967_/D
+ sky130_fd_sc_hd__a22o_1
X_15485_ _18566_/Q vssd1 vssd1 vccd1 vccd1 _15487_/A sky130_fd_sc_hd__inv_2
XANTENNA__15906__A2 _15896_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17310__S _19498_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17224_ _17223_/X _14035_/Y _17544_/S vssd1 vssd1 vccd1 vccd1 _17224_/X sky130_fd_sc_hd__mux2_1
XPHY_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11648_ _11648_/A vssd1 vssd1 vccd1 vccd1 _15311_/A sky130_fd_sc_hd__buf_2
XANTENNA__09046__B1 hold300/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14436_ _14438_/A vssd1 vssd1 vccd1 vccd1 _14436_/X sky130_fd_sc_hd__clkbuf_2
Xinput12 input12/A vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__buf_1
XFILLER_11_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput23 input23/A vssd1 vssd1 vccd1 vccd1 input23/X sky130_fd_sc_hd__buf_1
XPHY_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput34 HRESETn vssd1 vssd1 vccd1 vccd1 input34/X sky130_fd_sc_hd__buf_6
XPHY_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput45 input45/A vssd1 vssd1 vccd1 vccd1 input45/X sky130_fd_sc_hd__clkbuf_4
XFILLER_7_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17155_ _16484_/X _08930_/Y _17566_/S vssd1 vssd1 vccd1 vccd1 _17155_/X sky130_fd_sc_hd__mux2_1
X_11579_ _11579_/A _11579_/B vssd1 vssd1 vccd1 vccd1 _11603_/A sky130_fd_sc_hd__or2_1
X_14367_ _14368_/A vssd1 vssd1 vccd1 vccd1 _14367_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_156_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput56 input56/A vssd1 vssd1 vccd1 vccd1 input56/X sky130_fd_sc_hd__clkbuf_4
XFILLER_183_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16867__A0 _15768_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput67 input67/A vssd1 vssd1 vccd1 vccd1 input67/X sky130_fd_sc_hd__buf_4
Xinput78 input78/A vssd1 vssd1 vccd1 vccd1 input78/X sky130_fd_sc_hd__buf_1
XFILLER_183_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16106_ _18077_/Q vssd1 vssd1 vccd1 vccd1 _16106_/Y sky130_fd_sc_hd__inv_2
X_13318_ _18841_/Q vssd1 vssd1 vccd1 vccd1 _13464_/A sky130_fd_sc_hd__inv_4
XFILLER_6_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17086_ _17085_/X _13875_/Y _17545_/S vssd1 vssd1 vccd1 vccd1 _17086_/X sky130_fd_sc_hd__mux2_1
X_14298_ _18450_/Q _14289_/A _13682_/X _14290_/A vssd1 vssd1 vccd1 vccd1 _18450_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18156__CLK _20123_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_182_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19401__CLK _19976_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16037_ _17979_/Q vssd1 vssd1 vccd1 vccd1 _16037_/Y sky130_fd_sc_hd__inv_2
X_13249_ _18874_/Q _13242_/A _12538_/X _13243_/A vssd1 vssd1 vccd1 vccd1 _18874_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10903__A1 _19685_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19747__RESET_B repeater205/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_229_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16600__D _16600_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17988_ _19851_/CLK _17988_/D vssd1 vssd1 vccd1 vccd1 _17988_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12105__B1 _12104_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19727_ _20055_/CLK _19727_/D repeater205/X vssd1 vssd1 vccd1 vccd1 _19727_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__09064__A _12030_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16939_ _19483_/Q hold174/X _16946_/S vssd1 vssd1 vccd1 vccd1 _16939_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12656__A1 _18994_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17044__A0 _17473_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_225_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19658_ _19668_/CLK _19658_/D repeater270/X vssd1 vssd1 vccd1 vccd1 _19658_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__10131__A2 _10130_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09411_ _19368_/Q vssd1 vssd1 vccd1 vccd1 _09411_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18609_ _19566_/CLK _18609_/D repeater255/X vssd1 vssd1 vccd1 vccd1 _18609_/Q sky130_fd_sc_hd__dfrtp_1
X_19589_ _19610_/CLK _19589_/D hold343/X vssd1 vssd1 vccd1 vccd1 _19589_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_225_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09342_ _09255_/X _20036_/Q _09342_/S vssd1 vssd1 vccd1 vccd1 _20036_/D sky130_fd_sc_hd__mux2_1
XFILLER_206_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09273_ _20056_/Q _09269_/X _09086_/X _09271_/X vssd1 vssd1 vccd1 vccd1 _20056_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_221_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17220__S _17385_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16344__B _16344_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11919__B1 _11918_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_181_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12592__B1 _12353_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17283__A0 _17473_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19488__RESET_B repeater260/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_hold181_A HADDR[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08988_ _19518_/Q vssd1 vssd1 vccd1 vccd1 _10819_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_57_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19417__RESET_B repeater210/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_217_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10950_ _10950_/A vssd1 vssd1 vccd1 vccd1 _11772_/A sky130_fd_sc_hd__buf_2
XFILLER_217_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17586__A1 _19717_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09609_ _09609_/A vssd1 vssd1 vccd1 vccd1 _09609_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10881_ hold237/X vssd1 vssd1 vccd1 vccd1 _14277_/A sky130_fd_sc_hd__buf_4
XFILLER_44_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12620_ _19020_/Q _12613_/X _12384_/X _12616_/X vssd1 vssd1 vccd1 vccd1 _19020_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09276__B1 _09098_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_244_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12551_ _12551_/A _12553_/A _12551_/C vssd1 vssd1 vccd1 vccd1 _12551_/X sky130_fd_sc_hd__or3_2
XPHY_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11502_ _11482_/A _11502_/A2 _11528_/A _11500_/Y vssd1 vssd1 vccd1 vccd1 _19602_/D
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__17130__S _17490_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15270_ _15270_/A _15270_/B _15270_/C vssd1 vssd1 vccd1 vccd1 _15271_/B sky130_fd_sc_hd__or3_1
XANTENNA__09028__B1 _09027_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12482_ _19097_/Q _12478_/X _12232_/X _12479_/X vssd1 vssd1 vccd1 vccd1 _19097_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_200_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14221_ _18491_/Q _18490_/Q vssd1 vssd1 vccd1 vccd1 _14222_/B sky130_fd_sc_hd__or2_1
X_11433_ _11417_/X _11433_/B _11433_/C _11433_/D vssd1 vssd1 vccd1 vccd1 _11457_/C
+ sky130_fd_sc_hd__and4b_1
XPHY_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14152_ _19093_/Q vssd1 vssd1 vccd1 vccd1 _14152_/Y sky130_fd_sc_hd__inv_2
X_11364_ _11521_/A vssd1 vssd1 vccd1 vccd1 _11504_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_164_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13103_ _19187_/Q _13088_/A _16667_/A _18911_/Q vssd1 vssd1 vccd1 vccd1 _13103_/X
+ sky130_fd_sc_hd__o22a_1
X_10315_ _19870_/Q _10314_/X _10293_/Y vssd1 vssd1 vccd1 vccd1 _19870_/D sky130_fd_sc_hd__o21a_1
X_18960_ _19600_/CLK _18960_/D hold273/X vssd1 vssd1 vccd1 vccd1 _18960_/Q sky130_fd_sc_hd__dfrtp_4
X_14083_ _19065_/Q _14007_/A _14081_/Y _18675_/Q _14082_/X vssd1 vssd1 vccd1 vccd1
+ _14093_/A sky130_fd_sc_hd__o221a_1
XFILLER_4_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11295_ _19021_/Q vssd1 vssd1 vccd1 vccd1 _16716_/A sky130_fd_sc_hd__inv_2
XANTENNA__08988__A _19518_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17911_ _15786_/Y _15787_/Y _15788_/Y _15789_/Y _17913_/S0 _19632_/Q vssd1 vssd1
+ vccd1 vccd1 _17911_/X sky130_fd_sc_hd__mux4_2
X_13034_ _18912_/Q vssd1 vssd1 vccd1 vccd1 _13084_/A sky130_fd_sc_hd__inv_2
X_10246_ _10246_/A _10246_/B _10246_/C _10246_/D vssd1 vssd1 vccd1 vccd1 _10247_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_140_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18891_ _19964_/CLK _18891_/D hold372/X vssd1 vssd1 vccd1 vccd1 _18891_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_239_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19840__RESET_B repeater272/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10897__B1 _10882_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17842_ _16406_/Y _16407_/Y _16408_/Y _16409_/Y _17913_/S0 _19632_/Q vssd1 vssd1
+ vccd1 vccd1 _17842_/X sky130_fd_sc_hd__mux4_1
X_10177_ _19881_/Q _10174_/X _09098_/X _10175_/X vssd1 vssd1 vccd1 vccd1 _19881_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19158__RESET_B repeater212/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17773_ _18291_/Q _18283_/Q _18275_/Q _18443_/Q _17923_/S0 _19646_/Q vssd1 vssd1
+ vccd1 vccd1 _17773_/X sky130_fd_sc_hd__mux4_2
X_14985_ _18062_/Q _14976_/X _14791_/X _14979_/X vssd1 vssd1 vccd1 vccd1 _18062_/D
+ sky130_fd_sc_hd__a22o_1
X_19512_ _19513_/CLK hold225/X repeater259/X vssd1 vssd1 vccd1 vccd1 _19512_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__09503__B2 _19317_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15614__A _15643_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17305__S _17546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16724_ _16779_/X _15887_/X _16778_/X _16591_/X vssd1 vssd1 vccd1 vccd1 _16728_/A
+ sky130_fd_sc_hd__o22ai_2
XFILLER_47_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13936_ _18721_/Q _13935_/Y _13821_/B _13925_/X vssd1 vssd1 vccd1 vccd1 _18721_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_235_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19443_ _19992_/CLK _19443_/D repeater198/X vssd1 vssd1 vccd1 vccd1 _19443_/Q sky130_fd_sc_hd__dfrtp_1
X_16655_ _16909_/X _16597_/X _16914_/X _16598_/X vssd1 vssd1 vccd1 vccd1 _16656_/D
+ sky130_fd_sc_hd__a22o_2
XFILLER_235_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13867_ _13867_/A _13867_/B _13867_/C _13867_/D vssd1 vssd1 vccd1 vccd1 _13898_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_90_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13599__C1 _13560_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15606_ _15606_/A _15606_/B vssd1 vssd1 vccd1 vccd1 _15606_/Y sky130_fd_sc_hd__nor2_1
X_12818_ _18831_/Q vssd1 vssd1 vccd1 vccd1 _13554_/A sky130_fd_sc_hd__inv_2
X_19374_ _19971_/CLK _19374_/D repeater241/X vssd1 vssd1 vccd1 vccd1 _19374_/Q sky130_fd_sc_hd__dfrtp_4
X_16586_ _16586_/A _16615_/B vssd1 vssd1 vccd1 vccd1 _16586_/Y sky130_fd_sc_hd__nor2_1
XFILLER_34_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13798_ _18708_/Q vssd1 vssd1 vccd1 vccd1 _13945_/A sky130_fd_sc_hd__inv_2
XFILLER_203_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18793__RESET_B repeater261/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18325_ _19637_/CLK _18325_/D vssd1 vssd1 vccd1 vccd1 _18325_/Q sky130_fd_sc_hd__dfxtp_1
X_15537_ _15537_/A _15537_/B vssd1 vssd1 vccd1 vccd1 _15538_/A sky130_fd_sc_hd__or2_1
XFILLER_188_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12749_ _19251_/Q vssd1 vssd1 vccd1 vccd1 _16668_/A sky130_fd_sc_hd__inv_2
XFILLER_231_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17040__S _17493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18722__RESET_B repeater253/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18256_ _20081_/CLK _18256_/D vssd1 vssd1 vccd1 vccd1 _18256_/Q sky130_fd_sc_hd__dfxtp_1
X_15468_ _15471_/B _15467_/Y _15459_/X vssd1 vssd1 vccd1 vccd1 _15468_/X sky130_fd_sc_hd__o21a_1
X_17207_ _17206_/X _09407_/Y _17413_/S vssd1 vssd1 vccd1 vccd1 _17207_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14419_ _14727_/A vssd1 vssd1 vccd1 vccd1 _14419_/X sky130_fd_sc_hd__buf_2
X_18187_ _18460_/CLK _18187_/D vssd1 vssd1 vccd1 vccd1 _18187_/Q sky130_fd_sc_hd__dfxtp_1
X_15399_ _18532_/Q _13219_/B _13220_/B vssd1 vssd1 vccd1 vccd1 _15399_/X sky130_fd_sc_hd__a21bo_1
XFILLER_144_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12574__B1 _12396_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17138_ _16550_/Y _15501_/Y _17513_/S vssd1 vssd1 vccd1 vccd1 _17138_/X sky130_fd_sc_hd__mux2_1
XANTENNA__17501__A1 _08946_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19928__RESET_B repeater230/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09960_ _09960_/A vssd1 vssd1 vccd1 vccd1 _09960_/Y sky130_fd_sc_hd__inv_2
X_17069_ _16670_/Y _19390_/Q _17413_/S vssd1 vssd1 vccd1 vccd1 _17069_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12326__B1 _12080_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20080_ _20081_/CLK _20080_/D repeater204/X vssd1 vssd1 vccd1 vccd1 _20080_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_69_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09891_ _19336_/Q vssd1 vssd1 vccd1 vccd1 _09891_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16068__B2 _15915_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10888__B1 _10863_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14079__B1 _19078_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_214_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17017__A0 _17016_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17215__S _17566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17568__A1 _17914_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_225_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09325_ _15723_/A vssd1 vssd1 vccd1 vccd1 _09325_/Y sky130_fd_sc_hd__inv_2
XFILLER_159_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09256_ _11936_/A vssd1 vssd1 vccd1 vccd1 _12257_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_138_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09187_ _20124_/Q vssd1 vssd1 vccd1 vccd1 _10133_/B sky130_fd_sc_hd__buf_1
XFILLER_193_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12565__B1 _12380_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10100_ _19910_/Q _10103_/A _10097_/A _10026_/X vssd1 vssd1 vccd1 vccd1 _19910_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_161_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11080_ _19226_/Q vssd1 vssd1 vccd1 vccd1 _15222_/A sky130_fd_sc_hd__inv_2
XFILLER_248_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10031_ _10023_/C _10051_/B _10023_/A vssd1 vssd1 vccd1 vccd1 _10032_/C sky130_fd_sc_hd__o21a_1
XFILLER_0_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_1_1_0_HCLK_A clkbuf_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11962__A _11977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17125__S _17547_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14770_ _14819_/A _14975_/B _15082_/C vssd1 vssd1 vccd1 vccd1 _14772_/A sky130_fd_sc_hd__or3_4
XFILLER_91_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11982_ _19371_/Q _11977_/X _11981_/X _11979_/X vssd1 vssd1 vccd1 vccd1 _19371_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_217_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13721_ _13721_/A _13721_/B _13721_/C _13721_/D vssd1 vssd1 vccd1 vccd1 _13721_/Y
+ sky130_fd_sc_hd__nor4_2
XFILLER_232_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10933_ _10933_/A _10933_/B vssd1 vssd1 vccd1 vccd1 _10933_/X sky130_fd_sc_hd__and2_1
XANTENNA__16964__S _17482_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16440_ _19692_/Q vssd1 vssd1 vccd1 vccd1 _16440_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10864_ _19704_/Q _10855_/X _10863_/X _10857_/X vssd1 vssd1 vccd1 vccd1 _19704_/D
+ sky130_fd_sc_hd__a22o_1
X_13652_ _16952_/X _13644_/A _18789_/Q _13646_/A vssd1 vssd1 vccd1 vccd1 _18789_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_220_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12603_ _19030_/Q _12598_/X _12602_/X _12600_/X vssd1 vssd1 vccd1 vccd1 _19030_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16371_ _19691_/Q vssd1 vssd1 vccd1 vccd1 _16371_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13583_ _13583_/A vssd1 vssd1 vccd1 vccd1 _13583_/Y sky130_fd_sc_hd__inv_2
X_10795_ _19734_/Q vssd1 vssd1 vccd1 vccd1 _10801_/A sky130_fd_sc_hd__inv_2
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18110_ _18137_/CLK _18110_/D vssd1 vssd1 vccd1 vccd1 _18110_/Q sky130_fd_sc_hd__dfxtp_1
X_15322_ _15322_/A _15322_/B _15322_/C vssd1 vssd1 vccd1 vccd1 _15322_/X sky130_fd_sc_hd__and3_1
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19090_ _19609_/CLK _19090_/D hold343/X vssd1 vssd1 vccd1 vccd1 _19090_/Q sky130_fd_sc_hd__dfrtp_4
X_12534_ _19065_/Q _12528_/X _12533_/X _12529_/X vssd1 vssd1 vccd1 vccd1 _19065_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_169_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18041_ _18142_/CLK _18041_/D vssd1 vssd1 vccd1 vccd1 _18041_/Q sky130_fd_sc_hd__dfxtp_1
X_15253_ _19777_/Q vssd1 vssd1 vccd1 vccd1 _15253_/Y sky130_fd_sc_hd__inv_2
XFILLER_149_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12465_ _12479_/A vssd1 vssd1 vccd1 vccd1 _12465_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_repeater149_A _15963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14204_ _19098_/Q vssd1 vssd1 vccd1 vccd1 _14204_/Y sky130_fd_sc_hd__inv_2
X_11416_ _19565_/Q _19145_/Q _11578_/A _11415_/Y vssd1 vssd1 vccd1 vccd1 _11416_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_153_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12396_ hold296/X vssd1 vssd1 vccd1 vccd1 _12396_/X sky130_fd_sc_hd__buf_2
X_15184_ _17935_/Q _14250_/X _10446_/A _14252_/X vssd1 vssd1 vccd1 vccd1 _17935_/D
+ sky130_fd_sc_hd__a22o_1
X_11347_ _11347_/A _11347_/B _11347_/C _11347_/D vssd1 vssd1 vccd1 vccd1 _11362_/C
+ sky130_fd_sc_hd__and4_1
X_14135_ _14135_/A _14135_/B _14135_/C vssd1 vssd1 vccd1 vccd1 _18682_/D sky130_fd_sc_hd__nor3_1
X_19992_ _19992_/CLK _19992_/D repeater192/X vssd1 vssd1 vccd1 vccd1 _19992_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_153_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12308__B1 _12241_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19339__RESET_B repeater245/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11278_ _19602_/Q _16665_/A _11461_/A _18994_/Q vssd1 vssd1 vccd1 vccd1 _11278_/X
+ sky130_fd_sc_hd__o22a_1
X_14066_ _19083_/Q _14024_/A _19083_/Q _14024_/A vssd1 vssd1 vccd1 vccd1 _14066_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_113_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18943_ _18947_/CLK _18943_/D repeater213/X vssd1 vssd1 vccd1 vccd1 _18943_/Q sky130_fd_sc_hd__dfrtp_4
X_10229_ _19827_/Q _10224_/X _19829_/Q _10956_/D _10228_/X vssd1 vssd1 vccd1 vccd1
+ _10246_/A sky130_fd_sc_hd__o221a_1
X_13017_ _13017_/A vssd1 vssd1 vccd1 vccd1 _13017_/Y sky130_fd_sc_hd__inv_2
X_18874_ _20048_/CLK _18874_/D repeater208/X vssd1 vssd1 vccd1 vccd1 _18874_/Q sky130_fd_sc_hd__dfrtp_1
X_17825_ _18335_/Q _18215_/Q _18207_/Q _18199_/Q _17918_/S0 _18750_/Q vssd1 vssd1
+ vccd1 vccd1 _17825_/X sky130_fd_sc_hd__mux4_1
XFILLER_239_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17893__S1 _19632_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17035__S _17488_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17756_ _17753_/S _12058_/A _17756_/S vssd1 vssd1 vccd1 vccd1 _17756_/X sky130_fd_sc_hd__mux2_1
XFILLER_208_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14968_ _18072_/Q _14964_/X _14806_/X _14966_/X vssd1 vssd1 vccd1 vccd1 _18072_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_48_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16707_ _19394_/Q vssd1 vssd1 vccd1 vccd1 _16707_/Y sky130_fd_sc_hd__inv_4
XFILLER_207_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13919_ _13927_/A vssd1 vssd1 vccd1 vccd1 _13919_/X sky130_fd_sc_hd__buf_2
X_17687_ _15484_/X _19448_/Q _17696_/S vssd1 vssd1 vccd1 vccd1 _18565_/D sky130_fd_sc_hd__mux2_1
XANTENNA__16874__S _17541_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14899_ _18113_/Q _14896_/X _14699_/X _14898_/X vssd1 vssd1 vccd1 vccd1 _18113_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_222_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19426_ _19997_/CLK _19426_/D repeater185/X vssd1 vssd1 vccd1 vccd1 _19426_/Q sky130_fd_sc_hd__dfrtp_1
X_16638_ _16638_/A vssd1 vssd1 vccd1 vccd1 _16638_/X sky130_fd_sc_hd__buf_1
XFILLER_222_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19357_ _19968_/CLK _19357_/D hold371/X vssd1 vssd1 vccd1 vccd1 _19357_/Q sky130_fd_sc_hd__dfrtp_1
X_16569_ _19455_/Q vssd1 vssd1 vccd1 vccd1 _16569_/Y sky130_fd_sc_hd__inv_2
XFILLER_200_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09110_ _20090_/Q vssd1 vssd1 vccd1 vccd1 _09127_/A sky130_fd_sc_hd__inv_2
XFILLER_31_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18308_ _18431_/CLK _18308_/D vssd1 vssd1 vccd1 vccd1 _18308_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19288_ _19288_/CLK _19288_/D repeater211/X vssd1 vssd1 vccd1 vccd1 _19288_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__11102__A1_N _19634_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09041_ _09041_/A vssd1 vssd1 vccd1 vccd1 _09041_/X sky130_fd_sc_hd__clkbuf_2
X_18239_ _20077_/CLK _18239_/D vssd1 vssd1 vccd1 vccd1 _18239_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_176_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_175_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16622__B _16622_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17486__A0 _17486_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10951__A _11772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09943_ _19362_/Q vssd1 vssd1 vccd1 vccd1 _09943_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17238__A0 _15768_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20063_ _20064_/CLK _20063_/D repeater200/X vssd1 vssd1 vccd1 vccd1 _20063_/Q sky130_fd_sc_hd__dfrtp_1
X_09874_ _09874_/A _09957_/A vssd1 vssd1 vccd1 vccd1 _09875_/B sky130_fd_sc_hd__or2_2
XFILLER_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_246_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17884__S1 _19634_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater240 repeater241/X vssd1 vssd1 vccd1 vccd1 repeater240/X sky130_fd_sc_hd__buf_6
XFILLER_39_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrepeater251 hold366/A vssd1 vssd1 vccd1 vccd1 hold350/A sky130_fd_sc_hd__buf_8
XANTENNA__11782__A _15772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater262 repeater263/X vssd1 vssd1 vccd1 vccd1 repeater262/X sky130_fd_sc_hd__buf_8
XANTENNA__16461__B2 _15999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater273 repeater274/X vssd1 vssd1 vccd1 vccd1 repeater273/X sky130_fd_sc_hd__buf_6
XFILLER_73_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater284 hold356/A vssd1 vssd1 vccd1 vccd1 hold358/A sky130_fd_sc_hd__buf_4
XPHY_4427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_241_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16784__S _17513_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18837__CLK _18866_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_210_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09308_ _20048_/Q vssd1 vssd1 vccd1 vccd1 _09308_/Y sky130_fd_sc_hd__inv_2
X_10580_ _19806_/Q vssd1 vssd1 vccd1 vccd1 _10581_/A sky130_fd_sc_hd__inv_2
XANTENNA_hold311_A HWDATA[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09239_ _19884_/Q _15712_/A _19884_/Q _15712_/A vssd1 vssd1 vccd1 vccd1 _09239_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_167_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12250_ hold242/X _12556_/A _17612_/X vssd1 vssd1 vccd1 vccd1 _12250_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_182_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11201_ _19019_/Q vssd1 vssd1 vccd1 vccd1 _11201_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17477__A0 _17486_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12181_ _12187_/A _12309_/A vssd1 vssd1 vccd1 vccd1 _12182_/S sky130_fd_sc_hd__or2_1
XFILLER_79_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10861__A _12232_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11132_ _19629_/Q _19628_/Q vssd1 vssd1 vccd1 vccd1 _12253_/B sky130_fd_sc_hd__nand2_1
XANTENNA__16959__S _17542_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11063_ _19631_/Q vssd1 vssd1 vccd1 vccd1 _11064_/B sky130_fd_sc_hd__inv_2
X_15940_ _18123_/Q vssd1 vssd1 vccd1 vccd1 _15940_/Y sky130_fd_sc_hd__inv_2
XANTENNA__09706__B2 _19429_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10014_ _10085_/A _10084_/A _10083_/A _10101_/A vssd1 vssd1 vccd1 vccd1 _10016_/C
+ sky130_fd_sc_hd__or4_4
XFILLER_76_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15871_ _19261_/Q _15878_/B vssd1 vssd1 vccd1 vccd1 _15871_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__17875__S1 _18759_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15255__A2 _15253_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17610_ _15233_/Y _15202_/Y _17614_/S vssd1 vssd1 vccd1 vccd1 _17610_/X sky130_fd_sc_hd__mux2_1
X_14822_ _14822_/A vssd1 vssd1 vccd1 vccd1 _14822_/X sky130_fd_sc_hd__clkbuf_2
X_18590_ _19437_/CLK _18590_/D repeater269/X vssd1 vssd1 vccd1 vccd1 _18590_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_236_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17541_ _17540_/X _12901_/Y _17541_/S vssd1 vssd1 vccd1 vccd1 _17541_/X sky130_fd_sc_hd__mux2_1
X_14753_ _18198_/Q _14744_/X _14723_/X _14747_/X vssd1 vssd1 vccd1 vccd1 _18198_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_217_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11965_ _19381_/Q _11962_/X _09058_/X _11963_/X vssd1 vssd1 vccd1 vccd1 _19381_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_151_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11842__D _11842_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13704_ _13704_/A _13704_/B vssd1 vssd1 vccd1 vccd1 _13710_/B sky130_fd_sc_hd__nor2_4
X_10916_ _18511_/Q _18510_/Q vssd1 vssd1 vccd1 vccd1 _10923_/A sky130_fd_sc_hd__or2_2
X_17472_ _17471_/X _17894_/X _17568_/S vssd1 vssd1 vccd1 vccd1 _17472_/X sky130_fd_sc_hd__mux2_1
XFILLER_232_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14684_ _14684_/A vssd1 vssd1 vccd1 vccd1 _14684_/X sky130_fd_sc_hd__clkbuf_2
X_11896_ _19419_/Q _11891_/X _09049_/X _11892_/X vssd1 vssd1 vccd1 vccd1 _19419_/D
+ sky130_fd_sc_hd__a22o_1
X_19211_ _19214_/CLK _19211_/D hold367/X vssd1 vssd1 vccd1 vccd1 _19211_/Q sky130_fd_sc_hd__dfrtp_1
X_16423_ _18241_/Q vssd1 vssd1 vccd1 vccd1 _16423_/Y sky130_fd_sc_hd__inv_2
XFILLER_232_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13635_ _13635_/A _13637_/A _13637_/B vssd1 vssd1 vccd1 vccd1 _13635_/X sky130_fd_sc_hd__or3_2
X_10847_ _19715_/Q _10843_/X _10448_/X _10845_/X vssd1 vssd1 vccd1 vccd1 _19715_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_220_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_repeater266_A repeater267/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19142_ _19582_/CLK _19142_/D hold348/A vssd1 vssd1 vccd1 vccd1 _19142_/Q sky130_fd_sc_hd__dfrtp_4
X_16354_ _18224_/Q vssd1 vssd1 vccd1 vccd1 _16354_/Y sky130_fd_sc_hd__inv_2
X_13566_ _13566_/A vssd1 vssd1 vccd1 vccd1 _13566_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17704__A1 _19756_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10778_ _17627_/X _10772_/X _19746_/Q _10774_/X vssd1 vssd1 vccd1 vccd1 _19746_/D
+ sky130_fd_sc_hd__a22o_1
X_15305_ _18632_/Q _18629_/Q _15305_/C vssd1 vssd1 vccd1 vccd1 _15305_/X sky130_fd_sc_hd__or3_2
XFILLER_12_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12517_ _19074_/Q _12512_/X hold256/X _12513_/X vssd1 vssd1 vccd1 vccd1 _19074_/D
+ sky130_fd_sc_hd__a22o_1
X_19073_ _19610_/CLK _19073_/D hold343/X vssd1 vssd1 vccd1 vccd1 _19073_/Q sky130_fd_sc_hd__dfrtp_1
X_16285_ _18263_/Q vssd1 vssd1 vccd1 vccd1 _16285_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12028__A _12028_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13497_ _14613_/A vssd1 vssd1 vccd1 vccd1 _13618_/B sky130_fd_sc_hd__inv_2
XFILLER_172_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18024_ _18142_/CLK _18024_/D vssd1 vssd1 vccd1 vccd1 _18024_/Q sky130_fd_sc_hd__dfxtp_1
X_15236_ _15227_/Y _18637_/Q _18636_/Q vssd1 vssd1 vccd1 vccd1 _15388_/B sky130_fd_sc_hd__a21oi_2
X_12448_ _19121_/Q _12441_/X _12384_/X _12444_/X vssd1 vssd1 vccd1 vccd1 _19121_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_154_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18623__SET_B hold351/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15167_ _17946_/Q _15159_/A _14713_/A _15160_/A vssd1 vssd1 vccd1 vccd1 _17946_/D
+ sky130_fd_sc_hd__a22o_1
X_12379_ _19157_/Q _12374_/X _12375_/X _12378_/X vssd1 vssd1 vccd1 vccd1 _19157_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_114_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19173__RESET_B hold370/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14118_ _14118_/A vssd1 vssd1 vccd1 vccd1 _14118_/X sky130_fd_sc_hd__buf_2
X_15098_ _17993_/Q _15095_/X _14802_/A _15097_/X vssd1 vssd1 vccd1 vccd1 _17993_/D
+ sky130_fd_sc_hd__a22o_1
X_19975_ _19984_/CLK _19975_/D repeater244/X vssd1 vssd1 vccd1 vccd1 _19975_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__16869__S _17548_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20078__RESET_B repeater205/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14049_ _14049_/A _14049_/B _14045_/X _14048_/X vssd1 vssd1 vccd1 vccd1 _14094_/A
+ sky130_fd_sc_hd__or4bb_4
X_18926_ _19283_/CLK _18926_/D repeater216/X vssd1 vssd1 vccd1 vccd1 _18926_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12701__B1 _12602_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_126_HCLK_A clkbuf_4_4_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20007__RESET_B repeater241/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18857_ _18866_/CLK _18857_/D repeater231/X vssd1 vssd1 vccd1 vccd1 _18857_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17866__S1 _18759_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12698__A _12698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09590_ _20023_/Q _09589_/Y _09585_/X _09484_/B vssd1 vssd1 vccd1 vccd1 _20023_/D
+ sky130_fd_sc_hd__o211a_1
X_17808_ _18475_/Q _18451_/Q _18459_/Q _18059_/Q _17918_/S0 _18750_/Q vssd1 vssd1
+ vccd1 vccd1 _17808_/X sky130_fd_sc_hd__mux4_1
X_18788_ _19647_/CLK _18788_/D repeater260/X vssd1 vssd1 vccd1 vccd1 _18788_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_95_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14454__B1 _14437_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17739_ _15370_/X _19706_/Q _18508_/D vssd1 vssd1 vccd1 vccd1 _17739_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16617__B _16621_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19409_ _19984_/CLK _19409_/D repeater243/X vssd1 vssd1 vccd1 vccd1 _19409_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_189_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19943__RESET_B repeater244/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16633__A _16633_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09024_ _20120_/Q _09015_/X hold288/X _09019_/X vssd1 vssd1 vccd1 vccd1 _20120_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_148_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_50_HCLK clkbuf_opt_1_HCLK/A vssd1 vssd1 vccd1 vccd1 _19780_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold220 hold220/A vssd1 vssd1 vccd1 vccd1 hold220/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold231 hold231/A vssd1 vssd1 vccd1 vccd1 hold231/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold242 input73/X vssd1 vssd1 vccd1 vccd1 hold242/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 hold253/A vssd1 vssd1 vccd1 vccd1 hold253/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11743__A1 _15749_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold264 input60/X vssd1 vssd1 vccd1 vccd1 hold264/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11743__B2 _11738_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12940__B1 _12937_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold275 sda_i_S4 vssd1 vssd1 vccd1 vccd1 input77/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold286 input57/X vssd1 vssd1 vccd1 vccd1 hold286/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16779__S _17513_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold297 HWDATA[23] vssd1 vssd1 vccd1 vccd1 input53/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20115_ _20115_/CLK _20115_/D repeater238/X vssd1 vssd1 vccd1 vccd1 _20115_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_172_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09926_ _19961_/Q _16649_/A _09869_/A _19353_/Q vssd1 vssd1 vccd1 vccd1 _09926_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_58_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_219_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20046_ _20048_/CLK _20046_/D repeater209/X vssd1 vssd1 vccd1 vccd1 _20046_/Q sky130_fd_sc_hd__dfrtp_1
X_09857_ _09857_/A _09857_/B _09857_/C vssd1 vssd1 vccd1 vccd1 _09858_/B sky130_fd_sc_hd__or3_1
XANTENNA__17857__S1 _18759_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18825__RESET_B repeater217/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_hold261_A HWDATA[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14445__B1 _14415_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12401__A hold315/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09788_ _09788_/A _09805_/A vssd1 vssd1 vccd1 vccd1 _09803_/A sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_48_HCLK_A clkbuf_opt_2_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17403__S _17567_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ _11771_/A vssd1 vssd1 vccd1 vccd1 _11750_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_242_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10701_ _19776_/Q vssd1 vssd1 vccd1 vccd1 _10701_/Y sky130_fd_sc_hd__inv_2
XFILLER_53_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11681_ _10525_/B _11674_/X _10516_/B _11675_/X vssd1 vssd1 vccd1 vccd1 _19536_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_230_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14328__A hold264/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13420_ _13528_/B vssd1 vssd1 vccd1 vccd1 _13443_/A sky130_fd_sc_hd__clkbuf_2
XPHY_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10632_ _10631_/Y _10598_/A _10617_/X _10595_/B _10618_/A vssd1 vssd1 vccd1 vccd1
+ _10633_/A sky130_fd_sc_hd__o32a_1
XPHY_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10563_ _10595_/A _10595_/D _19801_/Q _10595_/B vssd1 vssd1 vccd1 vccd1 _15297_/A
+ sky130_fd_sc_hd__and4bb_1
X_13351_ _13351_/A vssd1 vssd1 vccd1 vccd1 _13352_/C sky130_fd_sc_hd__inv_2
XFILLER_154_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17793__S0 _17923_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12302_ _14279_/A vssd1 vssd1 vccd1 vccd1 _12302_/X sky130_fd_sc_hd__buf_2
X_16070_ _16637_/A vssd1 vssd1 vccd1 vccd1 _16070_/X sky130_fd_sc_hd__buf_1
X_10494_ _19538_/Q _19537_/Q _19540_/Q _19539_/Q vssd1 vssd1 vccd1 vccd1 _11654_/B
+ sky130_fd_sc_hd__or4_4
X_13282_ _14247_/A vssd1 vssd1 vccd1 vccd1 _13746_/A sky130_fd_sc_hd__inv_2
XFILLER_154_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_182_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15021_ _18042_/Q _15011_/A _15020_/X _15012_/A vssd1 vssd1 vccd1 vccd1 _18042_/D
+ sky130_fd_sc_hd__a22o_1
X_12233_ _19231_/Q _12228_/X _12232_/X _12229_/X vssd1 vssd1 vccd1 vccd1 _19231_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_5_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12164_ _12171_/A vssd1 vssd1 vccd1 vccd1 _12164_/X sky130_fd_sc_hd__buf_1
XFILLER_162_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11115_ _19638_/Q _11114_/X _19638_/Q _11114_/X vssd1 vssd1 vccd1 vccd1 _19638_/D
+ sky130_fd_sc_hd__o2bb2a_1
X_16972_ _15963_/X _12741_/Y _17534_/S vssd1 vssd1 vccd1 vccd1 _16972_/X sky130_fd_sc_hd__mux2_1
X_19760_ _19772_/CLK _19760_/D repeater228/X vssd1 vssd1 vccd1 vccd1 _19760_/Q sky130_fd_sc_hd__dfrtp_1
X_12095_ hold315/X vssd1 vssd1 vccd1 vccd1 _12095_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_122_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11046_ _11039_/A _10266_/B _17752_/X _19645_/Q vssd1 vssd1 vccd1 vccd1 _19645_/D
+ sky130_fd_sc_hd__o22a_1
X_15923_ _17987_/Q vssd1 vssd1 vccd1 vccd1 _15923_/Y sky130_fd_sc_hd__inv_2
X_18711_ _18718_/CLK _18711_/D repeater253/X vssd1 vssd1 vccd1 vccd1 _18711_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_237_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19691_ _19772_/CLK _19691_/D repeater201/X vssd1 vssd1 vccd1 vccd1 _19691_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17848__S1 _18759_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15228__A2 _15226_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18642_ _18642_/CLK _18642_/D repeater219/X vssd1 vssd1 vccd1 vccd1 _18642_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__18566__RESET_B repeater271/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15854_ _15854_/A vssd1 vssd1 vccd1 vccd1 _15854_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_65_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10170__B1 _09079_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12311__A _15776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14805_ _18169_/Q _14801_/X _14802_/X _14804_/X vssd1 vssd1 vccd1 vccd1 _18169_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_206_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18573_ _19462_/CLK _18573_/D repeater273/X vssd1 vssd1 vccd1 vccd1 _18573_/Q sky130_fd_sc_hd__dfrtp_4
X_15785_ _18114_/Q vssd1 vssd1 vccd1 vccd1 _15785_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12997_ _12997_/A vssd1 vssd1 vccd1 vccd1 _12997_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17313__S _17564_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17524_ _17523_/X _09848_/A _17524_/S vssd1 vssd1 vccd1 vccd1 _17524_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14736_ _18208_/Q _14732_/X _14604_/X _14734_/X vssd1 vssd1 vccd1 vccd1 _18208_/D
+ sky130_fd_sc_hd__a22o_1
X_11948_ _11955_/A vssd1 vssd1 vccd1 vccd1 _11948_/X sky130_fd_sc_hd__buf_1
XFILLER_221_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_178_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17455_ _15768_/Y _14177_/Y _17546_/S vssd1 vssd1 vccd1 vccd1 _17455_/X sky130_fd_sc_hd__mux2_1
XFILLER_205_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14667_ _18765_/Q vssd1 vssd1 vccd1 vccd1 _15121_/A sky130_fd_sc_hd__buf_1
XFILLER_60_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11879_ _19432_/Q _11875_/X _09016_/X _11878_/X vssd1 vssd1 vccd1 vccd1 _19432_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_20_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16406_ _18169_/Q vssd1 vssd1 vccd1 vccd1 _16406_/Y sky130_fd_sc_hd__inv_2
X_13618_ _15195_/A _13618_/B vssd1 vssd1 vccd1 vccd1 _15193_/A sky130_fd_sc_hd__or2_1
X_17386_ _17385_/X _18808_/Q _17386_/S vssd1 vssd1 vccd1 vccd1 _17386_/X sky130_fd_sc_hd__mux2_2
XANTENNA__19508__CLK _19510_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14598_ _14598_/A _14598_/B _14598_/C vssd1 vssd1 vccd1 vccd1 _14601_/A sky130_fd_sc_hd__or3_4
Xclkbuf_leaf_73_HCLK clkbuf_opt_4_HCLK/A vssd1 vssd1 vccd1 vccd1 _18856_/CLK sky130_fd_sc_hd__clkbuf_16
X_19125_ _19208_/CLK _19125_/D hold370/X vssd1 vssd1 vccd1 vccd1 _19125_/Q sky130_fd_sc_hd__dfrtp_2
X_16337_ _18016_/Q vssd1 vssd1 vccd1 vccd1 _16337_/Y sky130_fd_sc_hd__inv_2
X_13549_ _13549_/A _13549_/B vssd1 vssd1 vccd1 vccd1 _13573_/A sky130_fd_sc_hd__or2_1
XFILLER_146_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19354__RESET_B hold370/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17784__S0 _19647_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19056_ _19157_/CLK _19056_/D repeater268/X vssd1 vssd1 vccd1 vccd1 _19056_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__15164__B2 _15160_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16268_ _19636_/Q _15936_/Y _19635_/Q _15799_/Y vssd1 vssd1 vccd1 vccd1 _16268_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_134_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18007_ _18416_/CLK _18007_/D vssd1 vssd1 vccd1 vccd1 _18007_/Q sky130_fd_sc_hd__dfxtp_1
X_15219_ _19722_/Q vssd1 vssd1 vccd1 vccd1 _15219_/Y sky130_fd_sc_hd__inv_2
XFILLER_114_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16199_ _17968_/Q _17967_/Q _17966_/Q _17965_/Q vssd1 vssd1 vccd1 vccd1 _16199_/Y
+ sky130_fd_sc_hd__nor4_2
XFILLER_142_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09067__A _12032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14124__C1 _14112_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19958_ _19964_/CLK _19958_/D hold373/X vssd1 vssd1 vccd1 vccd1 _19958_/Q sky130_fd_sc_hd__dfrtp_1
X_09711_ _09668_/A _09710_/Y _20002_/Q _19431_/Q vssd1 vssd1 vccd1 vccd1 _09711_/X
+ sky130_fd_sc_hd__a22o_1
X_18909_ _19293_/CLK _18909_/D repeater188/X vssd1 vssd1 vccd1 vccd1 _18909_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__17839__S1 _18761_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19889_ _20050_/CLK _19889_/D repeater206/X vssd1 vssd1 vccd1 vccd1 _19889_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_56_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13317__A _19260_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09642_ _19981_/Q vssd1 vssd1 vccd1 vccd1 _09793_/A sky130_fd_sc_hd__inv_2
XFILLER_110_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10161__B1 _09098_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14427__B1 _14351_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_243_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09573_ _09492_/A _09492_/B _09571_/Y _09604_/B vssd1 vssd1 vccd1 vccd1 _20032_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_82_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17223__S _17546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_224_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_224_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10676__A _10676_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17775__S0 _17923_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09007_ _19514_/Q _19513_/Q _19504_/Q vssd1 vssd1 vccd1 vccd1 _11832_/B sky130_fd_sc_hd__or3_1
XFILLER_247_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14666__B1 hold320/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_219_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09909_ _09857_/A _19341_/Q _09867_/A _19351_/Q vssd1 vssd1 vccd1 vccd1 _09909_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_120_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20029_ _20035_/CLK _20029_/D repeater240/X vssd1 vssd1 vccd1 vccd1 _20029_/Q sky130_fd_sc_hd__dfrtp_1
X_12920_ _19291_/Q _18948_/Q _19291_/Q _18948_/Q vssd1 vssd1 vccd1 vccd1 _12920_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_19_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10152__A0 _10147_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14418__B1 _14417_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12851_ _18933_/Q vssd1 vssd1 vccd1 vccd1 _12964_/C sky130_fd_sc_hd__inv_2
XPHY_4021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15091__B1 hold263/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_215_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11970__A _11979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17133__S _17543_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11802_ _19460_/Q _11800_/X hold314/X _11801_/X vssd1 vssd1 vccd1 vccd1 _19460_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15570_ _18586_/Q _15566_/A _15569_/Y _15566_/Y vssd1 vssd1 vccd1 vccd1 _15571_/B
+ sky130_fd_sc_hd__o22a_1
XPHY_4065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12782_ _12777_/Y _18822_/Q _19233_/Q _13534_/A _12781_/X vssd1 vssd1 vccd1 vccd1
+ _12783_/D sky130_fd_sc_hd__o221a_1
XPHY_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_96_HCLK clkbuf_4_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19964_/CLK sky130_fd_sc_hd__clkbuf_16
Xrebuffer90 _09850_/B vssd1 vssd1 vccd1 vccd1 _10002_/B1 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_4087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14521_ _18329_/Q _14518_/X _14437_/X _14520_/X vssd1 vssd1 vccd1 vccd1 _18329_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11733_ _19504_/Q _11730_/X _16936_/X _11731_/X vssd1 vssd1 vccd1 vccd1 hold227/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16972__S _17534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_214_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17240_ _17239_/X _11439_/Y _17548_/S vssd1 vssd1 vccd1 vccd1 _17240_/X sky130_fd_sc_hd__mux2_1
XFILLER_186_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14452_ _14452_/A vssd1 vssd1 vccd1 vccd1 _14453_/A sky130_fd_sc_hd__inv_2
XPHY_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11664_ _18520_/Q _11668_/A vssd1 vssd1 vccd1 vccd1 _11675_/A sky130_fd_sc_hd__or2_1
XPHY_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13403_ _20103_/Q vssd1 vssd1 vccd1 vccd1 _13403_/Y sky130_fd_sc_hd__inv_4
XFILLER_186_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10615_ _10615_/A _10933_/B _10942_/C vssd1 vssd1 vccd1 vccd1 _10616_/D sky130_fd_sc_hd__or3_2
X_17171_ _17170_/X _13403_/Y _17535_/S vssd1 vssd1 vccd1 vccd1 _17171_/X sky130_fd_sc_hd__mux2_1
XPHY_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14383_ _18409_/Q _14380_/X _12714_/X _14382_/X vssd1 vssd1 vccd1 vccd1 _18409_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_128_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11595_ _19573_/Q _11594_/Y _11547_/B _11594_/A _11588_/X vssd1 vssd1 vccd1 vccd1
+ _19573_/D sky130_fd_sc_hd__o221a_1
XPHY_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17766__S0 _17923_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16122_ _19028_/Q vssd1 vssd1 vccd1 vccd1 _16122_/Y sky130_fd_sc_hd__inv_2
XPHY_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13334_ _13464_/A _13463_/C _13334_/C _13334_/D vssd1 vssd1 vccd1 vccd1 _13431_/A
+ sky130_fd_sc_hd__or4_4
X_10546_ _19808_/Q _19807_/Q _10572_/C vssd1 vssd1 vccd1 vccd1 _10557_/C sky130_fd_sc_hd__or3_1
XFILLER_41_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_2_HCLK clkbuf_4_0_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _18165_/CLK sky130_fd_sc_hd__clkbuf_16
X_16053_ _16053_/A vssd1 vssd1 vccd1 vccd1 _16053_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_155_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13265_ _18753_/Q vssd1 vssd1 vccd1 vccd1 _13274_/B sky130_fd_sc_hd__inv_2
X_10477_ _17701_/X _10471_/X _19818_/Q _10472_/X vssd1 vssd1 vccd1 vccd1 _19818_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_repeater229_A repeater230/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15004_ _18954_/Q vssd1 vssd1 vccd1 vccd1 _15004_/X sky130_fd_sc_hd__buf_2
XFILLER_124_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12216_ _19241_/Q _12212_/X _12028_/X _12213_/X vssd1 vssd1 vccd1 vccd1 _19241_/D
+ sky130_fd_sc_hd__a22o_1
X_13196_ _13196_/A vssd1 vssd1 vccd1 vccd1 _13199_/A sky130_fd_sc_hd__inv_2
XFILLER_123_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16720__B _16721_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19812_ _19812_/CLK _19812_/D repeater222/X vssd1 vssd1 vccd1 vccd1 _19812_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17308__S _17566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_0_HCLK_A HCLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12147_ _12147_/A1 _12143_/X _12088_/X _12144_/X vssd1 vssd1 vccd1 vccd1 _19286_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_151_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19743_ _20070_/CLK _19743_/D repeater207/X vssd1 vssd1 vccd1 vccd1 _19743_/Q sky130_fd_sc_hd__dfrtp_1
X_16955_ _17789_/X _18793_/Q _16957_/S vssd1 vssd1 vccd1 vccd1 _16955_/X sky130_fd_sc_hd__mux2_1
X_12078_ hold279/X vssd1 vssd1 vccd1 vccd1 _12078_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__13137__A _19169_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11029_ _11029_/A _11029_/B vssd1 vssd1 vccd1 vccd1 _11029_/Y sky130_fd_sc_hd__nand2_1
X_15906_ _17542_/X _15896_/X _17530_/X _15898_/X _15905_/X vssd1 vssd1 vccd1 vccd1
+ _15918_/C sky130_fd_sc_hd__o221a_2
XFILLER_238_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19674_ _19822_/CLK _19674_/D repeater218/X vssd1 vssd1 vccd1 vccd1 _19674_/Q sky130_fd_sc_hd__dfrtp_1
X_16886_ _16885_/X _15572_/Y _17513_/S vssd1 vssd1 vccd1 vccd1 _16886_/X sky130_fd_sc_hd__mux2_1
XFILLER_225_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18625_ _19814_/CLK _18625_/D repeater223/X vssd1 vssd1 vccd1 vccd1 _18625_/Q sky130_fd_sc_hd__dfrtp_1
X_15837_ _19693_/Q vssd1 vssd1 vccd1 vccd1 _15837_/Y sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_31_HCLK_A _18641_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17043__S _17474_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15768_ _15863_/B vssd1 vssd1 vccd1 vccd1 _15768_/Y sky130_fd_sc_hd__clkinv_16
X_18556_ _20066_/CLK _18556_/D repeater193/X vssd1 vssd1 vccd1 vccd1 _18556_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12435__A2 _12400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_94_HCLK_A clkbuf_4_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_221_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17507_ _17506_/X _12058_/A _17567_/S vssd1 vssd1 vccd1 vccd1 _17507_/X sky130_fd_sc_hd__mux2_1
X_14719_ _14719_/A vssd1 vssd1 vccd1 vccd1 _14719_/X sky130_fd_sc_hd__clkbuf_2
X_18487_ _19812_/CLK _18487_/D repeater222/X vssd1 vssd1 vccd1 vccd1 _18489_/D sky130_fd_sc_hd__dfstp_1
XFILLER_33_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15699_ _15697_/Y _15698_/X _15673_/X vssd1 vssd1 vccd1 vccd1 _15699_/X sky130_fd_sc_hd__o21a_1
XANTENNA__16882__S _17522_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19535__RESET_B repeater221/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_221_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17438_ _17437_/X _17884_/X _17568_/S vssd1 vssd1 vccd1 vccd1 _17438_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_193_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17369_ _16298_/Y _09324_/Y _19498_/Q vssd1 vssd1 vccd1 vccd1 _17369_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19108_ _19109_/CLK _19108_/D hold343/X vssd1 vssd1 vccd1 vccd1 _19108_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_174_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19039_ _19041_/CLK _19039_/D repeater266/X vssd1 vssd1 vccd1 vccd1 _19039_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_174_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20093__RESET_B repeater233/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput100 _16728_/X vssd1 vssd1 vccd1 vccd1 HRDATA[29] sky130_fd_sc_hd__clkbuf_2
Xoutput111 _18623_/Q vssd1 vssd1 vccd1 vccd1 HREADYOUT sky130_fd_sc_hd__clkbuf_2
Xoutput122 _15750_/X vssd1 vssd1 vccd1 vccd1 IRQ[4] sky130_fd_sc_hd__clkbuf_2
Xoutput133 _20038_/Q vssd1 vssd1 vccd1 vccd1 SCLK_S3 sky130_fd_sc_hd__clkbuf_2
XFILLER_126_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput144 _19671_/Q vssd1 vssd1 vccd1 vccd1 sda_oen_o_S4 sky130_fd_sc_hd__clkbuf_2
XFILLER_88_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17218__S _17542_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09625_ _09787_/B vssd1 vssd1 vccd1 vccd1 _09807_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__11882__B1 _09025_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09556_ _19319_/Q vssd1 vssd1 vccd1 vccd1 _09556_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09260__A _12370_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09487_ _09487_/A _09580_/A vssd1 vssd1 vccd1 vccd1 _09488_/B sky130_fd_sc_hd__or2_2
XANTENNA__16792__S _17490_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10400_ _10404_/A _10400_/B vssd1 vssd1 vccd1 vccd1 _10400_/X sky130_fd_sc_hd__or2_1
XFILLER_165_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11380_ _19138_/Q vssd1 vssd1 vccd1 vccd1 _11380_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19973__CLK _19984_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16325__B1 _17359_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10331_ _10331_/A _10340_/A vssd1 vssd1 vccd1 vccd1 _10332_/B sky130_fd_sc_hd__or2_1
XFILLER_109_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10262_ _15070_/A vssd1 vssd1 vccd1 vccd1 _14517_/A sky130_fd_sc_hd__buf_1
XFILLER_3_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13050_ _18896_/Q vssd1 vssd1 vccd1 vccd1 _13069_/B sky130_fd_sc_hd__inv_2
X_12001_ _12043_/A vssd1 vssd1 vccd1 vccd1 _12044_/A sky130_fd_sc_hd__inv_2
XANTENNA__15437__A _19773_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18840__RESET_B repeater233/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17128__S _17517_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_239_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10193_ _18796_/Q vssd1 vssd1 vccd1 vccd1 _13637_/A sky130_fd_sc_hd__inv_2
XFILLER_133_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17920__S0 _17923_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16967__S _17459_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16740_ _16793_/X _16509_/X _16837_/X _15896_/X _16739_/X vssd1 vssd1 vccd1 vccd1
+ _16743_/B sky130_fd_sc_hd__o221a_2
X_13952_ _18715_/Q _13951_/Y _13925_/A _13815_/B vssd1 vssd1 vccd1 vccd1 _18715_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_207_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12903_ _19283_/Q _12964_/A _12902_/Y _18946_/Q vssd1 vssd1 vccd1 vccd1 _12903_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_234_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16671_ _16671_/A _16718_/B vssd1 vssd1 vccd1 vccd1 _16671_/Y sky130_fd_sc_hd__nor2_1
X_13883_ _19204_/Q vssd1 vssd1 vccd1 vccd1 _13883_/Y sky130_fd_sc_hd__inv_2
XFILLER_235_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15622_ _15622_/A _15622_/B vssd1 vssd1 vccd1 vccd1 _15622_/Y sky130_fd_sc_hd__nor2_1
X_18410_ _18412_/CLK _18410_/D vssd1 vssd1 vccd1 vccd1 _18410_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16800__A1 _18916_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12834_ _12834_/A _12834_/B _12834_/C _12834_/D vssd1 vssd1 vccd1 vccd1 _13588_/A
+ sky130_fd_sc_hd__and4_2
X_19390_ _19933_/CLK _19390_/D repeater235/X vssd1 vssd1 vccd1 vccd1 _19390_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_62_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18341_ _18473_/CLK _18341_/D vssd1 vssd1 vccd1 vccd1 _18341_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15553_ _15557_/B _15552_/Y _15542_/X vssd1 vssd1 vccd1 vccd1 _15553_/X sky130_fd_sc_hd__o21a_1
X_12765_ _19257_/Q vssd1 vssd1 vccd1 vccd1 _12765_/Y sky130_fd_sc_hd__inv_2
XPHY_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_repeater179_A _17414_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14504_ _14504_/A vssd1 vssd1 vccd1 vccd1 _14505_/A sky130_fd_sc_hd__inv_2
XFILLER_203_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18272_ _20081_/CLK _18272_/D vssd1 vssd1 vccd1 vccd1 _18272_/Q sky130_fd_sc_hd__dfxtp_1
X_11716_ _11730_/A vssd1 vssd1 vccd1 vccd1 _11716_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_187_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15484_ _15487_/B _15482_/X _15483_/X vssd1 vssd1 vccd1 vccd1 _15484_/X sky130_fd_sc_hd__o21a_1
X_12696_ _18968_/Q _12691_/X hold259/X _12692_/X vssd1 vssd1 vccd1 vccd1 _18968_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16715__B _16715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17223_ _15768_/Y _14191_/Y _17546_/S vssd1 vssd1 vccd1 vccd1 _17223_/X sky130_fd_sc_hd__mux2_1
XPHY_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14435_ _14450_/A _14450_/B _14598_/C vssd1 vssd1 vccd1 vccd1 _14438_/A sky130_fd_sc_hd__or3_4
XPHY_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11647_ _15389_/A vssd1 vssd1 vccd1 vccd1 _11647_/Y sky130_fd_sc_hd__inv_2
XANTENNA__09046__A1 _20111_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput13 input13/A vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__clkbuf_1
XPHY_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput24 HADDR[30] vssd1 vssd1 vccd1 vccd1 input24/X sky130_fd_sc_hd__buf_1
X_17154_ _17153_/X _19953_/Q _17518_/S vssd1 vssd1 vccd1 vccd1 _17154_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput35 input35/A vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_hd__buf_1
XPHY_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14366_ _14366_/A _14366_/B _14784_/C vssd1 vssd1 vccd1 vccd1 _14368_/A sky130_fd_sc_hd__or3_4
XANTENNA__12050__B1 _11924_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11578_ _11578_/A _11606_/A vssd1 vssd1 vccd1 vccd1 _11579_/B sky130_fd_sc_hd__or2_2
Xinput46 input46/A vssd1 vssd1 vccd1 vccd1 input46/X sky130_fd_sc_hd__clkbuf_4
Xinput57 input57/A vssd1 vssd1 vccd1 vccd1 input57/X sky130_fd_sc_hd__buf_4
Xinput68 input68/A vssd1 vssd1 vccd1 vccd1 input68/X sky130_fd_sc_hd__clkbuf_4
X_16105_ _18133_/Q vssd1 vssd1 vccd1 vccd1 _16105_/Y sky130_fd_sc_hd__inv_2
X_13317_ _19260_/Q vssd1 vssd1 vccd1 vccd1 _13462_/A sky130_fd_sc_hd__inv_2
XFILLER_156_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10529_ _11649_/B _11651_/B _10529_/C _11653_/B vssd1 vssd1 vccd1 vccd1 _10532_/C
+ sky130_fd_sc_hd__or4_4
X_17085_ _17084_/X _14046_/Y _17544_/S vssd1 vssd1 vccd1 vccd1 _17085_/X sky130_fd_sc_hd__mux2_1
X_14297_ _18451_/Q _14289_/A _13680_/X _14290_/A vssd1 vssd1 vccd1 vccd1 _18451_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_171_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16036_ _18260_/Q vssd1 vssd1 vccd1 vccd1 _16036_/Y sky130_fd_sc_hd__inv_2
X_13248_ _18875_/Q _13241_/X _12536_/X _13243_/X vssd1 vssd1 vccd1 vccd1 _18875_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_143_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_103_HCLK clkbuf_4_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19293_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_131_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17038__S _17318_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18581__RESET_B repeater274/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11875__A _11891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13179_ _13179_/A vssd1 vssd1 vccd1 vccd1 _13179_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_229_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17911__S0 _17913_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16877__S _17529_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17987_ _19851_/CLK _17987_/D vssd1 vssd1 vccd1 vccd1 _17987_/Q sky130_fd_sc_hd__dfxtp_1
X_19726_ _20051_/CLK _19726_/D repeater207/X vssd1 vssd1 vccd1 vccd1 _19726_/Q sky130_fd_sc_hd__dfrtp_1
X_16938_ _19482_/Q hold162/X _16946_/S vssd1 vssd1 vccd1 vccd1 _16938_/X sky130_fd_sc_hd__mux2_1
XFILLER_96_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19787__RESET_B repeater203/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_237_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19657_ _19668_/CLK _19657_/D repeater270/X vssd1 vssd1 vccd1 vccd1 _19657_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__15055__B1 _15004_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16869_ _16868_/X _11415_/Y _17548_/S vssd1 vssd1 vccd1 vccd1 _16869_/X sky130_fd_sc_hd__mux2_1
X_09410_ _19908_/Q vssd1 vssd1 vccd1 vccd1 _10011_/B sky130_fd_sc_hd__inv_2
X_18608_ _19566_/CLK _18608_/D repeater255/X vssd1 vssd1 vccd1 vccd1 _18608_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_92_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19588_ _19610_/CLK _19588_/D hold343/X vssd1 vssd1 vccd1 vccd1 _19588_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_240_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09341_ _09339_/X _20037_/Q _09342_/S vssd1 vssd1 vccd1 vccd1 _20037_/D sky130_fd_sc_hd__mux2_1
X_18539_ _19825_/CLK _18539_/D repeater229/X vssd1 vssd1 vccd1 vccd1 _18539_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17501__S _17566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_221_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09272_ _20057_/Q _09269_/X _09082_/X _09271_/X vssd1 vssd1 vccd1 vccd1 _20057_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_20_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_221_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11919__A1 _19405_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12041__B1 _11911_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11785__A _11821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17902__S0 _17913_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09255__A _12313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16787__S _17473_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08987_ _10133_/A _08986_/Y _10132_/B _08986_/A vssd1 vssd1 vccd1 vccd1 _20123_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_69_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_3_7_0_HCLK_A clkbuf_3_7_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19457__RESET_B repeater272/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09608_ _09473_/A _09473_/B _09605_/Y _09607_/X vssd1 vssd1 vccd1 vccd1 _20012_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_113_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10880_ _15364_/A _10875_/X _10877_/X _10879_/X vssd1 vssd1 vccd1 vccd1 _19700_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_73_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09539_ _09489_/A _19319_/Q _09475_/A _19305_/Q vssd1 vssd1 vccd1 vccd1 _09539_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_189_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17411__S _17518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12550_ _12550_/A vssd1 vssd1 vccd1 vccd1 _19060_/D sky130_fd_sc_hd__inv_2
XPHY_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12280__B1 _12100_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_237_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11501_ _19603_/Q _11500_/Y _11490_/X _11484_/B vssd1 vssd1 vccd1 vccd1 _19603_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_185_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12481_ _19098_/Q _12478_/X _12302_/X _12479_/X vssd1 vssd1 vccd1 vccd1 _19098_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14220_ _14166_/X _14184_/X _14219_/X _18671_/Q _14112_/A vssd1 vssd1 vccd1 vccd1
+ _18671_/D sky130_fd_sc_hd__a32o_1
XPHY_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11432_ _19571_/Q _11428_/Y _19560_/Q _11429_/Y _11431_/X vssd1 vssd1 vccd1 vccd1
+ _11433_/D sky130_fd_sc_hd__o221a_1
XPHY_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_126_HCLK clkbuf_4_4_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19157_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_137_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14151_ _19122_/Q vssd1 vssd1 vccd1 vccd1 _16717_/A sky130_fd_sc_hd__inv_2
XFILLER_125_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11363_ _11523_/A vssd1 vssd1 vccd1 vccd1 _11521_/A sky130_fd_sc_hd__inv_2
XFILLER_152_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13102_ _19182_/Q vssd1 vssd1 vccd1 vccd1 _16667_/A sky130_fd_sc_hd__inv_2
X_10314_ _17928_/Q _10314_/B vssd1 vssd1 vccd1 vccd1 _10314_/X sky130_fd_sc_hd__and2_2
X_14082_ _19073_/Q _14014_/A _19081_/Q _14022_/A vssd1 vssd1 vccd1 vccd1 _14082_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_3_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11294_ _19001_/Q vssd1 vssd1 vccd1 vccd1 _11294_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17910_ _15782_/Y _15783_/Y _15784_/Y _15785_/Y _17913_/S0 _19632_/Q vssd1 vssd1
+ vccd1 vccd1 _17910_/X sky130_fd_sc_hd__mux4_2
XFILLER_98_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13033_ _18913_/Q vssd1 vssd1 vccd1 vccd1 _13085_/A sky130_fd_sc_hd__inv_2
X_10245_ _10240_/Y _19655_/Q _19828_/Q _10956_/C _10244_/X vssd1 vssd1 vccd1 vccd1
+ _10246_/D sky130_fd_sc_hd__o221a_1
XFILLER_78_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18890_ _19352_/CLK _18890_/D hold372/X vssd1 vssd1 vccd1 vccd1 _18890_/Q sky130_fd_sc_hd__dfrtp_1
X_17841_ _16402_/Y _16403_/Y _16404_/Y _16405_/Y _17913_/S0 _19632_/Q vssd1 vssd1
+ vccd1 vccd1 _17841_/X sky130_fd_sc_hd__mux4_2
X_10176_ _19882_/Q _10174_/X _09094_/X _10175_/X vssd1 vssd1 vccd1 vccd1 _19882_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14088__A1 _19069_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16482__C1 _16481_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12099__B1 _12098_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17772_ _18323_/Q _18003_/Q _18307_/Q _18299_/Q _17923_/S0 _19646_/Q vssd1 vssd1
+ vccd1 vccd1 _17772_/X sky130_fd_sc_hd__mux4_2
X_14984_ _18063_/Q _14976_/X hold244/X _14979_/X vssd1 vssd1 vccd1 vccd1 _18063_/D
+ sky130_fd_sc_hd__a22o_1
X_19511_ _19513_/CLK hold220/X repeater259/X vssd1 vssd1 vccd1 vccd1 _19511_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_219_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16723_ _19054_/Q _16723_/B vssd1 vssd1 vccd1 vccd1 _16723_/Y sky130_fd_sc_hd__nand2_1
X_13935_ _13935_/A vssd1 vssd1 vccd1 vccd1 _13935_/Y sky130_fd_sc_hd__inv_2
XFILLER_247_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11310__A2 _18991_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16654_ _17076_/X _16594_/X _16907_/X _16595_/X vssd1 vssd1 vccd1 vccd1 _16656_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_74_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19442_ _20064_/CLK _19442_/D repeater193/X vssd1 vssd1 vccd1 vccd1 _19442_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_235_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13866_ _13863_/Y _18704_/Q _13864_/Y _18719_/Q _13865_/X vssd1 vssd1 vccd1 vccd1
+ _13867_/D sky130_fd_sc_hd__o221a_1
XANTENNA__16785__A0 _17473_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15605_ _15605_/A vssd1 vssd1 vccd1 vccd1 _15605_/Y sky130_fd_sc_hd__inv_2
X_12817_ _18805_/Q vssd1 vssd1 vccd1 vccd1 _13529_/A sky130_fd_sc_hd__inv_2
X_19373_ _19971_/CLK _19373_/D repeater191/X vssd1 vssd1 vccd1 vccd1 _19373_/Q sky130_fd_sc_hd__dfrtp_1
X_16585_ _16585_/A _16615_/B vssd1 vssd1 vccd1 vccd1 _16585_/Y sky130_fd_sc_hd__nor2_1
X_13797_ _19125_/Q vssd1 vssd1 vccd1 vccd1 _13964_/A sky130_fd_sc_hd__inv_2
XANTENNA__17321__S _17543_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18324_ _18431_/CLK _18324_/D vssd1 vssd1 vccd1 vccd1 _18324_/Q sky130_fd_sc_hd__dfxtp_1
X_15536_ _18578_/Q vssd1 vssd1 vccd1 vccd1 _15536_/Y sky130_fd_sc_hd__inv_2
XFILLER_203_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12748_ _18833_/Q vssd1 vssd1 vccd1 vccd1 _13556_/A sky130_fd_sc_hd__clkinvlp_2
XANTENNA__12271__B1 _12083_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18255_ _20077_/CLK _18255_/D vssd1 vssd1 vccd1 vccd1 _18255_/Q sky130_fd_sc_hd__dfxtp_1
X_15467_ _15467_/A _15467_/B vssd1 vssd1 vccd1 vccd1 _15467_/Y sky130_fd_sc_hd__nor2_1
XPHY_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12679_ _18981_/Q _12677_/X hold315/X _12678_/X vssd1 vssd1 vccd1 vccd1 _18981_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_8_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17206_ _15963_/X _09497_/Y _17543_/S vssd1 vssd1 vccd1 vccd1 _17206_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14418_ _18389_/Q _14409_/X _14417_/X _14411_/X vssd1 vssd1 vccd1 vccd1 _18389_/D
+ sky130_fd_sc_hd__a22o_1
X_18186_ _18460_/CLK _18186_/D vssd1 vssd1 vccd1 vccd1 _18186_/Q sky130_fd_sc_hd__dfxtp_1
X_15398_ _15402_/A _17581_/X vssd1 vssd1 vccd1 vccd1 _18531_/D sky130_fd_sc_hd__and2_1
XANTENNA__11377__A2 _19132_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17137_ _17136_/X _15493_/Y _17513_/S vssd1 vssd1 vccd1 vccd1 _17137_/X sky130_fd_sc_hd__mux2_1
XFILLER_156_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14349_ _14352_/A vssd1 vssd1 vccd1 vccd1 _14349_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__18762__RESET_B repeater195/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17068_ _17067_/X _20024_/Q _17482_/S vssd1 vssd1 vccd1 vccd1 _17068_/X sky130_fd_sc_hd__mux2_2
X_16019_ _18340_/Q vssd1 vssd1 vccd1 vccd1 _16019_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09890_ _09874_/A _19358_/Q _19953_/Q _16548_/A _09889_/X vssd1 vssd1 vccd1 vccd1
+ _09895_/C sky130_fd_sc_hd__o221a_1
XFILLER_112_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09075__A hold250/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14079__A1 _19082_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_214_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19709_ _19720_/CLK _19709_/D repeater201/X vssd1 vssd1 vccd1 vccd1 _19709_/Q sky130_fd_sc_hd__dfstp_1
XPHY_4609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10949__A _10949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15028__B1 _14998_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_0_0_HCLK_A clkbuf_4_1_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19550__RESET_B repeater269/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_230_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17231__S _17546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09324_ _20045_/Q vssd1 vssd1 vccd1 vccd1 _09324_/Y sky130_fd_sc_hd__inv_2
XFILLER_167_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_149_HCLK clkbuf_4_1_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19867_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_159_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09255_ _12313_/A vssd1 vssd1 vccd1 vccd1 _09255_/X sky130_fd_sc_hd__buf_2
XANTENNA__10684__A _11842_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12014__B1 _09037_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14554__A2 _14547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09186_ _20074_/Q _09164_/A _09185_/X _09165_/A vssd1 vssd1 vccd1 vccd1 _20074_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_119_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12404__A hold301/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10030_ _10030_/A vssd1 vssd1 vccd1 vccd1 _10051_/B sky130_fd_sc_hd__inv_2
XFILLER_103_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19638__RESET_B repeater258/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16464__C1 _16462_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17406__S _17513_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_187_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11828__B1 _10868_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11981_ _14279_/A vssd1 vssd1 vccd1 vccd1 _11981_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__15019__B1 _15006_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13720_ _13708_/Y _13719_/X _13708_/Y _13719_/X vssd1 vssd1 vccd1 vccd1 _13721_/D
+ sky130_fd_sc_hd__a2bb2o_1
X_10932_ _17728_/X _10923_/A _19673_/Q _10924_/A vssd1 vssd1 vccd1 vccd1 _19673_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18146__CLK _19851_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13651_ _16953_/X _13644_/A _18790_/Q _13646_/X vssd1 vssd1 vccd1 vccd1 _18790_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_232_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10863_ _12234_/A vssd1 vssd1 vccd1 vccd1 _10863_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_220_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17141__S _17546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12602_ _14279_/A vssd1 vssd1 vccd1 vccd1 _12602_/X sky130_fd_sc_hd__buf_4
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16370_ _19031_/Q vssd1 vssd1 vccd1 vccd1 _16370_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13582_ _13545_/A _13545_/B _13571_/X _13580_/Y vssd1 vssd1 vccd1 vccd1 _18822_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_169_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10794_ _19738_/Q _10794_/B _19733_/Q vssd1 vssd1 vccd1 vccd1 _10807_/A sky130_fd_sc_hd__or3b_4
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15321_ _15321_/A _15321_/B vssd1 vssd1 vccd1 vccd1 _15321_/Y sky130_fd_sc_hd__nor2_1
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12533_ hold325/X vssd1 vssd1 vccd1 vccd1 _12533_/X sky130_fd_sc_hd__buf_4
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18040_ _19851_/CLK _18040_/D vssd1 vssd1 vccd1 vccd1 _18040_/Q sky130_fd_sc_hd__dfxtp_1
X_15252_ _18629_/Q vssd1 vssd1 vccd1 vccd1 _15256_/A sky130_fd_sc_hd__inv_2
XANTENNA__12005__B1 _09021_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12464_ _12478_/A vssd1 vssd1 vccd1 vccd1 _12464_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_172_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14203_ _19108_/Q vssd1 vssd1 vccd1 vccd1 _14203_/Y sky130_fd_sc_hd__inv_2
X_11415_ _19145_/Q vssd1 vssd1 vccd1 vccd1 _11415_/Y sky130_fd_sc_hd__inv_2
X_15183_ _18488_/D _10658_/C _18489_/D _17936_/Q _15182_/X vssd1 vssd1 vccd1 vccd1
+ _17936_/D sky130_fd_sc_hd__a32o_1
X_12395_ _19150_/Q _12388_/X _12394_/X _12390_/X vssd1 vssd1 vccd1 vccd1 _19150_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09421__B2 _09420_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08999__A _15890_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14134_ _14012_/B _14134_/A2 _14012_/A vssd1 vssd1 vccd1 vccd1 _14135_/C sky130_fd_sc_hd__o21a_1
X_11346_ _19588_/Q _11344_/Y _11463_/A _18964_/Q _11345_/X vssd1 vssd1 vccd1 vccd1
+ _11347_/D sky130_fd_sc_hd__o221a_1
X_19991_ _19992_/CLK _19991_/D repeater192/X vssd1 vssd1 vccd1 vccd1 _19991_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_165_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14065_ _19071_/Q vssd1 vssd1 vccd1 vccd1 _14065_/Y sky130_fd_sc_hd__inv_2
XANTENNA_repeater211_A repeater212/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18942_ _18947_/CLK _18942_/D repeater213/X vssd1 vssd1 vccd1 vccd1 _18942_/Q sky130_fd_sc_hd__dfrtp_1
X_11277_ _19580_/Q vssd1 vssd1 vccd1 vccd1 _11461_/A sky130_fd_sc_hd__inv_2
XANTENNA__12314__A _15774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13016_ _13004_/A _13004_/B _13014_/Y _12986_/A vssd1 vssd1 vccd1 vccd1 _18925_/D
+ sky130_fd_sc_hd__a211oi_2
X_10228_ _10226_/Y _19663_/Q _10227_/Y _19656_/Q vssd1 vssd1 vccd1 vccd1 _10228_/X
+ sky130_fd_sc_hd__o22a_1
X_18873_ _20049_/CLK _18873_/D repeater208/X vssd1 vssd1 vccd1 vccd1 _18873_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_95_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19379__RESET_B repeater230/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17316__S _17564_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17824_ _17820_/X _17821_/X _17822_/X _17823_/X _18751_/Q _18752_/Q vssd1 vssd1 vccd1
+ vccd1 _17824_/X sky130_fd_sc_hd__mux4_2
X_10159_ _19893_/Q _10154_/X _09090_/X _10156_/X vssd1 vssd1 vccd1 vccd1 _19893_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_181_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11819__B1 _09079_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14967_ _18073_/Q _14964_/X _14802_/X _14966_/X vssd1 vssd1 vccd1 vccd1 _18073_/D
+ sky130_fd_sc_hd__a22o_1
X_17755_ _17754_/S _11059_/Y _17755_/S vssd1 vssd1 vccd1 vccd1 _17755_/X sky130_fd_sc_hd__mux2_2
XFILLER_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16706_ _20119_/Q vssd1 vssd1 vccd1 vccd1 _16706_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13918_ _18731_/Q _13917_/Y _13830_/B _13917_/A _13901_/X vssd1 vssd1 vccd1 vccd1
+ _18731_/D sky130_fd_sc_hd__o221a_1
X_17686_ _15488_/X _19449_/Q _17696_/S vssd1 vssd1 vccd1 vccd1 _18566_/D sky130_fd_sc_hd__mux2_1
X_14898_ _14898_/A vssd1 vssd1 vccd1 vccd1 _14898_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_62_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19425_ _19997_/CLK _19425_/D repeater274/X vssd1 vssd1 vccd1 vccd1 _19425_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_222_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16637_ _16637_/A vssd1 vssd1 vccd1 vccd1 _16637_/X sky130_fd_sc_hd__clkbuf_2
X_13849_ _19199_/Q _13947_/A _19213_/Q _13909_/B vssd1 vssd1 vccd1 vccd1 _13849_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__15360__A _15364_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17051__S _17548_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19356_ _19968_/CLK _19356_/D hold371/X vssd1 vssd1 vccd1 vccd1 _19356_/Q sky130_fd_sc_hd__dfrtp_1
X_16568_ _16504_/X _16562_/X _16565_/X _16567_/X vssd1 vssd1 vccd1 vccd1 _16568_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_31_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18307_ _19847_/CLK _18307_/D vssd1 vssd1 vccd1 vccd1 _18307_/Q sky130_fd_sc_hd__dfxtp_1
X_15519_ _15523_/B vssd1 vssd1 vccd1 vccd1 _15526_/B sky130_fd_sc_hd__inv_2
XANTENNA__16890__S _17544_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16499_ _16487_/X _16504_/A _16492_/X _16496_/X _16498_/X vssd1 vssd1 vccd1 vccd1
+ _16499_/Y sky130_fd_sc_hd__o2111ai_4
X_19287_ _19288_/CLK _19287_/D repeater211/X vssd1 vssd1 vccd1 vccd1 _19287_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_200_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09040_ _20113_/Q _09029_/X _09039_/X _09031_/X vssd1 vssd1 vccd1 vccd1 _20113_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_148_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_149_HCLK_A clkbuf_4_1_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18238_ _20077_/CLK _18238_/D vssd1 vssd1 vccd1 vccd1 _18238_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_190_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18169_ _18169_/CLK _18169_/D vssd1 vssd1 vccd1 vccd1 _18169_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09942_ _19347_/Q vssd1 vssd1 vccd1 vccd1 _09942_/Y sky130_fd_sc_hd__inv_2
XANTENNA__09715__A2 _19418_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20062_ _20064_/CLK _20062_/D repeater200/X vssd1 vssd1 vccd1 vccd1 _20062_/Q sky130_fd_sc_hd__dfrtp_1
X_09873_ _09873_/A _09873_/B vssd1 vssd1 vccd1 vccd1 _09957_/A sky130_fd_sc_hd__or2_1
XFILLER_100_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17226__S _17473_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16997__A0 _15963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater230 repeater233/X vssd1 vssd1 vccd1 vccd1 repeater230/X sky130_fd_sc_hd__buf_8
XANTENNA__10730__B1 _10427_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater241 repeater242/X vssd1 vssd1 vccd1 vccd1 repeater241/X sky130_fd_sc_hd__buf_8
XFILLER_239_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18169__CLK _18169_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater252 repeater253/X vssd1 vssd1 vccd1 vccd1 repeater252/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__11782__B _11933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrepeater263 repeater266/X vssd1 vssd1 vccd1 vccd1 repeater263/X sky130_fd_sc_hd__buf_6
XFILLER_54_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrepeater274 hold348/A vssd1 vssd1 vccd1 vccd1 repeater274/X sky130_fd_sc_hd__buf_8
XFILLER_241_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater285 hold354/A vssd1 vssd1 vccd1 vccd1 hold356/A sky130_fd_sc_hd__buf_6
XFILLER_38_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12483__B1 _12234_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_242_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_214_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12235__B1 _12234_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold137_A HADDR[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09307_ _20049_/Q _15727_/A _20049_/Q _15727_/A vssd1 vssd1 vccd1 vccd1 _09333_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_70_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18684__RESET_B repeater252/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09238_ _09238_/A _09238_/B vssd1 vssd1 vccd1 vccd1 _15712_/A sky130_fd_sc_hd__or2_1
XANTENNA_hold304_A HWDATA[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14527__A2 _14519_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09169_ _14703_/A _09163_/X _09168_/X _09165_/X vssd1 vssd1 vccd1 vccd1 _20080_/D
+ sky130_fd_sc_hd__a22o_1
X_11200_ _19010_/Q vssd1 vssd1 vccd1 vccd1 _11200_/Y sky130_fd_sc_hd__inv_2
XFILLER_107_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12180_ _12313_/A vssd1 vssd1 vccd1 vccd1 _12180_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11131_ _19630_/Q vssd1 vssd1 vccd1 vccd1 _12253_/A sky130_fd_sc_hd__inv_2
XFILLER_134_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09706__A2 _19405_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11062_ _19632_/Q vssd1 vssd1 vccd1 vccd1 _11064_/A sky130_fd_sc_hd__inv_2
XFILLER_122_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19472__RESET_B repeater260/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10013_ _10013_/A vssd1 vssd1 vccd1 vccd1 _10101_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__17136__S _17512_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15445__A _15571_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15870_ _18951_/Q vssd1 vssd1 vccd1 vccd1 _15870_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_209_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19401__RESET_B hold371/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input22_A HADDR[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14821_ _14821_/A vssd1 vssd1 vccd1 vccd1 _14822_/A sky130_fd_sc_hd__inv_2
XFILLER_236_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16975__S _17544_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14752_ _18199_/Q _14744_/X _14751_/X _14747_/X vssd1 vssd1 vccd1 vccd1 _18199_/D
+ sky130_fd_sc_hd__a22o_1
X_17540_ _17539_/X _13135_/Y _17543_/S vssd1 vssd1 vccd1 vccd1 _17540_/X sky130_fd_sc_hd__mux2_1
X_11964_ _19382_/Q _11962_/X hold276/X _11963_/X vssd1 vssd1 vccd1 vccd1 _19382_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_17_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12474__B1 _12356_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13703_ _17761_/X vssd1 vssd1 vccd1 vccd1 _13706_/A sky130_fd_sc_hd__inv_2
X_10915_ _19683_/Q _10914_/A _10913_/Y _10914_/Y _18510_/Q vssd1 vssd1 vccd1 vccd1
+ _19683_/D sky130_fd_sc_hd__a221o_1
XFILLER_17_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17471_ _17470_/X _11093_/Y _17567_/S vssd1 vssd1 vccd1 vccd1 _17471_/X sky130_fd_sc_hd__mux2_1
XFILLER_204_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14683_ _14683_/A vssd1 vssd1 vccd1 vccd1 _14684_/A sky130_fd_sc_hd__inv_2
XFILLER_71_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11895_ _19420_/Q _11891_/X hold317/X _11892_/X vssd1 vssd1 vccd1 vccd1 _19420_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_output109_A _16482_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19210_ _19214_/CLK _19210_/D hold367/X vssd1 vssd1 vccd1 vccd1 _19210_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__12226__B1 _12225_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13634_ _13634_/A vssd1 vssd1 vccd1 vccd1 _18799_/D sky130_fd_sc_hd__inv_2
XFILLER_60_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16422_ _18257_/Q vssd1 vssd1 vccd1 vccd1 _16422_/Y sky130_fd_sc_hd__inv_2
X_10846_ _19716_/Q _10843_/X _10446_/X _10845_/X vssd1 vssd1 vccd1 vccd1 _19716_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_44_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_232_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19141_ _19561_/CLK _19141_/D repeater274/X vssd1 vssd1 vccd1 vccd1 _19141_/Q sky130_fd_sc_hd__dfrtp_4
X_16353_ _18240_/Q vssd1 vssd1 vccd1 vccd1 _16353_/Y sky130_fd_sc_hd__inv_2
X_13565_ _13555_/A _13555_/B _13597_/A _13563_/Y vssd1 vssd1 vccd1 vccd1 _18832_/D
+ sky130_fd_sc_hd__a211oi_2
X_10777_ _17626_/X _10772_/X _19747_/Q _10774_/X vssd1 vssd1 vccd1 vccd1 _19747_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_repeater161_A _17547_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater259_A repeater260/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12309__A _12309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15304_ _15304_/A _15305_/C vssd1 vssd1 vccd1 vccd1 _15304_/Y sky130_fd_sc_hd__nand2_1
XFILLER_157_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12516_ _19075_/Q _12512_/X hold281/X _12513_/X vssd1 vssd1 vccd1 vccd1 _19075_/D
+ sky130_fd_sc_hd__a22o_1
X_19072_ _19610_/CLK _19072_/D hold343/X vssd1 vssd1 vccd1 vccd1 _19072_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_200_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16284_ _18079_/Q vssd1 vssd1 vccd1 vccd1 _16284_/Y sky130_fd_sc_hd__inv_2
XFILLER_185_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13496_ _18836_/Q _15320_/A _13496_/C vssd1 vssd1 vccd1 vccd1 _14613_/A sky130_fd_sc_hd__or3_1
X_18023_ _18145_/CLK _18023_/D vssd1 vssd1 vccd1 vccd1 _18023_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15235_ _18622_/D vssd1 vssd1 vccd1 vccd1 _18624_/D sky130_fd_sc_hd__buf_1
XFILLER_172_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18641__D _18641_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12447_ _19122_/Q _12441_/X _12382_/X _12444_/X vssd1 vssd1 vccd1 vccd1 _19122_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_output90_A _16006_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15166_ _17947_/Q _15159_/A _14711_/A _15160_/A vssd1 vssd1 vccd1 vccd1 _17947_/D
+ sky130_fd_sc_hd__a22o_1
X_12378_ _12402_/A vssd1 vssd1 vccd1 vccd1 _12378_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_125_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14117_ _18693_/Q _14115_/Y _14116_/X _14117_/C1 vssd1 vssd1 vccd1 vccd1 _18693_/D
+ sky130_fd_sc_hd__o211a_1
X_11329_ _11468_/A _18970_/Q _11478_/A _18980_/Q vssd1 vssd1 vccd1 vccd1 _11329_/X
+ sky130_fd_sc_hd__o22a_1
X_15097_ _15097_/A vssd1 vssd1 vccd1 vccd1 _15097_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_99_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19974_ _19984_/CLK _19974_/D repeater244/X vssd1 vssd1 vccd1 vccd1 _19974_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_141_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14048_ _14046_/Y _18679_/Q _19066_/Q _14008_/A _14047_/X vssd1 vssd1 vccd1 vccd1
+ _14048_/X sky130_fd_sc_hd__o221a_1
X_18925_ _19283_/CLK _18925_/D repeater211/X vssd1 vssd1 vccd1 vccd1 _18925_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_122_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_228_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17046__S _17546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18856_ _18856_/CLK _18856_/D repeater231/X vssd1 vssd1 vccd1 vccd1 _18856_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_95_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19142__RESET_B hold348/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17807_ _18355_/Q _17995_/Q _18411_/Q _18395_/Q _17918_/S0 _18750_/Q vssd1 vssd1
+ vccd1 vccd1 _17807_/X sky130_fd_sc_hd__mux4_2
Xclkbuf_4_4_0_HCLK clkbuf_4_5_0_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_4_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_18787_ _19865_/CLK _18787_/D repeater263/X vssd1 vssd1 vccd1 vccd1 _18787_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__16885__S _17512_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15999_ _15999_/A vssd1 vssd1 vccd1 vccd1 _15999_/X sky130_fd_sc_hd__buf_2
XFILLER_236_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17738_ _15371_/X _19707_/Q _18508_/D vssd1 vssd1 vccd1 vccd1 _17738_/X sky130_fd_sc_hd__mux2_1
XFILLER_208_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20047__RESET_B repeater208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_224_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17669_ _15560_/X _19466_/Q _17683_/S vssd1 vssd1 vccd1 vccd1 _18583_/D sky130_fd_sc_hd__mux2_1
XFILLER_196_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19408_ _19984_/CLK _19408_/D repeater193/X vssd1 vssd1 vccd1 vccd1 _19408_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12217__B1 _12030_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17156__A0 _15963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19339_ _19352_/CLK _19339_/D repeater245/X vssd1 vssd1 vccd1 vccd1 _19339_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12219__A _12228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09023_ hold289/X vssd1 vssd1 vccd1 vccd1 hold288/A sky130_fd_sc_hd__buf_4
Xhold210 input37/X vssd1 vssd1 vccd1 vccd1 hold210/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__19983__RESET_B repeater192/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold221 hold221/A vssd1 vssd1 vccd1 vccd1 hold221/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold232 hold232/A vssd1 vssd1 vccd1 vccd1 hold232/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_160_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold243 RsRx_S0 vssd1 vssd1 vccd1 vccd1 input73/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11743__A2 _11737_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12940__A1 _12936_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold254 input75/X vssd1 vssd1 vccd1 vccd1 hold254/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold265 HWDATA[2] vssd1 vssd1 vccd1 vccd1 input60/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold276 hold276/A vssd1 vssd1 vccd1 vccd1 hold276/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold287 HWDATA[27] vssd1 vssd1 vccd1 vccd1 input57/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20114_ _20120_/CLK _20114_/D repeater217/X vssd1 vssd1 vccd1 vccd1 _20114_/Q sky130_fd_sc_hd__dfrtp_4
Xhold298 input52/X vssd1 vssd1 vccd1 vccd1 hold298/X sky130_fd_sc_hd__dlygate4sd3_1
X_09925_ _19353_/Q vssd1 vssd1 vccd1 vccd1 _16649_/A sky130_fd_sc_hd__inv_2
XFILLER_59_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11793__A _11800_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20045_ _20048_/CLK _20045_/D repeater209/X vssd1 vssd1 vccd1 vccd1 _20045_/Q sky130_fd_sc_hd__dfrtp_1
X_09856_ _09856_/A _09856_/B vssd1 vssd1 vccd1 vccd1 _09857_/C sky130_fd_sc_hd__or2_2
XFILLER_219_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16795__S _17545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09787_ _09807_/A _09787_/B _09787_/C vssd1 vssd1 vccd1 vccd1 _09805_/A sky130_fd_sc_hd__or3_1
XFILLER_45_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12456__B1 _12398_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18865__RESET_B repeater233/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10700_ _18879_/Q vssd1 vssd1 vccd1 vccd1 _15404_/A sky130_fd_sc_hd__clkbuf_2
XPHY_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12208__B1 _12098_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ _19537_/Q _11668_/X _11652_/B _11669_/X vssd1 vssd1 vccd1 vccd1 _19537_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10631_ _18554_/Q vssd1 vssd1 vccd1 vccd1 _10631_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17147__A0 _17486_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13350_ _13350_/A _13350_/B vssd1 vssd1 vccd1 vccd1 _13351_/A sky130_fd_sc_hd__or2_1
XFILLER_167_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10562_ _19802_/Q vssd1 vssd1 vccd1 vccd1 _10595_/B sky130_fd_sc_hd__inv_2
XANTENNA__11431__B2 _19155_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16543__B _16544_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12301_ _19199_/Q _12298_/X _12299_/X _12300_/X vssd1 vssd1 vccd1 vccd1 _19199_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_194_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17793__S1 _19646_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_132_HCLK_A clkbuf_4_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13281_ _18869_/Q _13654_/A _15190_/A vssd1 vssd1 vccd1 vccd1 _14247_/A sky130_fd_sc_hd__or3_4
X_10493_ _10493_/A _10493_/B vssd1 vssd1 vccd1 vccd1 _10736_/B sky130_fd_sc_hd__nand2_1
X_15020_ _18952_/Q vssd1 vssd1 vccd1 vccd1 _15020_/X sky130_fd_sc_hd__buf_2
XFILLER_6_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12232_ _12232_/A vssd1 vssd1 vccd1 vccd1 _12232_/X sky130_fd_sc_hd__buf_4
XFILLER_108_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12163_ _19274_/Q _12157_/X _12032_/X _12158_/X vssd1 vssd1 vccd1 vccd1 _19274_/D
+ sky130_fd_sc_hd__a22o_1
X_11114_ _11091_/X _11113_/B _17754_/S _11113_/Y _17755_/X vssd1 vssd1 vccd1 vccd1
+ _11114_/X sky130_fd_sc_hd__o221a_1
X_12094_ _12094_/A vssd1 vssd1 vccd1 vccd1 _12094_/X sky130_fd_sc_hd__clkbuf_2
X_16971_ _16970_/X _09873_/A _17524_/S vssd1 vssd1 vccd1 vccd1 _16971_/X sky130_fd_sc_hd__mux2_1
XFILLER_77_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08996__B _12130_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18710_ _18718_/CLK _18710_/D repeater253/X vssd1 vssd1 vccd1 vccd1 _18710_/Q sky130_fd_sc_hd__dfrtp_1
X_15922_ _18115_/Q vssd1 vssd1 vccd1 vccd1 _15922_/Y sky130_fd_sc_hd__inv_2
X_11045_ _17752_/X _10268_/B _11044_/X vssd1 vssd1 vccd1 vccd1 _19646_/D sky130_fd_sc_hd__a21oi_1
XFILLER_39_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19690_ _19772_/CLK _19690_/D repeater201/X vssd1 vssd1 vccd1 vccd1 _19690_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12695__B1 hold267/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18641_ _18641_/CLK _18641_/D repeater204/X vssd1 vssd1 vccd1 vccd1 _18641_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_37_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15853_ _18872_/Q vssd1 vssd1 vccd1 vccd1 _15853_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12311__B _12316_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14804_ _14804_/A vssd1 vssd1 vccd1 vccd1 _14804_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__12447__B1 _12382_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18572_ _19462_/CLK _18572_/D repeater273/X vssd1 vssd1 vccd1 vccd1 _18572_/Q sky130_fd_sc_hd__dfrtp_1
X_12996_ _12964_/C _12875_/B _12994_/Y _12986_/X vssd1 vssd1 vccd1 vccd1 _18933_/D
+ sky130_fd_sc_hd__a211oi_2
X_15784_ _18026_/Q vssd1 vssd1 vccd1 vccd1 _15784_/Y sky130_fd_sc_hd__inv_2
XFILLER_91_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16718__B _16718_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17523_ _17522_/X _09680_/Y _17523_/S vssd1 vssd1 vccd1 vccd1 _17523_/X sky130_fd_sc_hd__mux2_1
X_11947_ _19393_/Q _11939_/X _09027_/X _11942_/X vssd1 vssd1 vccd1 vccd1 _19393_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_45_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14735_ _18209_/Q _14732_/X _14600_/X _14734_/X vssd1 vssd1 vccd1 vccd1 _18209_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14519__A _14519_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_221_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14666_ _18242_/Q _14657_/A hold320/X _14658_/A vssd1 vssd1 vccd1 vccd1 _18242_/D
+ sky130_fd_sc_hd__a22o_1
X_17454_ _17453_/X _13062_/A _17488_/S vssd1 vssd1 vccd1 vccd1 _17454_/X sky130_fd_sc_hd__mux2_1
X_11878_ _11892_/A vssd1 vssd1 vccd1 vccd1 _11878_/X sky130_fd_sc_hd__clkbuf_2
X_16405_ _18057_/Q vssd1 vssd1 vccd1 vccd1 _16405_/Y sky130_fd_sc_hd__inv_2
X_13617_ _13617_/A vssd1 vssd1 vccd1 vccd1 _13617_/Y sky130_fd_sc_hd__inv_2
X_10829_ _19720_/Q vssd1 vssd1 vccd1 vccd1 _10829_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_4_12_0_HCLK clkbuf_3_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_12_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
X_17385_ _16211_/Y _20095_/Q _17385_/S vssd1 vssd1 vccd1 vccd1 _17385_/X sky130_fd_sc_hd__mux2_1
X_14597_ _18282_/Q _14588_/A hold320/X _14589_/A vssd1 vssd1 vccd1 vccd1 _18282_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_186_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19124_ _19609_/CLK _19124_/D hold355/X vssd1 vssd1 vccd1 vccd1 _19124_/Q sky130_fd_sc_hd__dfrtp_1
X_13548_ _13548_/A _13577_/A vssd1 vssd1 vccd1 vccd1 _13549_/B sky130_fd_sc_hd__or2_1
X_16336_ _18168_/Q vssd1 vssd1 vccd1 vccd1 _16336_/Y sky130_fd_sc_hd__inv_2
XFILLER_173_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17784__S1 _19648_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11878__A _11892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19055_ _19577_/CLK _19055_/D repeater268/X vssd1 vssd1 vccd1 vccd1 _19055_/Q sky130_fd_sc_hd__dfrtp_1
X_16267_ _18047_/Q vssd1 vssd1 vccd1 vccd1 _16267_/Y sky130_fd_sc_hd__inv_2
X_13479_ _13479_/A vssd1 vssd1 vccd1 vccd1 _13479_/Y sky130_fd_sc_hd__inv_2
XFILLER_173_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15164__A2 _15158_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15218_ _18638_/Q vssd1 vssd1 vccd1 vccd1 _15218_/Y sky130_fd_sc_hd__inv_2
X_18006_ _18416_/CLK _18006_/D vssd1 vssd1 vccd1 vccd1 _18006_/Q sky130_fd_sc_hd__dfxtp_1
X_16198_ _18748_/Q _16114_/Y _16043_/Y _16196_/Y vssd1 vssd1 vccd1 vccd1 _16198_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_142_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_54_HCLK_A clkbuf_opt_2_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15149_ _17960_/Q _15146_/X _14699_/A _15148_/X vssd1 vssd1 vccd1 vccd1 _17960_/D
+ sky130_fd_sc_hd__a22o_1
X_19957_ _19965_/CLK _19957_/D hold371/X vssd1 vssd1 vccd1 vccd1 _19957_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_68_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_206_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09710_ _19431_/Q vssd1 vssd1 vccd1 vccd1 _09710_/Y sky130_fd_sc_hd__inv_2
XFILLER_101_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18908_ _18908_/CLK _18908_/D repeater188/X vssd1 vssd1 vccd1 vccd1 _18908_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_206_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12686__B1 hold277/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19888_ _20050_/CLK _19888_/D repeater206/X vssd1 vssd1 vccd1 vccd1 _19888_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_28_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09641_ _09791_/A _09790_/A _09789_/A _09807_/A vssd1 vssd1 vccd1 vccd1 _09647_/C
+ sky130_fd_sc_hd__or4_4
X_18839_ _20107_/CLK _18839_/D repeater233/X vssd1 vssd1 vccd1 vccd1 _18839_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_56_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_243_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_222_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17504__S _17564_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12438__A0 _12313_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09572_ _20033_/Q _09571_/Y _09567_/X _09494_/B vssd1 vssd1 vccd1 vccd1 _20033_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_243_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18546__D _18546_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12610__A0 _12313_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17775__S1 _19646_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09006_ _10186_/A _10430_/A vssd1 vssd1 vccd1 vccd1 _10842_/A sky130_fd_sc_hd__or2_4
XANTENNA__14363__B1 _14329_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09258__A _19516_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15560__C1 _15512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19752__CLK _19900_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09908_ _19337_/Q vssd1 vssd1 vccd1 vccd1 _09908_/Y sky130_fd_sc_hd__inv_2
XFILLER_116_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09839_ _19947_/Q vssd1 vssd1 vccd1 vccd1 _09856_/A sky130_fd_sc_hd__inv_2
X_20028_ _20035_/CLK _20028_/D repeater242/X vssd1 vssd1 vccd1 vccd1 _20028_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_47_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12131__B _15895_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17414__S _17414_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11028__A _19873_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12850_ _18934_/Q vssd1 vssd1 vccd1 vccd1 _12876_/A sky130_fd_sc_hd__inv_2
XANTENNA__12429__B1 _12299_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11801_ _11801_/A vssd1 vssd1 vccd1 vccd1 _11801_/X sky130_fd_sc_hd__buf_1
XPHY_4044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12781_ _12779_/Y _18814_/Q _16619_/A _18824_/Q vssd1 vssd1 vccd1 vccd1 _12781_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_4055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer80 _14032_/B vssd1 vssd1 vccd1 vccd1 _14100_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_4077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14520_ _14520_/A vssd1 vssd1 vccd1 vccd1 _14520_/X sky130_fd_sc_hd__clkbuf_2
Xrebuffer91 _09850_/B vssd1 vssd1 vccd1 vccd1 _10000_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_4088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11732_ _19505_/Q _11730_/X _16937_/X _11731_/X vssd1 vssd1 vccd1 vccd1 hold221/A
+ sky130_fd_sc_hd__a22o_1
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14451_ _14452_/A vssd1 vssd1 vccd1 vccd1 _14451_/X sky130_fd_sc_hd__clkbuf_2
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11663_ _11674_/A vssd1 vssd1 vccd1 vccd1 _11668_/A sky130_fd_sc_hd__inv_2
XPHY_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13402_ _13389_/X _13402_/B _13402_/C _13402_/D vssd1 vssd1 vccd1 vccd1 _13418_/C
+ sky130_fd_sc_hd__and4b_1
XPHY_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10614_ _10614_/A _10614_/B _10614_/C vssd1 vssd1 vccd1 vccd1 _10942_/C sky130_fd_sc_hd__or3_1
X_17170_ _15963_/X _12793_/Y _17534_/S vssd1 vssd1 vccd1 vccd1 _17170_/X sky130_fd_sc_hd__mux2_1
XPHY_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12601__B1 _12599_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11404__B2 _19147_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14382_ _14382_/A vssd1 vssd1 vccd1 vccd1 _14382_/X sky130_fd_sc_hd__clkbuf_2
XPHY_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11594_ _11594_/A vssd1 vssd1 vccd1 vccd1 _11594_/Y sky130_fd_sc_hd__inv_2
XPHY_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16121_ _19442_/Q vssd1 vssd1 vccd1 vccd1 _16121_/Y sky130_fd_sc_hd__inv_2
X_13333_ _13469_/A _13468_/A _13333_/C _13470_/A vssd1 vssd1 vccd1 vccd1 _13334_/D
+ sky130_fd_sc_hd__or4_4
XFILLER_195_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17766__S1 _19646_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10545_ _19802_/Q _19801_/Q _10561_/A vssd1 vssd1 vccd1 vccd1 _10572_/C sky130_fd_sc_hd__or3_1
XFILLER_194_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16052_ _19695_/Q vssd1 vssd1 vccd1 vccd1 _16052_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14354__B1 _14351_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13264_ _13255_/Y _13263_/X _13255_/Y _13263_/X vssd1 vssd1 vccd1 vccd1 _13278_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_10476_ _17700_/X _10471_/X _19819_/Q _10472_/X vssd1 vssd1 vccd1 vccd1 _19819_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_170_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15003_ _18053_/Q _14991_/X _15002_/X _14994_/X vssd1 vssd1 vccd1 vccd1 _18053_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_124_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12215_ _19242_/Q _12212_/X _12026_/X _12213_/X vssd1 vssd1 vccd1 vccd1 _19242_/D
+ sky130_fd_sc_hd__a22o_1
X_13195_ _13071_/A _13195_/A2 _13193_/Y _13182_/X vssd1 vssd1 vccd1 vccd1 _18899_/D
+ sky130_fd_sc_hd__a211oi_2
X_19811_ _19812_/CLK _19811_/D repeater222/X vssd1 vssd1 vccd1 vccd1 _19811_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_123_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12146_ _19287_/Q _12143_/X _12086_/X _12144_/X vssd1 vssd1 vccd1 vccd1 _19287_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_111_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19742_ _20070_/CLK _19742_/D repeater207/X vssd1 vssd1 vccd1 vccd1 _19742_/Q sky130_fd_sc_hd__dfrtp_1
X_12077_ _19323_/Q _12068_/X _12076_/X _12072_/X vssd1 vssd1 vccd1 vccd1 _19323_/D
+ sky130_fd_sc_hd__a22o_1
X_16954_ _17784_/X _18792_/Q _16957_/S vssd1 vssd1 vccd1 vccd1 _16954_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12668__B1 hold279/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11028_ _19873_/Q _15294_/A vssd1 vssd1 vccd1 vccd1 _11029_/B sky130_fd_sc_hd__or2_1
X_15905_ _17568_/X _16506_/A _17548_/X _15904_/X vssd1 vssd1 vccd1 vccd1 _15905_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_110_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19673_ _19822_/CLK _19673_/D repeater218/X vssd1 vssd1 vccd1 vccd1 _19673_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_64_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16885_ _17473_/A0 _16737_/Y _17512_/S vssd1 vssd1 vccd1 vccd1 _16885_/X sky130_fd_sc_hd__mux2_1
XANTENNA__17324__S _17534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18624_ _19867_/CLK _18624_/D repeater262/X vssd1 vssd1 vccd1 vccd1 _18624_/Q sky130_fd_sc_hd__dfrtp_1
X_15836_ _15836_/A vssd1 vssd1 vccd1 vccd1 _15836_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__18716__RESET_B repeater253/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_225_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_40_HCLK clkbuf_opt_1_HCLK/A vssd1 vssd1 vccd1 vccd1 _19813_/CLK sky130_fd_sc_hd__clkbuf_16
X_18555_ _19810_/CLK _18555_/D repeater226/X vssd1 vssd1 vccd1 vccd1 _18555_/Q sky130_fd_sc_hd__dfrtp_1
X_15767_ _18871_/Q _18514_/Q vssd1 vssd1 vccd1 vccd1 _15767_/X sky130_fd_sc_hd__and2_2
X_12979_ _13060_/B vssd1 vssd1 vccd1 vccd1 _12980_/A sky130_fd_sc_hd__clkbuf_2
X_17506_ _17505_/X _10218_/Y _17566_/S vssd1 vssd1 vccd1 vccd1 _17506_/X sky130_fd_sc_hd__mux2_1
XFILLER_233_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14718_ _14718_/A vssd1 vssd1 vccd1 vccd1 _14719_/A sky130_fd_sc_hd__inv_2
X_18486_ _19812_/CLK _18486_/D repeater222/X vssd1 vssd1 vccd1 vccd1 _18488_/D sky130_fd_sc_hd__dfstp_2
XFILLER_221_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15698_ _18616_/Q _15693_/A _18617_/Q vssd1 vssd1 vccd1 vccd1 _15698_/X sky130_fd_sc_hd__o21a_1
X_17437_ _17436_/X _11059_/Y _17567_/S vssd1 vssd1 vccd1 vccd1 _17437_/X sky130_fd_sc_hd__mux2_1
XFILLER_221_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19625__CLK _19920_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14649_ _18254_/Q _14643_/X _09177_/X _14645_/X vssd1 vssd1 vccd1 vccd1 _18254_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_221_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17368_ _17367_/X _11381_/Y _17548_/S vssd1 vssd1 vccd1 vccd1 _17368_/X sky130_fd_sc_hd__mux2_1
XANTENNA__19575__RESET_B hold346/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19107_ _19109_/CLK _19107_/D hold343/X vssd1 vssd1 vccd1 vccd1 _19107_/Q sky130_fd_sc_hd__dfrtp_1
X_16319_ _16311_/Y _15828_/X _16313_/X _16318_/X vssd1 vssd1 vccd1 vccd1 _16319_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_119_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17299_ _15963_/X _12799_/Y _17534_/S vssd1 vssd1 vccd1 vccd1 _17299_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14345__B1 _14312_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19038_ _19867_/CLK _19038_/D repeater263/X vssd1 vssd1 vccd1 vccd1 _19038_/Q sky130_fd_sc_hd__dfrtp_1
Xoutput101 _16077_/Y vssd1 vssd1 vccd1 vccd1 HRDATA[2] sky130_fd_sc_hd__clkbuf_2
XFILLER_173_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput112 _16747_/Y vssd1 vssd1 vccd1 vccd1 IRQ[0] sky130_fd_sc_hd__clkbuf_2
Xoutput123 _15767_/X vssd1 vssd1 vccd1 vccd1 IRQ[5] sky130_fd_sc_hd__clkbuf_2
Xoutput134 _15731_/Y vssd1 vssd1 vccd1 vccd1 SSn_S2 sky130_fd_sc_hd__clkbuf_2
Xoutput145 _19764_/Q vssd1 vssd1 vccd1 vccd1 sda_oen_o_S5 sky130_fd_sc_hd__clkbuf_2
XFILLER_99_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12232__A _12232_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17234__S _17543_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09624_ _19364_/Q vssd1 vssd1 vccd1 vccd1 _09787_/B sky130_fd_sc_hd__inv_2
XANTENNA__11882__A1 _19429_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09555_ _19302_/Q vssd1 vssd1 vccd1 vccd1 _16471_/A sky130_fd_sc_hd__inv_2
XFILLER_71_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10687__A _15839_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09260__B _12130_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_212_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09486_ _09486_/A _09486_/B vssd1 vssd1 vccd1 vccd1 _09580_/A sky130_fd_sc_hd__or2_1
XPHY_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14584__B1 _14567_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16325__B2 _16003_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10330_ _10330_/A _10343_/A vssd1 vssd1 vccd1 vccd1 _10340_/A sky130_fd_sc_hd__or2_1
XFILLER_164_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17409__S _17543_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10261_ _19644_/Q vssd1 vssd1 vccd1 vccd1 _15070_/A sky130_fd_sc_hd__inv_2
XFILLER_3_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12000_ _12016_/A vssd1 vssd1 vccd1 vccd1 _12000_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_121_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10192_ _18797_/Q vssd1 vssd1 vccd1 vccd1 _13635_/A sky130_fd_sc_hd__inv_2
XFILLER_239_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17920__S1 _19646_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_219_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_63_HCLK clkbuf_opt_3_HCLK/A vssd1 vssd1 vccd1 vccd1 _20091_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_247_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13951_ _13951_/A _13951_/B vssd1 vssd1 vccd1 vccd1 _13951_/Y sky130_fd_sc_hd__nor2_2
XFILLER_46_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17144__S _17534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11981__A _14279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12902_ _19289_/Q vssd1 vssd1 vccd1 vccd1 _12902_/Y sky130_fd_sc_hd__inv_2
X_13882_ _13882_/A _13882_/B _13882_/C _13882_/D vssd1 vssd1 vccd1 vccd1 _13898_/C
+ sky130_fd_sc_hd__and4_1
X_16670_ _16670_/A _16718_/B vssd1 vssd1 vccd1 vccd1 _16670_/Y sky130_fd_sc_hd__nor2_1
XFILLER_235_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12833_ _12833_/A _12833_/B _12833_/C _12833_/D vssd1 vssd1 vccd1 vccd1 _12834_/D
+ sky130_fd_sc_hd__and4_1
X_15621_ _15621_/A vssd1 vssd1 vccd1 vccd1 _15621_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18340_ _18954_/CLK _18340_/D vssd1 vssd1 vccd1 vccd1 _18340_/Q sky130_fd_sc_hd__dfxtp_1
X_12764_ _19229_/Q _13530_/A _12760_/Y _18806_/Q _12763_/X vssd1 vssd1 vccd1 vccd1
+ _12764_/X sky130_fd_sc_hd__a221o_1
X_15552_ _15552_/A _15552_/B vssd1 vssd1 vccd1 vccd1 _15552_/Y sky130_fd_sc_hd__nor2_1
XPHY_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11715_ _19516_/Q _11708_/X _16948_/X _16950_/S vssd1 vssd1 vccd1 vccd1 hold215/A
+ sky130_fd_sc_hd__a22o_1
X_14503_ _14504_/A vssd1 vssd1 vccd1 vccd1 _14503_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_15483_ _15512_/A vssd1 vssd1 vccd1 vccd1 _15483_/X sky130_fd_sc_hd__clkbuf_2
X_18271_ _20077_/CLK _18271_/D vssd1 vssd1 vccd1 vccd1 _18271_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12695_ _18969_/Q _12691_/X hold267/X _12692_/X vssd1 vssd1 vccd1 vccd1 _18969_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16564__B2 _16683_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17222_ _16484_/X _10226_/Y _17566_/S vssd1 vssd1 vccd1 vccd1 _17222_/X sky130_fd_sc_hd__mux2_1
XPHY_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14434_ _18378_/Q _14425_/A _14405_/X _14426_/A vssd1 vssd1 vccd1 vccd1 _18378_/D
+ sky130_fd_sc_hd__a22o_1
X_11646_ _11639_/A _11639_/B _19546_/Q _11567_/A _11588_/X vssd1 vssd1 vccd1 vccd1
+ _19546_/D sky130_fd_sc_hd__o221a_1
XPHY_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09450__A1_N _10039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput14 input14/A vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__buf_1
XPHY_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14365_ _18418_/Q _14352_/A _14314_/X _14353_/A vssd1 vssd1 vccd1 vccd1 _18418_/D
+ sky130_fd_sc_hd__a22o_1
Xinput25 HADDR[31] vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__buf_1
XPHY_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17153_ _16548_/Y _19415_/Q _17541_/S vssd1 vssd1 vccd1 vccd1 _17153_/X sky130_fd_sc_hd__mux2_1
XFILLER_183_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11577_ _11577_/A _11577_/B vssd1 vssd1 vccd1 vccd1 _11606_/A sky130_fd_sc_hd__or2_1
Xinput36 HTRANS[0] vssd1 vssd1 vccd1 vccd1 input36/X sky130_fd_sc_hd__buf_1
XPHY_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12050__B2 _12017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput47 input47/A vssd1 vssd1 vccd1 vccd1 input47/X sky130_fd_sc_hd__clkbuf_4
X_13316_ _18849_/Q vssd1 vssd1 vccd1 vccd1 _13428_/D sky130_fd_sc_hd__inv_6
XFILLER_155_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14327__B1 _14326_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput58 input58/A vssd1 vssd1 vccd1 vccd1 input58/X sky130_fd_sc_hd__buf_4
X_16104_ _18221_/Q vssd1 vssd1 vccd1 vccd1 _16104_/Y sky130_fd_sc_hd__inv_2
X_10528_ _10505_/C _19537_/Q _10528_/C vssd1 vssd1 vccd1 vccd1 _11653_/B sky130_fd_sc_hd__and3b_1
Xinput69 input69/A vssd1 vssd1 vccd1 vccd1 input69/X sky130_fd_sc_hd__clkbuf_4
X_17084_ _15768_/Y _14155_/Y _17546_/S vssd1 vssd1 vccd1 vccd1 _17084_/X sky130_fd_sc_hd__mux2_1
X_14296_ _18452_/Q _14289_/A _13678_/X _14290_/A vssd1 vssd1 vccd1 vccd1 _18452_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_143_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13247_ _18876_/Q _13241_/X _12533_/X _13243_/X vssd1 vssd1 vccd1 vccd1 _18876_/D
+ sky130_fd_sc_hd__a22o_1
X_16035_ _18076_/Q vssd1 vssd1 vccd1 vccd1 _16035_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17319__S _17517_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10459_ _18549_/Q vssd1 vssd1 vccd1 vccd1 _10460_/C sky130_fd_sc_hd__inv_2
XFILLER_171_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20005__CLK _20091_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13178_ _13081_/A _13178_/A2 _13175_/Y _13199_/B vssd1 vssd1 vccd1 vccd1 _18909_/D
+ sky130_fd_sc_hd__a211oi_2
X_12129_ _19294_/Q _12094_/A _11926_/X _12096_/A vssd1 vssd1 vccd1 vccd1 _19294_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17911__S1 _19632_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18052__CLK _19851_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17986_ _19851_/CLK _17986_/D vssd1 vssd1 vccd1 vccd1 _17986_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19725_ _20050_/CLK _19725_/D repeater206/X vssd1 vssd1 vccd1 vccd1 _19725_/Q sky130_fd_sc_hd__dfrtp_1
X_16937_ _19481_/Q hold168/X _16946_/S vssd1 vssd1 vccd1 vccd1 _16937_/X sky130_fd_sc_hd__mux2_1
XFILLER_65_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11891__A _11891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17054__S _17524_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19656_ _19668_/CLK _19656_/D repeater270/X vssd1 vssd1 vccd1 vccd1 _19656_/Q sky130_fd_sc_hd__dfrtp_1
X_16868_ _16867_/X _11305_/Y _17547_/S vssd1 vssd1 vccd1 vccd1 _16868_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_237_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18607_ _19041_/CLK _18607_/D repeater263/X vssd1 vssd1 vccd1 vccd1 _18607_/Q sky130_fd_sc_hd__dfrtp_1
X_15819_ _17961_/Q vssd1 vssd1 vccd1 vccd1 _15819_/Y sky130_fd_sc_hd__inv_2
X_19587_ _19610_/CLK _19587_/D hold346/X vssd1 vssd1 vccd1 vccd1 _19587_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__16893__S _17487_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16799_ _16718_/Y _19291_/Q _17541_/S vssd1 vssd1 vccd1 vccd1 _16799_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09340_ _10186_/A _09340_/B _15749_/C vssd1 vssd1 vccd1 vccd1 _09342_/S sky130_fd_sc_hd__or3_1
XFILLER_240_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18538_ _19825_/CLK _18538_/D repeater229/X vssd1 vssd1 vccd1 vccd1 _18538_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_179_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12813__B1 _19247_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16004__B1 _17485_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09271_ _09271_/A vssd1 vssd1 vccd1 vccd1 _09271_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_61_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18469_ _18959_/CLK _18469_/D vssd1 vssd1 vccd1 vccd1 _18469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14566__B1 _14513_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10954__B _10954_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16641__B _16641_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17229__S _17524_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_86_HCLK clkbuf_4_13_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20115_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_87_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17902__S1 _19632_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08986_ _08986_/A vssd1 vssd1 vccd1 vccd1 _08986_/Y sky130_fd_sc_hd__inv_2
XFILLER_229_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09607_ _09607_/A vssd1 vssd1 vccd1 vccd1 _09607_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_56_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09538_ _19320_/Q vssd1 vssd1 vccd1 vccd1 _09538_/Y sky130_fd_sc_hd__inv_2
XPHY_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19940__CLK _19976_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09469_ _09469_/A _09469_/B vssd1 vssd1 vccd1 vccd1 _09612_/A sky130_fd_sc_hd__or2_1
XPHY_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11500_ _11500_/A vssd1 vssd1 vccd1 vccd1 _11500_/Y sky130_fd_sc_hd__inv_2
XPHY_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12480_ _19099_/Q _12478_/X _12299_/X _12479_/X vssd1 vssd1 vccd1 vccd1 _19099_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_185_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13240__B _13252_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11431_ _11579_/A _19146_/Q _11560_/C _19155_/Q vssd1 vssd1 vccd1 vccd1 _11431_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_22_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14309__B1 _13674_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14150_ _18672_/Q _13927_/A _14148_/A _14112_/X vssd1 vssd1 vccd1 vccd1 _18672_/D
+ sky130_fd_sc_hd__o211a_1
X_11362_ _11362_/A _11362_/B _11362_/C _11362_/D vssd1 vssd1 vccd1 vccd1 _11523_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_137_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16551__B _16622_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11791__B1 _09025_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13101_ _19185_/Q vssd1 vssd1 vccd1 vccd1 _13101_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17139__S _17493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10313_ _15578_/B vssd1 vssd1 vccd1 vccd1 _10314_/B sky130_fd_sc_hd__inv_2
XFILLER_153_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14081_ _19064_/Q vssd1 vssd1 vccd1 vccd1 _14081_/Y sky130_fd_sc_hd__inv_2
XFILLER_180_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11293_ _19587_/Q vssd1 vssd1 vccd1 vccd1 _11468_/B sky130_fd_sc_hd__inv_2
X_13032_ _18914_/Q vssd1 vssd1 vccd1 vccd1 _13086_/A sky130_fd_sc_hd__inv_2
XFILLER_98_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10244_ _10242_/Y _10243_/Y _19841_/Q _19668_/Q vssd1 vssd1 vccd1 vccd1 _10244_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_152_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16978__S _17548_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17840_ _16398_/Y _16399_/Y _16400_/Y _16401_/Y _17913_/S0 _19632_/Q vssd1 vssd1
+ vccd1 vccd1 _17840_/X sky130_fd_sc_hd__mux4_2
X_10175_ _10175_/A vssd1 vssd1 vccd1 vccd1 _10175_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_248_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17771_ _18387_/Q _18379_/Q _18371_/Q _18363_/Q _17923_/S0 _19646_/Q vssd1 vssd1
+ vccd1 vccd1 _17771_/X sky130_fd_sc_hd__mux4_2
X_14983_ hold245/X vssd1 vssd1 vccd1 vccd1 hold244/A sky130_fd_sc_hd__buf_2
XFILLER_59_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19510_ _19510_/CLK hold217/X repeater256/X vssd1 vssd1 vccd1 vccd1 _19510_/Q sky130_fd_sc_hd__dfrtp_1
X_16722_ _19468_/Q _16723_/B vssd1 vssd1 vccd1 vccd1 _16722_/Y sky130_fd_sc_hd__nand2_1
X_13934_ _13910_/A _13821_/B _13932_/Y _13927_/X vssd1 vssd1 vccd1 vccd1 _18722_/D
+ sky130_fd_sc_hd__a211oi_4
XFILLER_19_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19441_ _20064_/CLK _19441_/D repeater193/X vssd1 vssd1 vccd1 vccd1 _19441_/Q sky130_fd_sc_hd__dfrtp_1
X_16653_ _16964_/X _16555_/X _16992_/X _16556_/X vssd1 vssd1 vccd1 vccd1 _16656_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA_repeater191_A repeater210/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13865_ _19224_/Q _13834_/Y _19216_/Q _13912_/C vssd1 vssd1 vccd1 vccd1 _13865_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__17602__S _17605_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15604_ _18595_/Q vssd1 vssd1 vccd1 vccd1 _15606_/A sky130_fd_sc_hd__inv_2
X_12816_ _19236_/Q vssd1 vssd1 vccd1 vccd1 _12816_/Y sky130_fd_sc_hd__inv_2
X_19372_ _19971_/CLK _19372_/D repeater241/X vssd1 vssd1 vccd1 vccd1 _19372_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14796__B1 hold263/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16584_ _16616_/A vssd1 vssd1 vccd1 vccd1 _16615_/B sky130_fd_sc_hd__buf_4
X_13796_ _18716_/Q vssd1 vssd1 vccd1 vccd1 _13909_/D sky130_fd_sc_hd__inv_2
X_18323_ _18431_/CLK _18323_/D vssd1 vssd1 vccd1 vccd1 _18323_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15535_ _15535_/A _15535_/B vssd1 vssd1 vccd1 vccd1 _15535_/Y sky130_fd_sc_hd__nor2_1
X_12747_ _18818_/Q vssd1 vssd1 vccd1 vccd1 _13541_/A sky130_fd_sc_hd__inv_1
XFILLER_15_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_179_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10282__B1 _12058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18254_ _20077_/CLK _18254_/D vssd1 vssd1 vccd1 vccd1 _18254_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12678_ _12678_/A vssd1 vssd1 vccd1 vccd1 _12678_/X sky130_fd_sc_hd__buf_1
X_15466_ _15466_/A vssd1 vssd1 vccd1 vccd1 _15471_/B sky130_fd_sc_hd__inv_2
XFILLER_187_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17205_ _17204_/X _09480_/A _17482_/S vssd1 vssd1 vccd1 vccd1 _17205_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14417_ hold331/X vssd1 vssd1 vccd1 vccd1 _14417_/X sky130_fd_sc_hd__buf_2
X_11629_ _11629_/A vssd1 vssd1 vccd1 vccd1 _11629_/Y sky130_fd_sc_hd__inv_2
X_18185_ _18198_/CLK _18185_/D vssd1 vssd1 vccd1 vccd1 _18185_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15397_ _18531_/Q _13218_/B _13219_/B vssd1 vssd1 vccd1 vccd1 _15397_/X sky130_fd_sc_hd__a21bo_1
XFILLER_8_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17136_ _17473_/A0 _16525_/Y _17512_/S vssd1 vssd1 vccd1 vccd1 _17136_/X sky130_fd_sc_hd__mux2_1
X_14348_ _14450_/A _14545_/B _14557_/C vssd1 vssd1 vccd1 vccd1 _14352_/A sky130_fd_sc_hd__or3_4
XFILLER_156_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17049__S _17546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17067_ _16620_/Y _19386_/Q _17529_/S vssd1 vssd1 vccd1 vccd1 _17067_/X sky130_fd_sc_hd__mux2_1
X_14279_ _14279_/A vssd1 vssd1 vccd1 vccd1 _14279_/X sky130_fd_sc_hd__buf_2
XANTENNA__18669__SET_B repeater222/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16018_ _18348_/Q vssd1 vssd1 vccd1 vccd1 _16018_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14720__B1 _14600_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16888__S _17474_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17896__S0 _17908_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17969_ _20123_/CLK _17969_/D vssd1 vssd1 vccd1 vccd1 _17969_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_109_HCLK_A clkbuf_4_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19708_ _19720_/CLK _19708_/D repeater201/X vssd1 vssd1 vccd1 vccd1 _19708_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_214_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_238_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19639_ _19849_/CLK _19639_/D repeater257/X vssd1 vssd1 vccd1 vccd1 _19639_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__16776__A1 _09391_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_214_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17512__S _17512_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09323_ _09320_/Y _15722_/A _20044_/Q _09322_/A vssd1 vssd1 vccd1 vccd1 _09323_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14539__B1 _14509_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09254_ hold322/X vssd1 vssd1 vccd1 vccd1 _12313_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_21_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17820__S0 _17918_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_239_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09185_ _14713_/A vssd1 vssd1 vccd1 vccd1 _09185_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_147_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18098__CLK _18198_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11222__C1 _11221_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18819__RESET_B repeater231/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16798__S _17386_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17887__S0 _17908_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_248_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08969_ _08969_/A _08969_/B _08969_/C _08969_/D vssd1 vssd1 vccd1 vccd1 _08970_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_124_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11980_ _19372_/Q _11977_/X _11978_/X _11979_/X vssd1 vssd1 vccd1 vccd1 _19372_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_124_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11828__B2 _11801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_217_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10931_ _17727_/X _10923_/A _19674_/Q _10924_/A vssd1 vssd1 vccd1 vccd1 _19674_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_84_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17422__S _17544_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19607__RESET_B hold359/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10862_ _19705_/Q _10855_/X _10861_/X _10857_/X vssd1 vssd1 vccd1 vccd1 _19705_/D
+ sky130_fd_sc_hd__a22o_1
X_13650_ _16954_/X _13644_/X _18791_/Q _13646_/X vssd1 vssd1 vccd1 vccd1 _18791_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_72_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14242__A2 _14236_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_232_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16546__B _16583_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12601_ _19031_/Q _12598_/X _12599_/X _12600_/X vssd1 vssd1 vccd1 vccd1 _19031_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_31_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13581_ _18823_/Q _13580_/Y _13574_/X _13547_/B vssd1 vssd1 vccd1 vccd1 _18823_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_169_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10793_ _19737_/Q _10793_/B vssd1 vssd1 vccd1 vccd1 _19737_/D sky130_fd_sc_hd__and2_1
XFILLER_197_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19260__RESET_B repeater241/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15320_ _15320_/A vssd1 vssd1 vccd1 vccd1 _15320_/Y sky130_fd_sc_hd__inv_2
X_12532_ hold326/X vssd1 vssd1 vccd1 vccd1 hold325/A sky130_fd_sc_hd__clkbuf_2
XFILLER_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17811__S0 _17918_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15251_ _19780_/Q vssd1 vssd1 vccd1 vccd1 _15268_/A sky130_fd_sc_hd__inv_2
X_12463_ _19110_/Q _12457_/X _12410_/X _12458_/X vssd1 vssd1 vccd1 vccd1 _19110_/D
+ sky130_fd_sc_hd__a22o_1
X_11414_ _19565_/Q vssd1 vssd1 vccd1 vccd1 _11578_/A sky130_fd_sc_hd__inv_2
X_14202_ _14199_/Y _18698_/Q _19122_/Q _14031_/A _14201_/X vssd1 vssd1 vccd1 vccd1
+ _14219_/C sky130_fd_sc_hd__o221a_1
XFILLER_126_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15182_ _15744_/B _18488_/Q vssd1 vssd1 vccd1 vccd1 _15182_/X sky130_fd_sc_hd__or2_1
XFILLER_137_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12394_ hold306/X vssd1 vssd1 vccd1 vccd1 _12394_/X sky130_fd_sc_hd__buf_2
X_14133_ _18683_/Q _14135_/A _14116_/X _14133_/C1 vssd1 vssd1 vccd1 vccd1 _18683_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__08999__B _11936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11345_ _11480_/A _18982_/Q _11480_/A _18982_/Q vssd1 vssd1 vccd1 vccd1 _11345_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_19990_ _19992_/CLK _19990_/D repeater192/X vssd1 vssd1 vccd1 vccd1 _19990_/Q sky130_fd_sc_hd__dfrtp_1
X_14064_ _14064_/A _14064_/B _14059_/X _14063_/X vssd1 vssd1 vccd1 vccd1 _14094_/B
+ sky130_fd_sc_hd__or4bb_4
X_18941_ _18947_/CLK _18941_/D repeater213/X vssd1 vssd1 vccd1 vccd1 _18941_/Q sky130_fd_sc_hd__dfrtp_1
X_11276_ _19016_/Q vssd1 vssd1 vccd1 vccd1 _16665_/A sky130_fd_sc_hd__inv_2
XFILLER_140_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12314__B _12316_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13015_ _18926_/Q _13014_/Y _13006_/B _12980_/X vssd1 vssd1 vccd1 vccd1 _18926_/D
+ sky130_fd_sc_hd__o211a_1
X_10227_ _19829_/Q vssd1 vssd1 vccd1 vccd1 _10227_/Y sky130_fd_sc_hd__inv_2
X_18872_ _20049_/CLK _18872_/D repeater208/X vssd1 vssd1 vccd1 vccd1 _18872_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17878__S0 _17908_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_repeater204_A repeater205/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18860__CLK _18866_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08932__B2 _08928_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17823_ _17932_/Q _18454_/Q _18462_/Q _18062_/Q _17918_/S0 _18750_/Q vssd1 vssd1
+ vccd1 vccd1 _17823_/X sky130_fd_sc_hd__mux4_2
XANTENNA__19986__CLK _19992_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10158_ _19894_/Q _10154_/X _09086_/X _10156_/X vssd1 vssd1 vccd1 vccd1 _19894_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_208_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17754_ _17755_/S _11093_/Y _17754_/S vssd1 vssd1 vccd1 vccd1 _17754_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10089_ _19917_/Q _10088_/Y _10026_/A _10034_/B vssd1 vssd1 vccd1 vccd1 _19917_/D
+ sky130_fd_sc_hd__o211a_1
X_14966_ _14966_/A vssd1 vssd1 vccd1 vccd1 _14966_/X sky130_fd_sc_hd__clkbuf_2
X_16705_ _16682_/X _16705_/B _16705_/C vssd1 vssd1 vccd1 vccd1 _16705_/Y sky130_fd_sc_hd__nand3b_4
XFILLER_81_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13917_ _13917_/A vssd1 vssd1 vccd1 vccd1 _13917_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17685_ _15492_/X _19450_/Q _17696_/S vssd1 vssd1 vccd1 vccd1 _18567_/D sky130_fd_sc_hd__mux2_1
XFILLER_63_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14897_ _14897_/A vssd1 vssd1 vccd1 vccd1 _14898_/A sky130_fd_sc_hd__inv_2
X_19424_ _19997_/CLK _19424_/D repeater271/X vssd1 vssd1 vccd1 vccd1 _19424_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17332__S _17488_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19348__RESET_B repeater245/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16636_ _16812_/X _16573_/X _16875_/X _16574_/X _16635_/X vssd1 vssd1 vccd1 vccd1
+ _16641_/B sky130_fd_sc_hd__o221a_4
XANTENNA__14769__B1 _14693_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13848_ _13844_/Y _18720_/Q _13845_/Y _18714_/Q _13847_/X vssd1 vssd1 vccd1 vccd1
+ _13850_/C sky130_fd_sc_hd__a221o_1
XFILLER_35_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_222_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19355_ _19968_/CLK _19355_/D hold370/X vssd1 vssd1 vccd1 vccd1 _19355_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_222_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16567_ _17146_/X _16512_/X _17129_/X _16513_/X _16566_/X vssd1 vssd1 vccd1 vccd1
+ _16567_/X sky130_fd_sc_hd__o221a_4
X_13779_ _18733_/Q vssd1 vssd1 vccd1 vccd1 _13831_/A sky130_fd_sc_hd__inv_2
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18306_ _18435_/CLK _18306_/D vssd1 vssd1 vccd1 vccd1 _18306_/Q sky130_fd_sc_hd__dfxtp_1
X_15518_ _18573_/Q _18574_/Q _15518_/C vssd1 vssd1 vccd1 vccd1 _15523_/B sky130_fd_sc_hd__or3_1
XFILLER_200_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17802__S0 _17918_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19286_ _19288_/CLK _19286_/D repeater211/X vssd1 vssd1 vccd1 vccd1 _19286_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_149_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16498_ _17208_/X _15898_/X _17214_/X _15889_/X _16497_/X vssd1 vssd1 vccd1 vccd1
+ _16498_/X sky130_fd_sc_hd__o221a_2
X_18237_ _18268_/CLK _18237_/D vssd1 vssd1 vccd1 vccd1 _18237_/Q sky130_fd_sc_hd__dfxtp_1
X_15449_ _18556_/Q vssd1 vssd1 vccd1 vccd1 _15450_/B sky130_fd_sc_hd__inv_2
XFILLER_191_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16930__A1 hold206/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16391__C1 _16390_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18168_ _18169_/CLK _18168_/D vssd1 vssd1 vccd1 vccd1 _18168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_190_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17119_ _17473_/A0 _16534_/Y _17512_/S vssd1 vssd1 vccd1 vccd1 _17119_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18912__RESET_B repeater188/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18099_ _18260_/CLK _18099_/D vssd1 vssd1 vccd1 vccd1 _18099_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09086__A _10448_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09941_ _09854_/A _19337_/Q _09863_/A _19347_/Q _09940_/X vssd1 vssd1 vccd1 vccd1
+ _09947_/C sky130_fd_sc_hd__o221a_1
XANTENNA__17507__S _17567_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20061_ _20064_/CLK _20061_/D repeater200/X vssd1 vssd1 vccd1 vccd1 _20061_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17869__S0 _18760_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09872_ _09872_/A _09960_/A vssd1 vssd1 vccd1 vccd1 _09873_/B sky130_fd_sc_hd__or2_2
XFILLER_97_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrepeater220 repeater223/X vssd1 vssd1 vccd1 vccd1 repeater220/X sky130_fd_sc_hd__buf_4
Xrepeater231 repeater232/X vssd1 vssd1 vccd1 vccd1 repeater231/X sky130_fd_sc_hd__buf_8
Xrepeater242 repeater243/X vssd1 vssd1 vccd1 vccd1 repeater242/X sky130_fd_sc_hd__buf_8
XANTENNA__12240__A hold322/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater253 hold365/A vssd1 vssd1 vccd1 vccd1 repeater253/X sky130_fd_sc_hd__buf_8
Xrepeater264 repeater265/X vssd1 vssd1 vccd1 vccd1 repeater264/X sky130_fd_sc_hd__buf_6
XPHY_4407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_116_HCLK clkbuf_opt_0_HCLK/A vssd1 vssd1 vccd1 vccd1 _19608_/CLK sky130_fd_sc_hd__clkbuf_16
Xrepeater275 hold363/A vssd1 vssd1 vccd1 vccd1 hold348/A sky130_fd_sc_hd__buf_8
Xrepeater286 input34/X vssd1 vssd1 vccd1 vccd1 hold354/A sky130_fd_sc_hd__buf_8
XPHY_4418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17242__S _17490_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_214_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_241_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14167__A _19114_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09306_ _18660_/Q _09305_/B _09305_/Y vssd1 vssd1 vccd1 vccd1 _15727_/A sky130_fd_sc_hd__o21ai_1
XFILLER_194_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17174__A1 _12948_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09237_ _15709_/A _09226_/X _18646_/Q _18647_/Q vssd1 vssd1 vccd1 vccd1 _09238_/B
+ sky130_fd_sc_hd__a31oi_1
XFILLER_186_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15185__B1 _10448_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09168_ _14699_/A vssd1 vssd1 vccd1 vccd1 _09168_/X sky130_fd_sc_hd__clkbuf_2
X_09099_ _20094_/Q _09084_/X _09098_/X _09087_/X vssd1 vssd1 vccd1 vccd1 _20094_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_134_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11130_ _11123_/A _11064_/B _17747_/X _19631_/Q vssd1 vssd1 vccd1 vccd1 _19631_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_162_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17417__S _17536_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11061_ _19633_/Q vssd1 vssd1 vccd1 vccd1 _11061_/X sky130_fd_sc_hd__buf_1
XFILLER_103_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10012_ _19912_/Q vssd1 vssd1 vccd1 vccd1 _10084_/A sky130_fd_sc_hd__inv_2
XFILLER_130_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14820_ _14821_/A vssd1 vssd1 vccd1 vccd1 _14820_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__14999__B1 _14998_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14751_ _14751_/A vssd1 vssd1 vccd1 vccd1 _14751_/X sky130_fd_sc_hd__buf_2
XFILLER_205_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11963_ _11979_/A vssd1 vssd1 vccd1 vccd1 _11963_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_leaf_155_HCLK_A clkbuf_4_1_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17152__S _17536_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13702_ _13700_/A _14641_/B _13700_/Y vssd1 vssd1 vccd1 vccd1 _18762_/D sky130_fd_sc_hd__a21oi_1
XANTENNA__19441__RESET_B repeater193/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10914_ _10914_/A vssd1 vssd1 vccd1 vccd1 _10914_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19389__CLK _20091_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17470_ _17469_/X _10240_/Y _17566_/S vssd1 vssd1 vccd1 vccd1 _17470_/X sky130_fd_sc_hd__mux2_1
X_14682_ _14683_/A vssd1 vssd1 vccd1 vccd1 _14682_/X sky130_fd_sc_hd__clkbuf_2
X_11894_ _19421_/Q _11891_/X hold300/X _11892_/X vssd1 vssd1 vccd1 vccd1 _19421_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_205_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_204_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16421_ _18273_/Q vssd1 vssd1 vccd1 vccd1 _16421_/Y sky130_fd_sc_hd__inv_2
X_10845_ _10845_/A vssd1 vssd1 vccd1 vccd1 _10845_/X sky130_fd_sc_hd__buf_1
XANTENNA__12226__A1 _19235_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13633_ _18799_/Q _10196_/B _13630_/X _10196_/A _13632_/Y vssd1 vssd1 vccd1 vccd1
+ _13634_/A sky130_fd_sc_hd__o32a_1
XFILLER_204_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16991__S _17487_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19140_ _19582_/CLK _19140_/D hold348/A vssd1 vssd1 vccd1 vccd1 _19140_/Q sky130_fd_sc_hd__dfrtp_1
X_16352_ _18256_/Q vssd1 vssd1 vccd1 vccd1 _16352_/Y sky130_fd_sc_hd__inv_2
X_13564_ _18833_/Q _13563_/Y _13560_/X _13557_/B vssd1 vssd1 vccd1 vccd1 _18833_/D
+ sky130_fd_sc_hd__o211a_1
X_10776_ _17625_/X _10772_/X _19748_/Q _10774_/X vssd1 vssd1 vccd1 vccd1 _19748_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_185_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11985__B1 _11922_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12309__B _12316_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15303_ _18631_/Q _18633_/Q _18634_/Q _18630_/Q vssd1 vssd1 vccd1 vccd1 _15305_/C
+ sky130_fd_sc_hd__or4_4
XFILLER_40_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12515_ _19076_/Q _12512_/X _12344_/X _12513_/X vssd1 vssd1 vccd1 vccd1 _19076_/D
+ sky130_fd_sc_hd__a22o_1
X_19071_ _19610_/CLK _19071_/D hold361/X vssd1 vssd1 vccd1 vccd1 _19071_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__15176__B1 _10698_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13495_ _15319_/B _13495_/B vssd1 vssd1 vccd1 vccd1 _15320_/A sky130_fd_sc_hd__nand2_2
X_16283_ _18135_/Q vssd1 vssd1 vccd1 vccd1 _16283_/Y sky130_fd_sc_hd__inv_2
XANTENNA_repeater154_A _17413_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18022_ _18142_/CLK _18022_/D vssd1 vssd1 vccd1 vccd1 _18022_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12446_ _19123_/Q _12441_/X _12380_/X _12444_/X vssd1 vssd1 vccd1 vccd1 _19123_/D
+ sky130_fd_sc_hd__a22o_1
X_15234_ _18622_/D hold213/X vssd1 vssd1 vccd1 vccd1 hold212/A sky130_fd_sc_hd__or2_1
XFILLER_172_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12377_ _12428_/A vssd1 vssd1 vccd1 vccd1 _12402_/A sky130_fd_sc_hd__buf_2
X_15165_ _17948_/Q _15158_/X _14709_/A _15160_/X vssd1 vssd1 vccd1 vccd1 _17948_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_output83_A _16541_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14116_ _14116_/A vssd1 vssd1 vccd1 vccd1 _14116_/X sky130_fd_sc_hd__clkbuf_2
X_11328_ _18966_/Q vssd1 vssd1 vccd1 vccd1 _11328_/Y sky130_fd_sc_hd__inv_2
XFILLER_180_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15096_ _15096_/A vssd1 vssd1 vccd1 vccd1 _15097_/A sky130_fd_sc_hd__inv_2
X_19973_ _19984_/CLK _19973_/D repeater244/X vssd1 vssd1 vccd1 vccd1 _19973_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17327__S _17534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18924_ _19283_/CLK _18924_/D repeater212/X vssd1 vssd1 vccd1 vccd1 _18924_/Q sky130_fd_sc_hd__dfrtp_1
X_11259_ _19596_/Q vssd1 vssd1 vccd1 vccd1 _11476_/A sky130_fd_sc_hd__inv_2
X_14047_ _14043_/Y _18701_/Q _19068_/Q _14010_/A vssd1 vssd1 vccd1 vccd1 _14047_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_95_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12162__B1 _12030_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_139_HCLK clkbuf_4_3_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19841_/CLK sky130_fd_sc_hd__clkbuf_16
X_18855_ _18856_/CLK _18855_/D repeater231/X vssd1 vssd1 vccd1 vccd1 _18855_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_79_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19529__RESET_B repeater221/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17806_ _18187_/Q _18179_/Q _18171_/Q _18155_/Q _17918_/S0 _18750_/Q vssd1 vssd1
+ vccd1 vccd1 _17806_/X sky130_fd_sc_hd__mux4_1
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18786_ _19041_/CLK _18786_/D repeater263/X vssd1 vssd1 vccd1 vccd1 _18786_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_94_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15998_ _16509_/A vssd1 vssd1 vccd1 vccd1 _15998_/X sky130_fd_sc_hd__buf_1
XFILLER_243_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_236_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17737_ _15372_/X _19708_/Q _18508_/D vssd1 vssd1 vccd1 vccd1 _17737_/X sky130_fd_sc_hd__mux2_1
X_14949_ _20074_/Q vssd1 vssd1 vccd1 vccd1 _14949_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__13662__B1 _12032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16467__A _16467_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17062__S _17493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17668_ _15564_/Y _19467_/Q _17683_/S vssd1 vssd1 vccd1 vccd1 _18584_/D sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_14_HCLK_A clkbuf_4_2_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19407_ _19984_/CLK _19407_/D repeater243/X vssd1 vssd1 vccd1 vccd1 _19407_/Q sky130_fd_sc_hd__dfrtp_1
X_16619_ _16619_/A _16621_/B vssd1 vssd1 vccd1 vccd1 _16619_/Y sky130_fd_sc_hd__nor2_1
XFILLER_196_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_77_HCLK_A clkbuf_opt_4_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17599_ _15337_/X _19704_/Q _17600_/S vssd1 vssd1 vccd1 vccd1 _17599_/X sky130_fd_sc_hd__mux2_1
XANTENNA__20087__RESET_B repeater205/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_2_HCLK_A clkbuf_4_0_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19338_ _19352_/CLK _19338_/D repeater245/X vssd1 vssd1 vccd1 vccd1 _19338_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_188_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11976__B1 _11975_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19269_ _19283_/CLK _19269_/D repeater216/X vssd1 vssd1 vccd1 vccd1 _19269_/Q sky130_fd_sc_hd__dfrtp_4
X_09022_ _20121_/Q _09015_/X _09021_/X _09019_/X vssd1 vssd1 vccd1 vccd1 _20121_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13717__A1 _18760_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold200 HADDR[2] vssd1 vssd1 vccd1 vccd1 input23/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold211 HTRANS[1] vssd1 vssd1 vccd1 vccd1 input37/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold222 hold222/A vssd1 vssd1 vccd1 vccd1 hold222/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold233 hold233/A vssd1 vssd1 vccd1 vccd1 hold233/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold244 hold244/A vssd1 vssd1 vccd1 vccd1 hold244/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 hold369/X vssd1 vssd1 vccd1 vccd1 input75/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_160_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold266 input33/X vssd1 vssd1 vccd1 vccd1 hold266/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold277 input45/X vssd1 vssd1 vccd1 vccd1 hold277/X sky130_fd_sc_hd__dlygate4sd3_1
X_20113_ _20115_/CLK _20113_/D repeater238/X vssd1 vssd1 vccd1 vccd1 _20113_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__17237__S _17318_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold288 hold288/A vssd1 vssd1 vccd1 vccd1 hold288/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold299 HWDATA[22] vssd1 vssd1 vccd1 vccd1 input52/A sky130_fd_sc_hd__dlygate4sd3_1
X_09924_ _19341_/Q vssd1 vssd1 vccd1 vccd1 _09924_/Y sky130_fd_sc_hd__inv_2
XFILLER_120_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12153__B1 _12098_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19952__RESET_B repeater244/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20044_ _20066_/CLK _20044_/D repeater209/X vssd1 vssd1 vccd1 vccd1 _20044_/Q sky130_fd_sc_hd__dfrtp_1
X_09855_ _09855_/A _09992_/A vssd1 vssd1 vccd1 vccd1 _09856_/B sky130_fd_sc_hd__or2_2
XANTENNA__11900__B1 hold276/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18286__CLK _19847_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09786_ _09740_/A _09740_/B _09784_/Y _09813_/C vssd1 vssd1 vccd1 vccd1 _19984_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_100_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16096__B _16096_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_241_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12208__A1 _19247_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10630_ _19803_/Q _10606_/A _10613_/B _10609_/X vssd1 vssd1 vccd1 vccd1 _19803_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_201_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11967__B1 _09064_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10561_ _10561_/A _10576_/C vssd1 vssd1 vccd1 vccd1 _10595_/D sky130_fd_sc_hd__or2_1
XANTENNA__18834__RESET_B repeater239/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11431__A2 _19146_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12300_ _12300_/A vssd1 vssd1 vccd1 vccd1 _12300_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_13280_ _13280_/A _15909_/A vssd1 vssd1 vccd1 vccd1 _13654_/A sky130_fd_sc_hd__or2_1
X_10492_ _11655_/A _19540_/Q _10492_/C _19539_/Q vssd1 vssd1 vccd1 vccd1 _10493_/B
+ sky130_fd_sc_hd__or4b_4
XFILLER_212_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12231_ _19232_/Q _12228_/X _11981_/X _12229_/X vssd1 vssd1 vccd1 vccd1 _19232_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_30_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12162_ _19275_/Q _12157_/X _12030_/X _12158_/X vssd1 vssd1 vccd1 vccd1 _19275_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_135_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11113_ _19637_/Q _11113_/B vssd1 vssd1 vccd1 vccd1 _11113_/Y sky130_fd_sc_hd__nor2_1
XFILLER_123_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17147__S _17543_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12093_ _19316_/Q _12082_/X _12092_/X _12084_/X vssd1 vssd1 vccd1 vccd1 _19316_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_150_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16970_ _16969_/X _09684_/Y _17523_/S vssd1 vssd1 vccd1 vccd1 _16970_/X sky130_fd_sc_hd__mux2_1
XFILLER_123_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18629__CLK _19780_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19693__RESET_B repeater208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15921_ _18027_/Q vssd1 vssd1 vccd1 vccd1 _15921_/Y sky130_fd_sc_hd__inv_2
X_11044_ _11039_/A _10266_/B _10266_/A vssd1 vssd1 vccd1 vccd1 _11044_/X sky130_fd_sc_hd__o21a_1
XFILLER_89_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12695__A1 _18969_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18640_ _19780_/CLK _18640_/D repeater226/X vssd1 vssd1 vccd1 vccd1 _18640_/Q sky130_fd_sc_hd__dfrtp_1
X_15852_ _19765_/Q vssd1 vssd1 vccd1 vccd1 _15852_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14803_ _14803_/A vssd1 vssd1 vccd1 vccd1 _14804_/A sky130_fd_sc_hd__inv_2
XFILLER_64_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12447__A1 _19122_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18571_ _19462_/CLK _18571_/D repeater273/X vssd1 vssd1 vccd1 vccd1 _18571_/Q sky130_fd_sc_hd__dfrtp_1
X_15783_ _18018_/Q vssd1 vssd1 vccd1 vccd1 _15783_/Y sky130_fd_sc_hd__inv_2
XANTENNA_output121_A _16752_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12995_ _18934_/Q _12994_/Y _12877_/B _12980_/X vssd1 vssd1 vccd1 vccd1 _18934_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_92_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10458__B1 _10427_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17522_ _17521_/X _09904_/Y _17522_/S vssd1 vssd1 vccd1 vccd1 _17522_/X sky130_fd_sc_hd__mux2_1
X_14734_ _14734_/A vssd1 vssd1 vccd1 vccd1 _14734_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_233_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11946_ _19394_/Q _11939_/X _09025_/X _11942_/X vssd1 vssd1 vccd1 vccd1 _19394_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_55_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17453_ _17452_/X _12922_/Y _17487_/S vssd1 vssd1 vccd1 vccd1 _17453_/X sky130_fd_sc_hd__mux2_1
X_14665_ _18243_/Q _14657_/A _14567_/X _14658_/A vssd1 vssd1 vccd1 vccd1 _18243_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_repeater271_A repeater272/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_221_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11877_ _11915_/A vssd1 vssd1 vccd1 vccd1 _11892_/A sky130_fd_sc_hd__buf_2
XANTENNA__17610__S _17614_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16404_ _18041_/Q vssd1 vssd1 vccd1 vccd1 _16404_/Y sky130_fd_sc_hd__inv_2
XFILLER_232_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13616_ _18800_/Q _13616_/B vssd1 vssd1 vccd1 vccd1 _13617_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09076__B1 _09075_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10828_ _19700_/Q vssd1 vssd1 vccd1 vccd1 _15349_/A sky130_fd_sc_hd__clkbuf_2
X_17384_ _17383_/X _20008_/Q _17414_/S vssd1 vssd1 vccd1 vccd1 _17384_/X sky130_fd_sc_hd__mux2_2
X_14596_ _18283_/Q _14588_/A _14567_/X _14589_/A vssd1 vssd1 vccd1 vccd1 _18283_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11958__B1 hold300/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_186_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19123_ _19609_/CLK _19123_/D hold355/X vssd1 vssd1 vccd1 vccd1 _19123_/Q sky130_fd_sc_hd__dfrtp_2
X_16335_ _18056_/Q vssd1 vssd1 vccd1 vccd1 _16335_/Y sky130_fd_sc_hd__inv_2
X_13547_ _13547_/A _13547_/B vssd1 vssd1 vccd1 vccd1 _13577_/A sky130_fd_sc_hd__or2_1
XFILLER_185_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18652__D hold341/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10759_ _19872_/Q _10759_/B _10759_/C vssd1 vssd1 vccd1 vccd1 _10765_/B sky130_fd_sc_hd__or3_1
XFILLER_187_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16897__A0 _17473_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19054_ _19577_/CLK _19054_/D repeater267/X vssd1 vssd1 vccd1 vccd1 _19054_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18504__RESET_B repeater222/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16266_ _18471_/Q vssd1 vssd1 vccd1 vccd1 _16266_/Y sky130_fd_sc_hd__inv_2
X_13478_ _13466_/A _13466_/B _13476_/Y _13437_/X vssd1 vssd1 vccd1 vccd1 _18843_/D
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__18159__CLK _18198_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18005_ _18416_/CLK _18005_/D vssd1 vssd1 vccd1 vccd1 _18005_/Q sky130_fd_sc_hd__dfxtp_1
X_15217_ _15217_/A vssd1 vssd1 vccd1 vccd1 _15217_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19404__CLK _19984_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12429_ _19132_/Q _12427_/X _12299_/X _12428_/X vssd1 vssd1 vccd1 vccd1 _19132_/D
+ sky130_fd_sc_hd__a22o_1
X_16197_ _16043_/Y _16196_/Y _18747_/Q vssd1 vssd1 vccd1 vccd1 _16197_/X sky130_fd_sc_hd__o21a_1
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12383__B1 _12382_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15148_ _15148_/A vssd1 vssd1 vccd1 vccd1 _15148_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_126_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17057__S _17547_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15079_ _18004_/Q _15072_/A hold263/X _15073_/A vssd1 vssd1 vccd1 vccd1 _18004_/D
+ sky130_fd_sc_hd__a22o_1
X_19956_ _19956_/CLK _19956_/D repeater245/X vssd1 vssd1 vccd1 vccd1 _19956_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_206_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18907_ _18908_/CLK _18907_/D repeater188/X vssd1 vssd1 vccd1 vccd1 _18907_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__16896__S _17474_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19887_ _20051_/CLK _19887_/D repeater200/X vssd1 vssd1 vccd1 vccd1 _19887_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_206_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09640_ _09640_/A vssd1 vssd1 vccd1 vccd1 _09807_/A sky130_fd_sc_hd__clkbuf_2
X_18838_ _20107_/CLK _18838_/D repeater234/X vssd1 vssd1 vccd1 vccd1 _18838_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_110_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09571_ _09571_/A vssd1 vssd1 vccd1 vccd1 _09571_/Y sky130_fd_sc_hd__inv_2
XFILLER_215_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12438__A1 _19125_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18769_ _20058_/CLK _18769_/D repeater194/X vssd1 vssd1 vccd1 vccd1 _18769_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_222_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10449__B1 _10448_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17377__A1 _17864_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11134__A _12053_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17520__S _17548_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16644__B _16647_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12610__A1 _19024_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10692__B _10718_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09005_ _19500_/Q _19499_/Q _11842_/D vssd1 vssd1 vccd1 vccd1 _10430_/A sky130_fd_sc_hd__or3_4
XFILLER_247_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_183_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_hold197_A HADDR[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12126__B1 _11920_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09907_ _19939_/Q _09904_/Y _09866_/A _19350_/Q _09906_/X vssd1 vssd1 vccd1 vccd1
+ _09911_/C sky130_fd_sc_hd__o221a_1
XFILLER_116_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20027_ _20115_/CLK _20027_/D repeater239/X vssd1 vssd1 vccd1 vccd1 _20027_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_247_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09838_ _19948_/Q vssd1 vssd1 vccd1 vccd1 _09857_/B sky130_fd_sc_hd__inv_2
XANTENNA__16812__A0 _16811_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19033__RESET_B repeater267/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12429__A1 _19132_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09769_ _09769_/A vssd1 vssd1 vccd1 vccd1 _09769_/Y sky130_fd_sc_hd__inv_2
XFILLER_132_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11800_ _11800_/A vssd1 vssd1 vccd1 vccd1 _11800_/X sky130_fd_sc_hd__buf_1
XPHY_4034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12780_ _19247_/Q vssd1 vssd1 vccd1 vccd1 _16619_/A sky130_fd_sc_hd__inv_2
XFILLER_27_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_203_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrebuffer70 _09729_/A vssd1 vssd1 vccd1 vccd1 _09767_/A sky130_fd_sc_hd__dlygate4sd1_1
XPHY_4067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer81 _13538_/B vssd1 vssd1 vccd1 vccd1 _13594_/A sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_14_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11731_ _11731_/A vssd1 vssd1 vccd1 vccd1 _11731_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_70_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrebuffer92 _13068_/B vssd1 vssd1 vccd1 vccd1 _13205_/C1 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_4089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16576__C1 _16575_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17430__S _17565_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10860__B1 _10451_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14450_ _14450_/A _14450_/B _14557_/C vssd1 vssd1 vccd1 vccd1 _14452_/A sky130_fd_sc_hd__or3_4
X_11662_ _10531_/X _11660_/Y _11661_/Y vssd1 vssd1 vccd1 vccd1 _11674_/A sky130_fd_sc_hd__o21ai_2
XPHY_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_60_HCLK_A clkbuf_4_12_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14051__B1 _19081_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13401_ _13397_/Y _18840_/Q _13398_/Y _18838_/Q _13400_/X vssd1 vssd1 vccd1 vccd1
+ _13402_/D sky130_fd_sc_hd__o221a_1
XFILLER_168_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10613_ _10613_/A _10613_/B _10613_/C _10584_/C vssd1 vssd1 vccd1 vccd1 _10933_/B
+ sky130_fd_sc_hd__or4b_4
XANTENNA__11979__A _11979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11593_ _19574_/Q _11591_/X _11592_/X _11586_/A vssd1 vssd1 vccd1 vccd1 _19574_/D
+ sky130_fd_sc_hd__o211a_1
X_14381_ _14381_/A vssd1 vssd1 vccd1 vccd1 _14382_/A sky130_fd_sc_hd__inv_2
XPHY_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14355__A hold237/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16879__A0 _15963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16120_ _19404_/Q vssd1 vssd1 vccd1 vccd1 _16120_/Y sky130_fd_sc_hd__inv_2
X_10544_ _19804_/Q _19803_/Q _10577_/B vssd1 vssd1 vccd1 vccd1 _10561_/A sky130_fd_sc_hd__or3_1
X_13332_ _18847_/Q vssd1 vssd1 vccd1 vccd1 _13470_/A sky130_fd_sc_hd__inv_2
XPHY_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16051_ _19687_/Q vssd1 vssd1 vccd1 vccd1 _16051_/Y sky130_fd_sc_hd__inv_2
X_10475_ _17699_/X _10471_/X _19820_/Q _10472_/X vssd1 vssd1 vccd1 vccd1 _19820_/D
+ sky130_fd_sc_hd__a22o_1
X_13263_ _13256_/X _13262_/B _15082_/A _18756_/Q _13737_/B vssd1 vssd1 vccd1 vccd1
+ _13263_/X sky130_fd_sc_hd__a32o_1
XANTENNA__12365__B1 _12232_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15002_ _18955_/Q vssd1 vssd1 vccd1 vccd1 _15002_/X sky130_fd_sc_hd__buf_2
X_12214_ _19243_/Q _12212_/X _12107_/X _12213_/X vssd1 vssd1 vccd1 vccd1 _19243_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_124_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13194_ _18900_/Q _13193_/Y _13180_/X _13194_/C1 vssd1 vssd1 vccd1 vccd1 _18900_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_136_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19803__RESET_B repeater222/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19810_ _19810_/CLK _19810_/D repeater224/X vssd1 vssd1 vccd1 vccd1 _19810_/Q sky130_fd_sc_hd__dfrtp_1
X_12145_ _19288_/Q _12143_/X _12083_/X _12144_/X vssd1 vssd1 vccd1 vccd1 _19288_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_150_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12117__B1 _12038_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16953_ _17779_/X _18791_/Q _16957_/S vssd1 vssd1 vccd1 vccd1 _16953_/X sky130_fd_sc_hd__mux2_1
X_12076_ hold289/X vssd1 vssd1 vccd1 vccd1 _12076_/X sky130_fd_sc_hd__buf_2
X_19741_ _20051_/CLK _19741_/D repeater200/X vssd1 vssd1 vccd1 vccd1 _19741_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_173_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11027_ _15296_/A _11027_/B vssd1 vssd1 vccd1 vccd1 _15294_/A sky130_fd_sc_hd__or2_1
XFILLER_77_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15904_ _15904_/A vssd1 vssd1 vccd1 vccd1 _15904_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__17605__S _17605_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19672_ _19812_/CLK _19672_/D repeater225/X vssd1 vssd1 vccd1 vccd1 _19672_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA__15914__A _15914_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16884_ _16883_/X _09879_/Y _17524_/S vssd1 vssd1 vccd1 vccd1 _16884_/X sky130_fd_sc_hd__mux2_1
X_18623_ _18623_/CLK _18623_/D hold351/X vssd1 vssd1 vccd1 vccd1 _18623_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_64_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15835_ _15971_/A vssd1 vssd1 vccd1 vccd1 _15836_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_46_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18554_ _18633_/CLK _18554_/D repeater224/X vssd1 vssd1 vccd1 vccd1 _18554_/Q sky130_fd_sc_hd__dfrtp_1
X_15766_ _15764_/Y _18523_/Q _11655_/X _15765_/X vssd1 vssd1 vccd1 vccd1 _18520_/D
+ sky130_fd_sc_hd__a31o_1
XANTENNA__09297__B1 _09101_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12978_ _12978_/A vssd1 vssd1 vccd1 vccd1 _12978_/Y sky130_fd_sc_hd__inv_2
XFILLER_233_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17505_ _17504_/X _15935_/Y _17565_/S vssd1 vssd1 vccd1 vccd1 _17505_/X sky130_fd_sc_hd__mux2_1
X_14717_ _14718_/A vssd1 vssd1 vccd1 vccd1 _14717_/X sky130_fd_sc_hd__clkbuf_2
X_18485_ _19545_/CLK _18485_/D repeater225/X vssd1 vssd1 vccd1 vccd1 _18485_/Q sky130_fd_sc_hd__dfrtp_1
X_11929_ _11841_/X _19400_/Q _11929_/S vssd1 vssd1 vccd1 vccd1 _19400_/D sky130_fd_sc_hd__mux2_1
XFILLER_17_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18756__RESET_B repeater195/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15697_ _15697_/A vssd1 vssd1 vccd1 vccd1 _15697_/Y sky130_fd_sc_hd__inv_2
XPHY_4590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17340__S _19498_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10851__B1 _10423_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17436_ _17435_/X _10227_/Y _17566_/S vssd1 vssd1 vccd1 vccd1 _17436_/X sky130_fd_sc_hd__mux2_1
X_14648_ _18255_/Q _14643_/X _09174_/X _14645_/X vssd1 vssd1 vccd1 vccd1 _18255_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_221_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17367_ _17366_/X _11311_/Y _17459_/S vssd1 vssd1 vccd1 vccd1 _17367_/X sky130_fd_sc_hd__mux2_1
X_14579_ _18294_/Q _14572_/X _14578_/X _14574_/X vssd1 vssd1 vccd1 vccd1 _18294_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_119_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19106_ _19109_/CLK _19106_/D hold361/X vssd1 vssd1 vccd1 vccd1 _19106_/Q sky130_fd_sc_hd__dfrtp_1
X_16318_ _16314_/Y _15971_/X _16315_/Y _15838_/X _16317_/X vssd1 vssd1 vccd1 vccd1
+ _16318_/X sky130_fd_sc_hd__o221a_1
XANTENNA__17531__A1 _13483_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17298_ _17297_/X _15487_/A _17524_/S vssd1 vssd1 vccd1 vccd1 _17298_/X sky130_fd_sc_hd__mux2_1
XFILLER_173_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19037_ _19041_/CLK _19037_/D repeater266/X vssd1 vssd1 vccd1 vccd1 _19037_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_134_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16249_ _11742_/A _16243_/X _16246_/Y _16248_/X vssd1 vssd1 vccd1 vccd1 _16249_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_115_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput102 _16735_/Y vssd1 vssd1 vccd1 vccd1 HRDATA[30] sky130_fd_sc_hd__clkbuf_2
Xoutput113 _15780_/X vssd1 vssd1 vccd1 vccd1 IRQ[10] sky130_fd_sc_hd__clkbuf_2
XFILLER_133_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput124 _15775_/X vssd1 vssd1 vccd1 vccd1 IRQ[6] sky130_fd_sc_hd__clkbuf_2
Xoutput135 _15732_/Y vssd1 vssd1 vccd1 vccd1 SSn_S3 sky130_fd_sc_hd__clkbuf_2
XANTENNA__19544__RESET_B repeater221/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09094__A _12232_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19939_ _19976_/CLK _19939_/D hold371/X vssd1 vssd1 vccd1 vccd1 _19939_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_229_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09524__B2 _19313_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17515__S _17548_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_229_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09623_ _20002_/Q vssd1 vssd1 vccd1 vccd1 _09668_/A sky130_fd_sc_hd__inv_2
XFILLER_228_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09554_ _09485_/A _19315_/Q _09474_/B _19303_/Q _09553_/X vssd1 vssd1 vccd1 vccd1
+ _09564_/B sky130_fd_sc_hd__o221a_1
XANTENNA__09288__B1 _09077_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14281__B1 _13674_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18497__RESET_B repeater203/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09485_ _09485_/A _09584_/A vssd1 vssd1 vccd1 vccd1 _09486_/B sky130_fd_sc_hd__or2_2
XPHY_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17250__S _17542_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12595__B1 hold259/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09269__A _09270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16325__A2 _16148_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12347__B1 hold281/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10260_ _19873_/Q vssd1 vssd1 vccd1 vccd1 _12058_/A sky130_fd_sc_hd__inv_2
XFILLER_3_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10191_ _18799_/Q vssd1 vssd1 vccd1 vccd1 _10196_/A sky130_fd_sc_hd__inv_2
XFILLER_78_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17425__S _17459_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13950_ _13950_/A _13954_/A vssd1 vssd1 vccd1 vccd1 _13951_/B sky130_fd_sc_hd__or2_2
XFILLER_120_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12901_ _19262_/Q vssd1 vssd1 vccd1 vccd1 _12901_/Y sky130_fd_sc_hd__inv_2
X_13881_ _13878_/Y _18721_/Q _13879_/Y _18716_/Q _13880_/X vssd1 vssd1 vccd1 vccd1
+ _13882_/D sky130_fd_sc_hd__o221a_1
XFILLER_219_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15620_ _18599_/Q vssd1 vssd1 vccd1 vccd1 _15622_/A sky130_fd_sc_hd__inv_2
XANTENNA__13254__A _18870_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12832_ _12827_/Y _18805_/Q _19243_/Q _13543_/A _12831_/X vssd1 vssd1 vccd1 vccd1
+ _12833_/D sky130_fd_sc_hd__o221a_1
XANTENNA__09279__B1 _09108_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_215_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15551_ _15555_/B vssd1 vssd1 vccd1 vccd1 _15557_/B sky130_fd_sc_hd__inv_2
X_12763_ _19240_/Q _18817_/Q _12761_/Y _13540_/A vssd1 vssd1 vccd1 vccd1 _12763_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17160__S _17529_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14502_ _14743_/A _14731_/B _14758_/C vssd1 vssd1 vccd1 vccd1 _14504_/A sky130_fd_sc_hd__or3_4
XPHY_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11714_ _12130_/B _11708_/X _16949_/X _16950_/S vssd1 vssd1 vccd1 vccd1 hold209/A
+ sky130_fd_sc_hd__a22o_1
X_18270_ _20077_/CLK _18270_/D vssd1 vssd1 vccd1 vccd1 _18270_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15482_ _18564_/Q _15474_/A _18565_/Q vssd1 vssd1 vccd1 vccd1 _15482_/X sky130_fd_sc_hd__o21a_1
XPHY_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16564__A2 _16687_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12694_ _18970_/Q _12691_/X hold250/X _12692_/X vssd1 vssd1 vccd1 vccd1 _18970_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_187_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17221_ _17220_/X _13537_/B _17386_/S vssd1 vssd1 vccd1 vccd1 _17221_/X sky130_fd_sc_hd__mux2_2
XPHY_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14433_ _18379_/Q _14425_/A _14403_/X _14426_/A vssd1 vssd1 vccd1 vccd1 _18379_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11645_ _11645_/A _11645_/B _11645_/C vssd1 vssd1 vccd1 vccd1 _19547_/D sky130_fd_sc_hd__nor3_4
XPHY_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12586__B1 _12344_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17152_ _17151_/X _09477_/A _17536_/S vssd1 vssd1 vccd1 vccd1 _17152_/X sky130_fd_sc_hd__mux2_2
XPHY_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14364_ _18419_/Q _14352_/A _14312_/X _14353_/A vssd1 vssd1 vccd1 vccd1 _18419_/D
+ sky130_fd_sc_hd__a22o_1
Xinput15 input15/A vssd1 vssd1 vccd1 vccd1 input15/X sky130_fd_sc_hd__clkbuf_1
XFILLER_183_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11576_ _11576_/A _11609_/A vssd1 vssd1 vccd1 vccd1 _11577_/B sky130_fd_sc_hd__or2_2
Xinput26 input26/A vssd1 vssd1 vccd1 vccd1 input26/X sky130_fd_sc_hd__buf_1
XPHY_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12050__A2 _12016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput37 input37/A vssd1 vssd1 vccd1 vccd1 input37/X sky130_fd_sc_hd__clkbuf_2
XPHY_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput48 input48/A vssd1 vssd1 vccd1 vccd1 input48/X sky130_fd_sc_hd__clkbuf_4
X_16103_ _18237_/Q vssd1 vssd1 vccd1 vccd1 _16103_/Y sky130_fd_sc_hd__inv_2
X_13315_ _18850_/Q vssd1 vssd1 vccd1 vccd1 _13428_/C sky130_fd_sc_hd__clkinvlp_4
Xinput59 input59/A vssd1 vssd1 vccd1 vccd1 input59/X sky130_fd_sc_hd__buf_4
X_10527_ _10527_/A _11652_/B _15270_/B vssd1 vssd1 vccd1 vccd1 _10529_/C sky130_fd_sc_hd__or3_1
X_17083_ _17082_/X _15606_/A _17474_/S vssd1 vssd1 vccd1 vccd1 _17083_/X sky130_fd_sc_hd__mux2_1
X_14295_ _18453_/Q _14288_/X _13676_/X _14290_/X vssd1 vssd1 vccd1 vccd1 _18453_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_109_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12338__B1 _12100_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16034_ _18132_/Q vssd1 vssd1 vccd1 vccd1 _16034_/Y sky130_fd_sc_hd__inv_2
X_13246_ _18877_/Q _13241_/X _12602_/X _13243_/X vssd1 vssd1 vccd1 vccd1 _18877_/D
+ sky130_fd_sc_hd__a22o_1
X_10458_ _19826_/Q _10450_/A _10427_/X _10452_/A vssd1 vssd1 vccd1 vccd1 _19826_/D
+ sky130_fd_sc_hd__a22o_1
X_10389_ _11065_/A vssd1 vssd1 vccd1 vccd1 _14490_/A sky130_fd_sc_hd__clkbuf_2
X_13177_ _18910_/Q _13175_/Y _13177_/B1 _13176_/X vssd1 vssd1 vccd1 vccd1 _18910_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__17991__CLK _18169_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12128_ _19295_/Q _12094_/A _11924_/X _12096_/A vssd1 vssd1 vccd1 vccd1 _19295_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_151_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17985_ _19825_/CLK _17985_/D vssd1 vssd1 vccd1 vccd1 _17985_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17335__S _17545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19724_ _19795_/CLK _19724_/D repeater226/X vssd1 vssd1 vccd1 vccd1 _19724_/Q sky130_fd_sc_hd__dfrtp_4
X_12059_ _11869_/A _13642_/D _12056_/Y _11853_/A _12056_/A vssd1 vssd1 vccd1 vccd1
+ _19329_/D sky130_fd_sc_hd__a32o_1
X_16936_ _19480_/Q hold177/X _16946_/S vssd1 vssd1 vccd1 vccd1 _16936_/X sky130_fd_sc_hd__mux2_1
XFILLER_77_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11313__A1 _11487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12510__B1 _12408_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_237_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16867_ _15768_/Y _11214_/Y _17546_/S vssd1 vssd1 vccd1 vccd1 _16867_/X sky130_fd_sc_hd__mux2_1
X_19655_ _19847_/CLK _19655_/D repeater264/X vssd1 vssd1 vccd1 vccd1 _19655_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_26_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18606_ _19041_/CLK _18606_/D repeater263/X vssd1 vssd1 vccd1 vccd1 _18606_/Q sky130_fd_sc_hd__dfrtp_1
X_15818_ _18767_/Q vssd1 vssd1 vccd1 vccd1 _16750_/A sky130_fd_sc_hd__inv_2
X_19586_ _19591_/CLK _19586_/D hold363/X vssd1 vssd1 vccd1 vccd1 _19586_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_65_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16798_ _16797_/X _13555_/A _17386_/S vssd1 vssd1 vccd1 vccd1 _16798_/X sky130_fd_sc_hd__mux2_2
XFILLER_46_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18537_ _19825_/CLK _18537_/D repeater228/X vssd1 vssd1 vccd1 vccd1 _18537_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_34_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18590__RESET_B repeater269/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15749_ _15749_/A _15749_/B _15749_/C vssd1 vssd1 vccd1 vccd1 _17550_/S sky130_fd_sc_hd__and3_1
XFILLER_33_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16004__B2 _16003_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17070__S _17414_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09270_ _09270_/A vssd1 vssd1 vccd1 vccd1 _09271_/A sky130_fd_sc_hd__inv_2
XFILLER_33_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18468_ _18954_/CLK _18468_/D vssd1 vssd1 vccd1 vccd1 _18468_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17752__A1 _12058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19742__CLK _20070_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17419_ _17418_/X _12937_/Y _17459_/S vssd1 vssd1 vccd1 vccd1 _17419_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18399_ _18416_/CLK _18399_/D vssd1 vssd1 vccd1 vccd1 _18399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09089__A hold245/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16712__C1 _16711_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14723__A _14791_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12329__B1 _12083_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08985_ _16986_/S _09198_/A _08980_/Y _08981_/Y _08984_/X vssd1 vssd1 vccd1 vccd1
+ _08986_/A sky130_fd_sc_hd__o311a_1
XANTENNA__17245__S _17386_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12501__B1 _12392_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18678__RESET_B repeater252/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10698__A _14791_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09606_ _09474_/B _09605_/A _20013_/Q _09605_/Y _09567_/X vssd1 vssd1 vccd1 vccd1
+ _20013_/D sky130_fd_sc_hd__o221a_1
XANTENNA__16243__B2 _15914_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_232_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14254__B1 _13682_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_189_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09537_ _09470_/A _19299_/Q _20007_/Q _09534_/Y _09536_/X vssd1 vssd1 vccd1 vccd1
+ _09545_/B sky130_fd_sc_hd__o221a_1
XFILLER_197_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09468_ _09468_/A _09615_/A vssd1 vssd1 vccd1 vccd1 _09469_/B sky130_fd_sc_hd__or2_2
XPHY_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold327_A HWDATA[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09399_ _19390_/Q vssd1 vssd1 vccd1 vccd1 _09399_/Y sky130_fd_sc_hd__inv_2
XPHY_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12568__B1 _12386_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11430_ _19575_/Q vssd1 vssd1 vccd1 vccd1 _11560_/C sky130_fd_sc_hd__inv_2
XFILLER_137_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11361_ _11350_/X _11361_/B _11361_/C _11361_/D vssd1 vssd1 vccd1 vccd1 _11362_/D
+ sky130_fd_sc_hd__and4b_1
XANTENNA__19466__RESET_B repeater274/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10312_ _18619_/Q _18618_/Q _15697_/A vssd1 vssd1 vccd1 vccd1 _15578_/B sky130_fd_sc_hd__or3_4
X_13100_ _19176_/Q _13077_/A _13097_/Y _18910_/Q _13099_/X vssd1 vssd1 vccd1 vccd1
+ _13109_/B sky130_fd_sc_hd__o221a_1
XFILLER_137_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14080_ _14067_/X _14080_/B _14080_/C _14080_/D vssd1 vssd1 vccd1 vccd1 _14080_/X
+ sky130_fd_sc_hd__and4b_1
X_11292_ _18994_/Q vssd1 vssd1 vccd1 vccd1 _11292_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_30_HCLK _18641_/CLK vssd1 vssd1 vccd1 vccd1 _20085_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_3_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10243_ _19668_/Q vssd1 vssd1 vccd1 vccd1 _10243_/Y sky130_fd_sc_hd__inv_2
X_13031_ _18915_/Q vssd1 vssd1 vccd1 vccd1 _13087_/A sky130_fd_sc_hd__inv_2
XFILLER_180_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10174_ _10174_/A vssd1 vssd1 vccd1 vccd1 _10174_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_78_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16482__A1 _15199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17155__S _17566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11992__A _15776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17770_ _18315_/Q _18435_/Q _18427_/Q _18419_/Q _17923_/S0 _19646_/Q vssd1 vssd1
+ vccd1 vccd1 _17770_/X sky130_fd_sc_hd__mux4_1
XANTENNA__16482__B2 _16476_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14982_ _18064_/Q _14976_/X hold236/X _14979_/X vssd1 vssd1 vccd1 vccd1 _18064_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_78_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16721_ _16721_/A _16721_/B vssd1 vssd1 vccd1 vccd1 _16721_/Y sky130_fd_sc_hd__nor2_1
X_13933_ _18723_/Q _13932_/Y _13907_/X _13823_/B vssd1 vssd1 vccd1 vccd1 _18723_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_219_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16994__S _17490_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19440_ _20066_/CLK _19440_/D repeater193/X vssd1 vssd1 vccd1 vccd1 _19440_/Q sky130_fd_sc_hd__dfrtp_1
X_16652_ _16966_/X _16563_/X _17018_/X _16591_/X vssd1 vssd1 vccd1 vccd1 _16656_/A
+ sky130_fd_sc_hd__o22ai_4
X_13864_ _19208_/Q vssd1 vssd1 vccd1 vccd1 _13864_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_234_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15603_ _15606_/B _15602_/Y _15590_/X vssd1 vssd1 vccd1 vccd1 _15603_/X sky130_fd_sc_hd__o21a_1
XFILLER_62_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12815_ _19248_/Q vssd1 vssd1 vccd1 vccd1 _12815_/Y sky130_fd_sc_hd__inv_2
X_19371_ _19971_/CLK _19371_/D repeater241/X vssd1 vssd1 vccd1 vccd1 _19371_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_16_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16583_ _16583_/A _16583_/B vssd1 vssd1 vccd1 vccd1 _16583_/Y sky130_fd_sc_hd__nor2_1
X_13795_ _18717_/Q vssd1 vssd1 vccd1 vccd1 _13909_/C sky130_fd_sc_hd__inv_2
X_18322_ _18435_/CLK _18322_/D vssd1 vssd1 vccd1 vccd1 _18322_/Q sky130_fd_sc_hd__dfxtp_1
X_15534_ _18577_/Q _15530_/A _15530_/B _15533_/Y _15530_/Y vssd1 vssd1 vccd1 vccd1
+ _15535_/B sky130_fd_sc_hd__o32a_1
X_12746_ _19254_/Q vssd1 vssd1 vccd1 vccd1 _12746_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16537__A2 _16687_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18253_ _20076_/CLK _18253_/D vssd1 vssd1 vccd1 vccd1 _18253_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_230_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15465_ _18561_/Q vssd1 vssd1 vccd1 vccd1 _15467_/A sky130_fd_sc_hd__inv_2
XPHY_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12677_ _12677_/A vssd1 vssd1 vccd1 vccd1 _12677_/X sky130_fd_sc_hd__clkbuf_2
XPHY_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12328__A _12335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17204_ _17203_/X _09436_/Y _17529_/S vssd1 vssd1 vccd1 vccd1 _17204_/X sky130_fd_sc_hd__mux2_1
XPHY_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14416_ _18390_/Q _14409_/X _14415_/X _14411_/X vssd1 vssd1 vccd1 vccd1 _18390_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11628_ _11626_/A _11626_/B _11617_/A _11626_/Y vssd1 vssd1 vccd1 vccd1 _19556_/D
+ sky130_fd_sc_hd__a211oi_2
X_18184_ _18198_/CLK _18184_/D vssd1 vssd1 vccd1 vccd1 _18184_/Q sky130_fd_sc_hd__dfxtp_1
X_15396_ _15402_/A _17582_/X vssd1 vssd1 vccd1 vccd1 _18530_/D sky130_fd_sc_hd__and2_1
XFILLER_184_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17135_ _17134_/X _09860_/A _17414_/S vssd1 vssd1 vccd1 vccd1 _17135_/X sky130_fd_sc_hd__mux2_1
X_14347_ _19644_/Q vssd1 vssd1 vccd1 vccd1 _14450_/A sky130_fd_sc_hd__buf_1
XFILLER_129_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11559_ _11570_/B _11559_/B _11559_/C vssd1 vssd1 vccd1 vccd1 _11590_/A sky130_fd_sc_hd__or3_1
XFILLER_195_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17066_ _16622_/Y _15529_/Y _17474_/S vssd1 vssd1 vccd1 vccd1 _17066_/X sky130_fd_sc_hd__mux2_1
X_14278_ _18464_/Q _14272_/X _14277_/X _14275_/X vssd1 vssd1 vccd1 vccd1 _18464_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_171_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16017_ _18148_/Q vssd1 vssd1 vccd1 vccd1 _16017_/Y sky130_fd_sc_hd__inv_2
X_13229_ _13231_/A vssd1 vssd1 vccd1 vccd1 _13230_/A sky130_fd_sc_hd__inv_2
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19295__CLK _20115_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17896__S1 _18759_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17065__S _17518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17968_ _19842_/CLK _17968_/D vssd1 vssd1 vccd1 vccd1 _17968_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_214_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19707_ _19720_/CLK _19707_/D repeater201/X vssd1 vssd1 vccd1 vccd1 _19707_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16919_ _16918_/X _09485_/A _17482_/S vssd1 vssd1 vccd1 vccd1 _16919_/X sky130_fd_sc_hd__mux2_1
XANTENNA__18771__RESET_B repeater271/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16225__A1 _15226_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17899_ _17895_/X _17896_/X _17897_/X _17898_/X _18760_/Q _18761_/Q vssd1 vssd1 vccd1
+ vccd1 _17899_/X sky130_fd_sc_hd__mux4_2
XFILLER_65_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18700__RESET_B hold359/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19638_ _19847_/CLK _19638_/D repeater258/X vssd1 vssd1 vccd1 vccd1 _19638_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_81_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_213_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19569_ _19576_/CLK _19569_/D repeater255/X vssd1 vssd1 vccd1 vccd1 _19569_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_80_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_222_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09322_ _09322_/A vssd1 vssd1 vccd1 vccd1 _15722_/A sky130_fd_sc_hd__inv_2
XFILLER_230_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19977__RESET_B repeater193/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16528__A2 _15904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15736__B1 _10660_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09253_ _18652_/Q _20059_/Q _09253_/S vssd1 vssd1 vccd1 vccd1 _20059_/D sky130_fd_sc_hd__mux2_1
XFILLER_194_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17820__S1 _18750_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09184_ _14713_/A _09164_/A _09183_/X _09165_/A vssd1 vssd1 vccd1 vccd1 _20075_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_182_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_53_HCLK clkbuf_4_9_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19720_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__17489__A0 _15768_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11773__A1 hold196/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19638__CLK _19847_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09718__B2 _19415_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18859__RESET_B repeater232/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17887__S1 _18759_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16464__A1 _11742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08968_ _19860_/Q _08962_/Y _08964_/X _18772_/Q _08967_/X vssd1 vssd1 vccd1 vccd1
+ _08969_/D sky130_fd_sc_hd__o221a_1
XFILLER_29_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14475__B1 _14474_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11828__A2 _11800_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_229_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11317__A _18973_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10930_ _17726_/X _10923_/A _19675_/Q _10924_/A vssd1 vssd1 vccd1 vccd1 _19675_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_17_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10861_ _12232_/A vssd1 vssd1 vccd1 vccd1 _10861_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_232_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12600_ _12600_/A vssd1 vssd1 vccd1 vccd1 _12600_/X sky130_fd_sc_hd__clkbuf_2
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13580_ _13580_/A vssd1 vssd1 vccd1 vccd1 _13580_/Y sky130_fd_sc_hd__inv_2
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_242_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10792_ _19738_/Q _10794_/B _10788_/Y vssd1 vssd1 vccd1 vccd1 _19738_/D sky130_fd_sc_hd__a21o_1
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19647__RESET_B repeater261/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12531_ _19066_/Q _12528_/X _12302_/X _12529_/X vssd1 vssd1 vccd1 vccd1 _19066_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17811__S1 _18750_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15250_ _19778_/Q vssd1 vssd1 vccd1 vccd1 _15250_/Y sky130_fd_sc_hd__inv_2
XPHY_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12462_ _19111_/Q _12457_/X _12408_/X _12458_/X vssd1 vssd1 vccd1 vccd1 _19111_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_166_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14201_ _14200_/Y _18684_/Q _19101_/Q _14011_/A vssd1 vssd1 vccd1 vccd1 _14201_/X
+ sky130_fd_sc_hd__o22a_1
X_11413_ _19566_/Q vssd1 vssd1 vccd1 vccd1 _11579_/A sky130_fd_sc_hd__inv_2
X_15181_ _18488_/D vssd1 vssd1 vccd1 vccd1 _15744_/B sky130_fd_sc_hd__inv_2
XANTENNA__15459__A _15512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12393_ _19151_/Q _12388_/X _12392_/X _12390_/X vssd1 vssd1 vccd1 vccd1 _19151_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_115_HCLK_A clkbuf_opt_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14132_ _14132_/A vssd1 vssd1 vccd1 vccd1 _14135_/A sky130_fd_sc_hd__clkinvlp_2
X_11344_ _18970_/Q vssd1 vssd1 vccd1 vccd1 _11344_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16989__S _17548_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18940_ _19325_/CLK _18940_/D repeater213/X vssd1 vssd1 vccd1 vccd1 _18940_/Q sky130_fd_sc_hd__dfrtp_1
X_14063_ _14060_/Y _18702_/Q _19091_/Q _14032_/A _14062_/X vssd1 vssd1 vccd1 vccd1
+ _14063_/X sky130_fd_sc_hd__o221a_1
XFILLER_153_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11275_ _19604_/Q vssd1 vssd1 vccd1 vccd1 _11484_/A sky130_fd_sc_hd__inv_2
XANTENNA__14702__B2 _14701_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13014_ _13014_/A vssd1 vssd1 vccd1 vccd1 _13014_/Y sky130_fd_sc_hd__inv_2
X_10226_ _19836_/Q vssd1 vssd1 vccd1 vccd1 _10226_/Y sky130_fd_sc_hd__inv_2
X_18871_ _20058_/CLK _18871_/D repeater198/X vssd1 vssd1 vccd1 vccd1 _18871_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17878__S1 _18759_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15194__A _18757_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10157_ _19895_/Q _10154_/X _09082_/X _10156_/X vssd1 vssd1 vccd1 vccd1 _19895_/D
+ sky130_fd_sc_hd__a22o_1
X_17822_ _18358_/Q _17998_/Q _18414_/Q _18398_/Q _17918_/S0 _18750_/Q vssd1 vssd1
+ vccd1 vccd1 _17822_/X sky130_fd_sc_hd__mux4_2
XFILLER_66_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14466__B1 _14437_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12611__A _15769_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13269__B2 _17918_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10088_ _10088_/A _10088_/B vssd1 vssd1 vccd1 vccd1 _10088_/Y sky130_fd_sc_hd__nor2_2
X_17753_ _15296_/Y _11153_/Y _17753_/S vssd1 vssd1 vccd1 vccd1 _17753_/X sky130_fd_sc_hd__mux2_1
X_14965_ _14965_/A vssd1 vssd1 vccd1 vccd1 _14966_/A sky130_fd_sc_hd__inv_2
XFILLER_181_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17613__S _17614_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16704_ _17089_/X _16687_/X _16839_/X _16688_/X _16703_/X vssd1 vssd1 vccd1 vccd1
+ _16705_/C sky130_fd_sc_hd__o221a_1
X_13916_ _13916_/A _13970_/C _13916_/C vssd1 vssd1 vccd1 vccd1 _18732_/D sky130_fd_sc_hd__nor3_1
X_17684_ _15496_/Y _19451_/Q _17696_/S vssd1 vssd1 vccd1 vccd1 _18568_/D sky130_fd_sc_hd__mux2_1
X_14896_ _14897_/A vssd1 vssd1 vccd1 vccd1 _14896_/X sky130_fd_sc_hd__clkbuf_2
X_16635_ _16872_/X _16633_/X _16919_/X _16634_/X vssd1 vssd1 vccd1 vccd1 _16635_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_63_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19423_ _19470_/CLK _19423_/D repeater274/X vssd1 vssd1 vccd1 vccd1 _19423_/Q sky130_fd_sc_hd__dfrtp_2
X_13847_ _19215_/Q _13912_/D _13846_/Y _18705_/Q vssd1 vssd1 vccd1 vccd1 _13847_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_204_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19354_ _19968_/CLK _19354_/D hold370/X vssd1 vssd1 vccd1 vccd1 _19354_/Q sky130_fd_sc_hd__dfrtp_4
X_16566_ _17175_/X _16684_/A _17158_/X _16003_/X vssd1 vssd1 vccd1 vccd1 _16566_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__17707__A1 _19770_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13778_ _18734_/Q vssd1 vssd1 vccd1 vccd1 _13832_/A sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_76_HCLK clkbuf_opt_4_HCLK/A vssd1 vssd1 vccd1 vccd1 _18827_/CLK sky130_fd_sc_hd__clkbuf_16
X_18305_ _18416_/CLK _18305_/D vssd1 vssd1 vccd1 vccd1 _18305_/Q sky130_fd_sc_hd__dfxtp_1
X_15517_ _18574_/Q vssd1 vssd1 vccd1 vccd1 _15517_/Y sky130_fd_sc_hd__inv_2
X_12729_ _14814_/A vssd1 vssd1 vccd1 vccd1 _12729_/X sky130_fd_sc_hd__clkbuf_2
X_19285_ _19288_/CLK _19285_/D repeater211/X vssd1 vssd1 vccd1 vccd1 _19285_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12058__A _12058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17802__S1 _18750_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16497_ _17229_/X _16148_/X _17227_/X _15908_/X vssd1 vssd1 vccd1 vccd1 _16497_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_230_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18236_ _20076_/CLK _18236_/D vssd1 vssd1 vccd1 vccd1 _18236_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15448_ _18557_/Q vssd1 vssd1 vccd1 vccd1 _15450_/A sky130_fd_sc_hd__inv_2
XFILLER_164_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16472__B _16544_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18167_ _18169_/CLK _18167_/D vssd1 vssd1 vccd1 vccd1 _18167_/Q sky130_fd_sc_hd__dfxtp_1
X_15379_ _19795_/Q _10655_/B _10655_/X vssd1 vssd1 vccd1 vccd1 _15379_/X sky130_fd_sc_hd__a21bo_1
XFILLER_144_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14273__A _14273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17118_ _17117_/X _18901_/Q _17542_/S vssd1 vssd1 vccd1 vccd1 _17118_/X sky130_fd_sc_hd__mux2_1
XFILLER_190_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18098_ _18198_/CLK _18098_/D vssd1 vssd1 vccd1 vccd1 _18098_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16899__S _17513_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17049_ _15768_/Y _11220_/Y _17546_/S vssd1 vssd1 vccd1 vccd1 _17049_/X sky130_fd_sc_hd__mux2_1
X_09940_ _19947_/Q _16472_/A _19964_/Q _09939_/Y vssd1 vssd1 vccd1 vccd1 _09940_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12704__B1 _12538_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20060_ _20064_/CLK _20060_/D repeater199/X vssd1 vssd1 vccd1 vccd1 _20060_/Q sky130_fd_sc_hd__dfrtp_1
X_09871_ _09871_/A _09871_/B vssd1 vssd1 vccd1 vccd1 _09960_/A sky130_fd_sc_hd__or2_1
XANTENNA__18952__RESET_B repeater257/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17869__S1 _18761_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14457__B1 _14415_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater210 repeater243/X vssd1 vssd1 vccd1 vccd1 repeater210/X sky130_fd_sc_hd__buf_8
Xrepeater221 repeater223/X vssd1 vssd1 vccd1 vccd1 repeater221/X sky130_fd_sc_hd__buf_8
Xrepeater232 repeater233/X vssd1 vssd1 vccd1 vccd1 repeater232/X sky130_fd_sc_hd__buf_6
Xrepeater243 repeater244/X vssd1 vssd1 vccd1 vccd1 repeater243/X sky130_fd_sc_hd__buf_6
Xrepeater254 hold364/A vssd1 vssd1 vccd1 vccd1 hold366/A sky130_fd_sc_hd__buf_8
Xrepeater265 repeater267/X vssd1 vssd1 vccd1 vccd1 repeater265/X sky130_fd_sc_hd__buf_6
Xrepeater276 hold345/A vssd1 vssd1 vccd1 vccd1 hold364/A sky130_fd_sc_hd__buf_6
XANTENNA__17523__S _17523_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16647__B _16647_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20018__CLK _20091_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09305_ _18660_/Q _09305_/B vssd1 vssd1 vccd1 vccd1 _09305_/Y sky130_fd_sc_hd__nand2_1
XFILLER_222_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19058__RESET_B repeater257/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09236_ _19881_/Q _15709_/A _09233_/Y _09234_/Y _09235_/Y vssd1 vssd1 vccd1 vccd1
+ _09236_/X sky130_fd_sc_hd__o221a_1
XFILLER_210_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09167_ _20080_/Q vssd1 vssd1 vccd1 vccd1 _14703_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_79_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09098_ _12234_/A vssd1 vssd1 vccd1 vccd1 _09098_/X sky130_fd_sc_hd__buf_4
XANTENNA__16685__A1 _16962_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11060_ _19634_/Q vssd1 vssd1 vccd1 vccd1 _11060_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18693__RESET_B hold359/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10011_ _10011_/A _10011_/B _10101_/C vssd1 vssd1 vccd1 vccd1 _10081_/C sky130_fd_sc_hd__or3_1
XFILLER_88_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_192_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14448__B1 _14403_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17433__S _17568_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14750_ _18200_/Q _14744_/X _14749_/X _14747_/X vssd1 vssd1 vccd1 vccd1 _18200_/D
+ sky130_fd_sc_hd__a22o_1
X_11962_ _11977_/A vssd1 vssd1 vccd1 vccd1 _11962_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_1_1_1_HCLK clkbuf_1_1_1_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_17_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19899__RESET_B repeater195/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_99_HCLK clkbuf_4_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19214_/CLK sky130_fd_sc_hd__clkbuf_16
X_13701_ _13700_/A _13506_/A _18763_/Q _13700_/Y vssd1 vssd1 vccd1 vccd1 _18763_/D
+ sky130_fd_sc_hd__o22a_1
X_10913_ _19683_/Q vssd1 vssd1 vccd1 vccd1 _10913_/Y sky130_fd_sc_hd__inv_2
X_14681_ _14681_/A _15196_/A vssd1 vssd1 vccd1 vccd1 _14683_/A sky130_fd_sc_hd__or2_4
XANTENNA__19828__RESET_B repeater270/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14358__A hold245/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11893_ _19422_/Q _11891_/X hold314/X _11892_/X vssd1 vssd1 vccd1 vccd1 _19422_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_244_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16420_ _17976_/Q vssd1 vssd1 vccd1 vccd1 _16420_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13262__A _18751_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13632_ _10196_/B _12058_/B _13637_/B vssd1 vssd1 vccd1 vccd1 _13632_/Y sky130_fd_sc_hd__a21oi_1
X_10844_ _10844_/A vssd1 vssd1 vccd1 vccd1 _10845_/A sky130_fd_sc_hd__inv_2
X_16351_ _18272_/Q vssd1 vssd1 vccd1 vccd1 _16351_/Y sky130_fd_sc_hd__inv_2
X_13563_ _13563_/A vssd1 vssd1 vccd1 vccd1 _13563_/Y sky130_fd_sc_hd__inv_2
X_10775_ _17624_/X _10772_/X _19749_/Q _10774_/X vssd1 vssd1 vccd1 vccd1 _19749_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_212_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16573__A _16683_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15302_ _18627_/Q vssd1 vssd1 vccd1 vccd1 _15302_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17796__S0 _17923_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12514_ _19077_/Q _12512_/X _12413_/X _12513_/X vssd1 vssd1 vccd1 vccd1 _19077_/D
+ sky130_fd_sc_hd__a22o_1
X_19070_ _19610_/CLK _19070_/D hold361/X vssd1 vssd1 vccd1 vccd1 _19070_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__19410__RESET_B repeater193/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16282_ _18223_/Q vssd1 vssd1 vccd1 vccd1 _16282_/Y sky130_fd_sc_hd__inv_2
XFILLER_146_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13494_ _13494_/A _20086_/Q vssd1 vssd1 vccd1 vccd1 _13495_/B sky130_fd_sc_hd__nor2_1
X_18021_ _18145_/CLK _18021_/D vssd1 vssd1 vccd1 vccd1 _18021_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_5_HCLK clkbuf_4_2_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19630_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_157_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15233_ _15233_/A _15233_/B vssd1 vssd1 vccd1 vccd1 _15233_/Y sky130_fd_sc_hd__nor2_1
X_12445_ _19124_/Q _12441_/X _12375_/X _12444_/X vssd1 vssd1 vccd1 vccd1 _19124_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_repeater147_A _17683_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15164_ _17949_/Q _15158_/X _14707_/A _15160_/X vssd1 vssd1 vccd1 vccd1 _17949_/D
+ sky130_fd_sc_hd__a22o_1
X_12376_ _12427_/A vssd1 vssd1 vccd1 vccd1 _12428_/A sky130_fd_sc_hd__inv_2
XFILLER_153_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14115_ _14115_/A vssd1 vssd1 vccd1 vccd1 _14115_/Y sky130_fd_sc_hd__clkinv_1
X_11327_ _19578_/Q _11324_/Y _11477_/A _18979_/Q _11326_/X vssd1 vssd1 vccd1 vccd1
+ _11331_/C sky130_fd_sc_hd__o221a_1
X_15095_ _15096_/A vssd1 vssd1 vccd1 vccd1 _15095_/X sky130_fd_sc_hd__clkbuf_2
X_19972_ _19976_/CLK _19972_/D hold371/X vssd1 vssd1 vccd1 vccd1 _19972_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_141_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14687__B1 _14606_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14046_ _19068_/Q vssd1 vssd1 vccd1 vccd1 _14046_/Y sky130_fd_sc_hd__inv_2
X_18923_ _18947_/CLK _18923_/D repeater211/X vssd1 vssd1 vccd1 vccd1 _18923_/Q sky130_fd_sc_hd__dfrtp_1
X_11258_ _19023_/Q vssd1 vssd1 vccd1 vccd1 _11258_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10209_ _10209_/A _10209_/B _10209_/C _10209_/D vssd1 vssd1 vccd1 vccd1 _10209_/X
+ sky130_fd_sc_hd__or4_4
X_18854_ _18856_/CLK _18854_/D repeater231/X vssd1 vssd1 vccd1 vccd1 _18854_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_79_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11189_ _17713_/X _11184_/X _19618_/Q _11185_/X vssd1 vssd1 vccd1 vccd1 _19618_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10173__B1 _09090_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17805_ _18331_/Q _18211_/Q _18203_/Q _18195_/Q _17918_/S0 _18750_/Q vssd1 vssd1
+ vccd1 vccd1 _17805_/X sky130_fd_sc_hd__mux4_2
X_18785_ _19157_/CLK _18785_/D repeater265/X vssd1 vssd1 vccd1 vccd1 _18785_/Q sky130_fd_sc_hd__dfrtp_1
X_15997_ _16530_/A vssd1 vssd1 vccd1 vccd1 _15997_/X sky130_fd_sc_hd__buf_1
XANTENNA__17343__S _17564_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17736_ _15373_/X _19709_/Q _18508_/D vssd1 vssd1 vccd1 vccd1 _17736_/X sky130_fd_sc_hd__mux2_1
X_14948_ _18083_/Q _14940_/A _14935_/X _14941_/A vssd1 vssd1 vccd1 vccd1 _18083_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_236_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19333__CLK _20013_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16467__B _16469_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17667_ _15568_/X _19468_/Q _17683_/S vssd1 vssd1 vccd1 vccd1 _18585_/D sky130_fd_sc_hd__mux2_1
X_14879_ _18124_/Q _14872_/A _14711_/X _14873_/A vssd1 vssd1 vccd1 vccd1 _18124_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19406_ _19984_/CLK _19406_/D repeater210/X vssd1 vssd1 vccd1 vccd1 _19406_/Q sky130_fd_sc_hd__dfrtp_4
X_16618_ _16618_/A _16621_/B vssd1 vssd1 vccd1 vccd1 _16618_/Y sky130_fd_sc_hd__nor2_1
XFILLER_211_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17598_ _15340_/X _19705_/Q _17600_/S vssd1 vssd1 vccd1 vccd1 _17598_/X sky130_fd_sc_hd__mux2_1
XFILLER_51_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14611__B1 _14567_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16549_ _16723_/B vssd1 vssd1 vccd1 vccd1 _16622_/B sky130_fd_sc_hd__buf_2
X_19337_ _20013_/CLK _19337_/D repeater242/X vssd1 vssd1 vccd1 vccd1 _19337_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__16483__A _17565_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17787__S0 _17923_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19268_ _19283_/CLK _19268_/D repeater212/X vssd1 vssd1 vccd1 vccd1 _19268_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_31_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09021_ hold291/X vssd1 vssd1 vccd1 vccd1 _09021_/X sky130_fd_sc_hd__buf_4
X_18219_ _18268_/CLK _18219_/D vssd1 vssd1 vccd1 vccd1 _18219_/Q sky130_fd_sc_hd__dfxtp_1
X_19199_ _19221_/CLK _19199_/D hold365/X vssd1 vssd1 vccd1 vccd1 _19199_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_157_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20056__RESET_B repeater204/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09097__A _14793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold201 hold201/A vssd1 vssd1 vccd1 vccd1 hold201/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold212 hold212/A vssd1 vssd1 vccd1 vccd1 hold212/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold223 hold223/A vssd1 vssd1 vccd1 vccd1 hold223/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17864__A0 _17860_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold234 input44/X vssd1 vssd1 vccd1 vccd1 hold234/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17518__S _17518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold245 input65/X vssd1 vssd1 vccd1 vccd1 hold245/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold256 hold256/A vssd1 vssd1 vccd1 vccd1 hold256/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold267 hold267/A vssd1 vssd1 vccd1 vccd1 hold267/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_161_HCLK_A clkbuf_4_0_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20112_ _20122_/CLK _20112_/D repeater217/X vssd1 vssd1 vccd1 vccd1 _20112_/Q sky130_fd_sc_hd__dfrtp_1
Xhold278 HWDATA[16] vssd1 vssd1 vccd1 vccd1 input45/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09923_ _19965_/Q _09921_/Y _09848_/A _19331_/Q _09922_/X vssd1 vssd1 vccd1 vccd1
+ _09928_/C sky130_fd_sc_hd__o221a_1
Xhold289 input59/X vssd1 vssd1 vccd1 vccd1 hold289/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_59_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20043_ _20051_/CLK _20043_/D repeater209/X vssd1 vssd1 vccd1 vccd1 _20043_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_59_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09854_ _09854_/A _09854_/B vssd1 vssd1 vccd1 vccd1 _09992_/A sky130_fd_sc_hd__or2_1
XFILLER_100_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10164__B1 _09108_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09785_ _19985_/Q _09784_/Y _09731_/A _09742_/B vssd1 vssd1 vccd1 vccd1 _19985_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__17253__S _17512_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19992__RESET_B repeater192/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14850__B1 _14808_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09560__A _19325_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19921__RESET_B repeater230/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19239__RESET_B repeater239/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_241_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17778__S0 _17923_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10560_ _19808_/Q _19807_/Q _10572_/B vssd1 vssd1 vccd1 vccd1 _10576_/C sky130_fd_sc_hd__or3_1
XANTENNA__18850__CLK _18866_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19976__CLK _19976_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09219_ _09217_/Y _15714_/A _09217_/Y _15714_/A vssd1 vssd1 vccd1 vccd1 _09242_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_6_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10491_ _11655_/A _10491_/B _19539_/Q _10492_/C vssd1 vssd1 vccd1 vccd1 _10493_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_155_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_182_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12230_ _19233_/Q _12228_/X _11978_/X _12229_/X vssd1 vssd1 vccd1 vccd1 _19233_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_136_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18874__RESET_B repeater208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_205_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17428__S _19498_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12161_ _19276_/Q _12157_/X _12028_/X _12158_/X vssd1 vssd1 vccd1 vccd1 _19276_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_163_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11112_ _11116_/A _11116_/B vssd1 vssd1 vccd1 vccd1 _11113_/B sky130_fd_sc_hd__and2_1
XFILLER_122_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12092_ hold298/X vssd1 vssd1 vccd1 vccd1 _12092_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_1_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13257__A _18750_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_20_HCLK_A clkbuf_4_3_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15920_ _18019_/Q vssd1 vssd1 vccd1 vccd1 _15920_/Y sky130_fd_sc_hd__inv_2
X_11043_ _11043_/A _11043_/B vssd1 vssd1 vccd1 vccd1 _19647_/D sky130_fd_sc_hd__nor2_1
XFILLER_104_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_83_HCLK_A clkbuf_4_13_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_237_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15851_ _15848_/Y _15864_/B _15849_/Y _15828_/X _15850_/X vssd1 vssd1 vccd1 vccd1
+ _15851_/X sky130_fd_sc_hd__o221a_1
XANTENNA__17163__S _17386_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14802_ _14802_/A vssd1 vssd1 vccd1 vccd1 _14802_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_218_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15782_ _18138_/Q vssd1 vssd1 vccd1 vccd1 _15782_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18570_ _19437_/CLK _18570_/D repeater273/X vssd1 vssd1 vccd1 vccd1 _18570_/Q sky130_fd_sc_hd__dfrtp_1
X_12994_ _12994_/A vssd1 vssd1 vccd1 vccd1 _12994_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19662__RESET_B repeater270/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14733_ _14733_/A vssd1 vssd1 vccd1 vccd1 _14734_/A sky130_fd_sc_hd__inv_2
X_17521_ _17520_/X _15874_/Y _17539_/S vssd1 vssd1 vccd1 vccd1 _17521_/X sky130_fd_sc_hd__mux2_1
X_11945_ _19395_/Q _11939_/X hold288/X _11942_/X vssd1 vssd1 vccd1 vccd1 _19395_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_output114_A _15781_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17452_ _17486_/A0 _13110_/Y _17522_/S vssd1 vssd1 vccd1 vccd1 _17452_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14664_ _18244_/Q _14657_/A _14582_/X _14658_/A vssd1 vssd1 vccd1 vccd1 _18244_/D
+ sky130_fd_sc_hd__a22o_1
X_11876_ _11914_/A vssd1 vssd1 vccd1 vccd1 _11915_/A sky130_fd_sc_hd__inv_2
X_16403_ _18073_/Q vssd1 vssd1 vccd1 vccd1 _16403_/Y sky130_fd_sc_hd__inv_2
XFILLER_221_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13615_ _13613_/Y _17762_/S _18801_/Q _13620_/A vssd1 vssd1 vccd1 vccd1 _13616_/B
+ sky130_fd_sc_hd__o22a_1
X_10827_ _10698_/X _17750_/X _17750_/S _10823_/Y _19721_/Q vssd1 vssd1 vccd1 vccd1
+ _19721_/D sky130_fd_sc_hd__a32o_1
XANTENNA__09076__A1 _20101_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17383_ _16212_/Y _19370_/Q _17413_/S vssd1 vssd1 vccd1 vccd1 _17383_/X sky130_fd_sc_hd__mux2_1
X_14595_ _18284_/Q _14588_/A _14582_/X _14589_/A vssd1 vssd1 vccd1 vccd1 _18284_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17769__S0 _19647_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19122_ _19609_/CLK _19122_/D hold357/X vssd1 vssd1 vccd1 vccd1 _19122_/Q sky130_fd_sc_hd__dfrtp_2
X_16334_ _18040_/Q vssd1 vssd1 vccd1 vccd1 _16334_/Y sky130_fd_sc_hd__inv_2
X_13546_ _13546_/A _13580_/A vssd1 vssd1 vccd1 vccd1 _13547_/B sky130_fd_sc_hd__or2_2
XFILLER_186_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15149__B2 _15148_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10758_ _19754_/Q _10758_/B vssd1 vssd1 vccd1 vccd1 _19754_/D sky130_fd_sc_hd__and2_1
XFILLER_146_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19053_ _19157_/CLK _19053_/D repeater267/X vssd1 vssd1 vccd1 vccd1 _19053_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_187_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16265_ _18407_/Q vssd1 vssd1 vccd1 vccd1 _16265_/Y sky130_fd_sc_hd__inv_2
X_13477_ _18844_/Q _13476_/Y _13468_/B _13443_/X vssd1 vssd1 vccd1 vccd1 _18844_/D
+ sky130_fd_sc_hd__o211a_1
X_10689_ _11830_/B vssd1 vssd1 vccd1 vccd1 _12370_/B sky130_fd_sc_hd__buf_1
XFILLER_185_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15216_ _18481_/Q _18638_/Q _15216_/C vssd1 vssd1 vccd1 vccd1 _15217_/A sky130_fd_sc_hd__and3_1
X_18004_ _18416_/CLK _18004_/D vssd1 vssd1 vccd1 vccd1 _18004_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09379__A2 _09374_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12428_ _12428_/A vssd1 vssd1 vccd1 vccd1 _12428_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_106_HCLK clkbuf_4_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _18727_/CLK sky130_fd_sc_hd__clkbuf_16
X_16196_ _13749_/Y _17962_/Q _16195_/X vssd1 vssd1 vccd1 vccd1 _16196_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__12383__A1 _19155_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17338__S _17548_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15147_ _15147_/A vssd1 vssd1 vccd1 vccd1 _15148_/A sky130_fd_sc_hd__inv_2
XANTENNA__18544__RESET_B repeater232/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12359_ _19166_/Q _12352_/X _12225_/X _12354_/X vssd1 vssd1 vccd1 vccd1 _19166_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_141_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15078_ _18005_/Q _15071_/X _14793_/X _15073_/X vssd1 vssd1 vccd1 vccd1 _18005_/D
+ sky130_fd_sc_hd__a22o_1
X_19955_ _19956_/CLK _19955_/D repeater245/X vssd1 vssd1 vccd1 vccd1 _19955_/Q sky130_fd_sc_hd__dfrtp_1
X_14029_ _14029_/A _14104_/A vssd1 vssd1 vccd1 vccd1 _14030_/B sky130_fd_sc_hd__or2_2
XFILLER_101_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18906_ _18908_/CLK _18906_/D repeater212/X vssd1 vssd1 vccd1 vccd1 _18906_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_206_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19886_ _20066_/CLK _19886_/D repeater200/X vssd1 vssd1 vccd1 vccd1 _19886_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__10697__A1 _10451_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18837_ _18866_/CLK _18837_/D repeater231/X vssd1 vssd1 vccd1 vccd1 _18837_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__11894__B1 hold300/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17073__S _17385_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15382__A _19717_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09570_ _09494_/A _09494_/B _09495_/Y _09604_/B vssd1 vssd1 vccd1 vccd1 _20034_/D
+ sky130_fd_sc_hd__a211oi_2
X_18768_ _20058_/CLK _18768_/D repeater194/X vssd1 vssd1 vccd1 vccd1 _18768_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_222_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10449__A1 _19832_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17719_ _15421_/X _19522_/Q _18546_/D vssd1 vssd1 vccd1 vccd1 _17719_/X sky130_fd_sc_hd__mux2_1
XFILLER_223_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18699_ _18701_/CLK _18699_/D hold351/X vssd1 vssd1 vccd1 vccd1 _18699_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_222_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19332__RESET_B repeater245/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_223_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09004_ _19502_/Q _19501_/Q vssd1 vssd1 vccd1 vccd1 _11842_/D sky130_fd_sc_hd__or2_4
XFILLER_118_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17248__S _17513_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09906_ _19967_/Q _09905_/Y _09875_/A _19359_/Q vssd1 vssd1 vccd1 vccd1 _09906_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_99_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_219_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20026_ _20032_/CLK _20026_/D repeater239/X vssd1 vssd1 vccd1 vccd1 _20026_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_58_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09837_ _19949_/Q vssd1 vssd1 vccd1 vccd1 _09857_/A sky130_fd_sc_hd__inv_2
XFILLER_246_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15076__B1 hold244/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09768_ _09752_/A _09752_/B _09767_/X _09765_/Y vssd1 vssd1 vccd1 vccd1 _19996_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14823__B1 _14745_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09699_ _19991_/Q _09697_/Y _09747_/A _19420_/Q _09698_/X vssd1 vssd1 vccd1 vccd1
+ _09703_/C sky130_fd_sc_hd__o221a_1
XPHY_4046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer60 _14009_/B vssd1 vssd1 vccd1 vccd1 _14141_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_215_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17711__S _18546_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrebuffer71 _09729_/A vssd1 vssd1 vccd1 vccd1 _09735_/B sky130_fd_sc_hd__dlygate4sd1_1
XPHY_4068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11730_ _11730_/A vssd1 vssd1 vccd1 vccd1 _11730_/X sky130_fd_sc_hd__clkbuf_2
Xrebuffer82 _13066_/B vssd1 vssd1 vccd1 vccd1 _13208_/B1 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_4079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrebuffer93 _13068_/B vssd1 vssd1 vccd1 vccd1 _13203_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_199_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11661_ _11661_/A vssd1 vssd1 vccd1 vccd1 _11661_/Y sky130_fd_sc_hd__inv_2
XPHY_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13400_ _13399_/Y _13354_/A _20121_/Q _18867_/Q vssd1 vssd1 vccd1 vccd1 _13400_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10612_ _18553_/Q vssd1 vssd1 vccd1 vccd1 _10612_/Y sky130_fd_sc_hd__inv_2
XPHY_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14380_ _14381_/A vssd1 vssd1 vccd1 vccd1 _14380_/X sky130_fd_sc_hd__clkbuf_2
XPHY_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11592_ _11592_/A vssd1 vssd1 vccd1 vccd1 _11592_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_129_HCLK clkbuf_4_4_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19561_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13331_ _18848_/Q vssd1 vssd1 vccd1 vccd1 _13333_/C sky130_fd_sc_hd__inv_2
XFILLER_168_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10543_ _19798_/Q _19797_/Q _19800_/Q _19799_/Q vssd1 vssd1 vccd1 vccd1 _10577_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_195_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_2_1_0_HCLK clkbuf_2_1_0_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_3_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XPHY_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11060__A _19634_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16050_ _19711_/Q vssd1 vssd1 vccd1 vccd1 _16050_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13262_ _18751_/Q _13262_/B vssd1 vssd1 vccd1 vccd1 _13737_/B sky130_fd_sc_hd__nand2_1
X_10474_ _17698_/X _10471_/X _19821_/Q _10472_/X vssd1 vssd1 vccd1 vccd1 _19821_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_155_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15001_ _18054_/Q _14991_/X _15000_/X _14994_/X vssd1 vssd1 vccd1 vccd1 _18054_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17158__S _17536_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13562__B1 _13597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12213_ _12229_/A vssd1 vssd1 vccd1 vccd1 _12213_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__09766__C1 _09759_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13193_ _13193_/A vssd1 vssd1 vccd1 vccd1 _13193_/Y sky130_fd_sc_hd__inv_2
XFILLER_163_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17923__S0 _17923_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10107__C _10107_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12144_ _12151_/A vssd1 vssd1 vccd1 vccd1 _12144_/X sky130_fd_sc_hd__buf_1
XFILLER_69_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16997__S _17534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19740_ _20051_/CLK _19740_/D repeater206/X vssd1 vssd1 vccd1 vccd1 _19740_/Q sky130_fd_sc_hd__dfrtp_1
X_12075_ _19324_/Q _12068_/X _12074_/X _12072_/X vssd1 vssd1 vccd1 vccd1 _19324_/D
+ sky130_fd_sc_hd__a22o_1
X_16952_ _17774_/X _18790_/Q _16957_/S vssd1 vssd1 vccd1 vccd1 _16952_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11026_ _11026_/A vssd1 vssd1 vccd1 vccd1 _11026_/Y sky130_fd_sc_hd__inv_2
X_15903_ _16494_/A vssd1 vssd1 vccd1 vccd1 _15904_/A sky130_fd_sc_hd__buf_1
X_19671_ _19812_/CLK _19671_/D repeater225/X vssd1 vssd1 vccd1 vccd1 _19671_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA__19843__RESET_B repeater270/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16883_ _16882_/X _09677_/Y _17523_/S vssd1 vssd1 vccd1 vccd1 _16883_/X sky130_fd_sc_hd__mux2_1
X_18622_ _19859_/CLK _18622_/D repeater262/X vssd1 vssd1 vccd1 vccd1 _18622_/Q sky130_fd_sc_hd__dfrtp_1
X_15834_ _19709_/Q vssd1 vssd1 vccd1 vccd1 _15834_/Y sky130_fd_sc_hd__inv_2
XFILLER_46_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18553_ _19810_/CLK _18553_/D repeater226/X vssd1 vssd1 vccd1 vccd1 _18553_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_18_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11628__B1 _11617_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15765_ _19764_/Q _19520_/Q _15765_/C vssd1 vssd1 vccd1 vccd1 _15765_/X sky130_fd_sc_hd__and3_1
X_12977_ _12885_/A _12885_/B _12975_/Y _13027_/C vssd1 vssd1 vccd1 vccd1 _18943_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_205_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17504_ _15939_/Y _15936_/Y _17564_/S vssd1 vssd1 vccd1 vccd1 _17504_/X sky130_fd_sc_hd__mux2_1
X_14716_ _14743_/A _14731_/B _15082_/C vssd1 vssd1 vccd1 vccd1 _14718_/A sky130_fd_sc_hd__or3_4
X_11928_ _11933_/A _12309_/A vssd1 vssd1 vccd1 vccd1 _11929_/S sky130_fd_sc_hd__or2_1
XFILLER_233_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18484_ _19545_/CLK _18484_/D repeater225/X vssd1 vssd1 vccd1 vccd1 _18484_/Q sky130_fd_sc_hd__dfrtp_1
X_15696_ _18617_/Q vssd1 vssd1 vccd1 vccd1 _15696_/Y sky130_fd_sc_hd__inv_2
XPHY_4580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17435_ _17434_/X _16094_/Y _17565_/S vssd1 vssd1 vccd1 vccd1 _17435_/X sky130_fd_sc_hd__mux2_1
X_14647_ _18256_/Q _14643_/X _09171_/X _14645_/X vssd1 vssd1 vccd1 vccd1 _18256_/D
+ sky130_fd_sc_hd__a22o_1
X_11859_ _12058_/B vssd1 vssd1 vccd1 vccd1 _13630_/A sky130_fd_sc_hd__inv_2
XFILLER_177_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14546__A _14547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14578_ _14791_/A vssd1 vssd1 vccd1 vccd1 _14578_/X sky130_fd_sc_hd__clkbuf_2
X_17366_ _15768_/Y _11280_/Y _17546_/S vssd1 vssd1 vccd1 vccd1 _17366_/X sky130_fd_sc_hd__mux2_1
XANTENNA__18796__RESET_B repeater258/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19105_ _19109_/CLK _19105_/D hold361/X vssd1 vssd1 vccd1 vccd1 _19105_/Q sky130_fd_sc_hd__dfrtp_1
X_13529_ _13529_/A _13610_/A vssd1 vssd1 vccd1 vccd1 _13530_/B sky130_fd_sc_hd__or2_2
X_16317_ _15250_/Y _15840_/A _16316_/Y _15842_/X vssd1 vssd1 vccd1 vccd1 _16317_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17297_ _17486_/A0 _16502_/Y _17517_/S vssd1 vssd1 vccd1 vccd1 _17297_/X sky130_fd_sc_hd__mux2_1
XANTENNA__18725__RESET_B repeater253/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19036_ _19157_/CLK _19036_/D repeater267/X vssd1 vssd1 vccd1 vccd1 _19036_/Q sky130_fd_sc_hd__dfrtp_1
X_16248_ _17390_/X _16595_/A _17399_/X _15999_/A vssd1 vssd1 vccd1 vccd1 _16248_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_173_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17068__S _17482_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput103 _16743_/Y vssd1 vssd1 vccd1 vccd1 HRDATA[31] sky130_fd_sc_hd__clkbuf_2
Xoutput114 _15781_/X vssd1 vssd1 vccd1 vccd1 IRQ[11] sky130_fd_sc_hd__clkbuf_2
X_16179_ _17949_/Q vssd1 vssd1 vccd1 vccd1 _16179_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput125 _15777_/X vssd1 vssd1 vccd1 vccd1 IRQ[7] sky130_fd_sc_hd__clkbuf_2
Xoutput136 _19610_/Q vssd1 vssd1 vccd1 vccd1 pwm_S6 sky130_fd_sc_hd__clkbuf_2
XANTENNA__17914__S0 _19633_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19938_ _20013_/CLK _19938_/D repeater243/X vssd1 vssd1 vccd1 vccd1 _19938_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_101_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19869_ _20050_/CLK _19869_/D repeater197/X vssd1 vssd1 vccd1 vccd1 _19869_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_229_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09622_ _20004_/Q _10079_/A _09618_/A _09581_/X vssd1 vssd1 vccd1 vccd1 _20004_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_83_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14805__B1 _14802_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09553_ _20005_/Q _09551_/Y _20031_/Q _09552_/Y vssd1 vssd1 vccd1 vccd1 _09553_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__17531__S _17537_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09484_ _09484_/A _09484_/B vssd1 vssd1 vccd1 vccd1 _09584_/A sky130_fd_sc_hd__or2_1
XANTENNA__12292__B1 _12035_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20071__RESET_B repeater207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20000__RESET_B repeater192/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09996__C1 _09964_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12347__A1 _19172_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_191_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17905__S0 _17908_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10190_ _11869_/A _19329_/Q vssd1 vssd1 vccd1 vccd1 _13642_/B sky130_fd_sc_hd__or2_2
XFILLER_87_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17706__S _18546_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11322__A2 _18986_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12900_ _12897_/Y _18930_/Q _19273_/Q _12870_/C _12899_/X vssd1 vssd1 vccd1 vccd1
+ _12908_/B sky130_fd_sc_hd__o221a_1
X_20009_ _20013_/CLK _20009_/D repeater240/X vssd1 vssd1 vccd1 vccd1 _20009_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_101_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13880_ _19215_/Q _13912_/D _19214_/Q _13909_/A vssd1 vssd1 vccd1 vccd1 _13880_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_247_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12831_ _19258_/Q _12829_/Y _19251_/Q _13551_/A vssd1 vssd1 vccd1 vccd1 _12831_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_36_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17441__S _17517_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15550_ _18581_/Q _15550_/B vssd1 vssd1 vccd1 vccd1 _15555_/B sky130_fd_sc_hd__or2_1
XFILLER_215_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12762_ _18817_/Q vssd1 vssd1 vccd1 vccd1 _13540_/A sky130_fd_sc_hd__inv_2
XFILLER_199_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_202_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14501_ _18338_/Q _14492_/A _14268_/X _14493_/A vssd1 vssd1 vccd1 vccd1 _18338_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_215_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11713_ _12370_/A _11708_/X _16950_/X _16950_/S vssd1 vssd1 vccd1 vccd1 hold205/A
+ sky130_fd_sc_hd__a22o_1
XPHY_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15481_ _15481_/A vssd1 vssd1 vccd1 vccd1 _15487_/B sky130_fd_sc_hd__inv_2
X_12693_ _18971_/Q _12691_/X hold239/X _12692_/X vssd1 vssd1 vccd1 vccd1 _18971_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_230_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17220_ _17219_/X _13377_/Y _17385_/S vssd1 vssd1 vccd1 vccd1 _17220_/X sky130_fd_sc_hd__mux2_1
XPHY_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14432_ _18380_/Q _14425_/A _14419_/X _14426_/A vssd1 vssd1 vccd1 vccd1 _18380_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11644_ _11639_/A _11639_/B _11639_/C vssd1 vssd1 vccd1 vccd1 _11645_/B sky130_fd_sc_hd__o21a_1
XPHY_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17151_ _17150_/X _09458_/Y _17529_/S vssd1 vssd1 vccd1 vccd1 _17151_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14363_ _18420_/Q _14352_/A _14329_/X _14353_/A vssd1 vssd1 vccd1 vccd1 _18420_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11575_ _11575_/A _11575_/B vssd1 vssd1 vccd1 vccd1 _11609_/A sky130_fd_sc_hd__or2_1
Xinput16 input16/A vssd1 vssd1 vccd1 vccd1 input16/X sky130_fd_sc_hd__clkbuf_1
XPHY_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput27 input27/A vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_hd__buf_1
XPHY_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16102_ _18253_/Q vssd1 vssd1 vccd1 vccd1 _16102_/Y sky130_fd_sc_hd__inv_2
X_13314_ _18851_/Q vssd1 vssd1 vccd1 vccd1 _13430_/B sky130_fd_sc_hd__inv_6
Xinput38 input38/A vssd1 vssd1 vccd1 vccd1 input38/X sky130_fd_sc_hd__buf_6
XFILLER_6_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10526_ _19532_/Q _10526_/B _19531_/Q vssd1 vssd1 vccd1 vccd1 _15270_/B sky130_fd_sc_hd__nor3b_4
Xinput49 input49/A vssd1 vssd1 vccd1 vccd1 input49/X sky130_fd_sc_hd__buf_4
X_17082_ _17473_/A0 _16439_/Y _17473_/S vssd1 vssd1 vccd1 vccd1 _17082_/X sky130_fd_sc_hd__mux2_1
X_14294_ _18454_/Q _14288_/X _13674_/X _14290_/X vssd1 vssd1 vccd1 vccd1 _18454_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_6_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16033_ _18220_/Q vssd1 vssd1 vccd1 vccd1 _16033_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19694__CLK _20051_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13245_ _18878_/Q _13241_/X _12599_/X _13243_/X vssd1 vssd1 vccd1 vccd1 _18878_/D
+ sky130_fd_sc_hd__a22o_1
X_10457_ _19827_/Q _10450_/X _10425_/X _10452_/X vssd1 vssd1 vccd1 vccd1 _19827_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_109_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12614__A _12650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13176_ _13180_/A vssd1 vssd1 vccd1 vccd1 _13176_/X sky130_fd_sc_hd__buf_2
X_10388_ _19851_/Q vssd1 vssd1 vccd1 vccd1 _11065_/A sky130_fd_sc_hd__inv_2
XFILLER_69_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12127_ _19296_/Q _12121_/X _11922_/X _12122_/X vssd1 vssd1 vccd1 vccd1 _19296_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_69_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17984_ _20124_/CLK _17984_/D vssd1 vssd1 vccd1 vccd1 _17984_/Q sky130_fd_sc_hd__dfxtp_1
X_19723_ _19795_/CLK _19723_/D repeater218/X vssd1 vssd1 vccd1 vccd1 _19723_/Q sky130_fd_sc_hd__dfrtp_1
X_12058_ _12058_/A _12058_/B vssd1 vssd1 vccd1 vccd1 _13642_/D sky130_fd_sc_hd__or2_1
X_16935_ _19479_/Q hold180/X _16946_/S vssd1 vssd1 vccd1 vccd1 _16935_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12510__A1 _19079_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11313__A2 _18989_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11009_ _11009_/A vssd1 vssd1 vccd1 vccd1 _11010_/B sky130_fd_sc_hd__inv_2
X_19654_ _19855_/CLK _19654_/D repeater264/X vssd1 vssd1 vccd1 vccd1 _19654_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_77_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16866_ _16865_/X _09866_/A _17524_/S vssd1 vssd1 vccd1 vccd1 _16866_/X sky130_fd_sc_hd__mux2_1
XFILLER_93_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18605_ _19041_/CLK _18605_/D repeater263/X vssd1 vssd1 vccd1 vccd1 _18605_/Q sky130_fd_sc_hd__dfrtp_4
X_15817_ _18106_/Q vssd1 vssd1 vccd1 vccd1 _15817_/Y sky130_fd_sc_hd__inv_2
X_19585_ _19585_/CLK _19585_/D hold361/X vssd1 vssd1 vccd1 vccd1 _19585_/Q sky130_fd_sc_hd__dfrtp_4
X_16797_ _16796_/X _16706_/Y _17535_/S vssd1 vssd1 vccd1 vccd1 _16797_/X sky130_fd_sc_hd__mux2_1
XFILLER_53_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17351__S _17543_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18536_ _19825_/CLK _18536_/D repeater228/X vssd1 vssd1 vccd1 vccd1 _18536_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12274__B1 _12090_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15748_ _15746_/Y _18485_/Q _10584_/D _15747_/X vssd1 vssd1 vccd1 vccd1 _18482_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_179_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16004__A2 _16002_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20051__CLK _20051_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10824__A1 _10446_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18467_ _18954_/CLK _18467_/D vssd1 vssd1 vccd1 vccd1 _18467_/Q sky130_fd_sc_hd__dfxtp_1
X_15679_ _15683_/B _15678_/X _15643_/X vssd1 vssd1 vccd1 vccd1 _15679_/X sky130_fd_sc_hd__o21a_1
XANTENNA__18906__RESET_B repeater212/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17418_ _17486_/A0 _13145_/Y _17543_/S vssd1 vssd1 vccd1 vccd1 _17418_/X sky130_fd_sc_hd__mux2_1
XANTENNA__16960__A0 _15963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18398_ _18416_/CLK _18398_/D vssd1 vssd1 vccd1 vccd1 _18398_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17349_ _17486_/A0 _16299_/Y _17517_/S vssd1 vssd1 vccd1 vccd1 _17349_/X sky130_fd_sc_hd__mux2_1
XFILLER_147_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19019_ _19609_/CLK _19019_/D hold357/X vssd1 vssd1 vccd1 vccd1 _19019_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_228_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17526__S _17548_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08984_ _20072_/Q _20071_/Q _20073_/Q _08983_/X vssd1 vssd1 vccd1 vccd1 _08984_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_114_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_244_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09605_ _09605_/A vssd1 vssd1 vccd1 vccd1 _09605_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16243__A2 _15883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15451__B1 _15571_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_232_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17261__S _17543_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09536_ _20027_/Q _09535_/Y _09476_/A _19306_/Q vssd1 vssd1 vccd1 vccd1 _09536_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12265__B1 _12074_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19399__D _19399_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09467_ _09467_/A _09467_/B vssd1 vssd1 vccd1 vccd1 _09615_/A sky130_fd_sc_hd__or2_1
XFILLER_240_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09398_ _19930_/Q vssd1 vssd1 vccd1 vccd1 _10046_/A sky130_fd_sc_hd__inv_2
XPHY_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13214__C1 _13176_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11360_ _11460_/A _18961_/Q _19594_/Q _11348_/Y _11359_/X vssd1 vssd1 vccd1 vccd1
+ _11361_/D sky130_fd_sc_hd__o221a_1
XFILLER_22_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10311_ _18617_/Q _18616_/Q _15693_/A vssd1 vssd1 vccd1 vccd1 _15697_/A sky130_fd_sc_hd__or3_4
XFILLER_125_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11291_ _19603_/Q _11286_/Y _11483_/A _19017_/Q _11290_/X vssd1 vssd1 vccd1 vccd1
+ _11298_/C sky130_fd_sc_hd__o221a_1
XFILLER_138_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17259__A1 _18977_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13030_ _18916_/Q vssd1 vssd1 vccd1 vccd1 _13088_/A sky130_fd_sc_hd__clkinvlp_2
X_10242_ _19841_/Q vssd1 vssd1 vccd1 vccd1 _10242_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17436__S _17566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10173_ _19883_/Q _10166_/X _09090_/X _10168_/X vssd1 vssd1 vccd1 vccd1 _19883_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10751__B1 _10427_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11992__B _11998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14981_ hold237/X vssd1 vssd1 vccd1 vccd1 hold236/A sky130_fd_sc_hd__buf_2
XFILLER_93_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16720_ _16720_/A _16721_/B vssd1 vssd1 vccd1 vccd1 _16720_/Y sky130_fd_sc_hd__nor2_1
XFILLER_247_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13932_ _13932_/A vssd1 vssd1 vccd1 vccd1 _13932_/Y sky130_fd_sc_hd__inv_2
XFILLER_93_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17431__A1 _08952_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_234_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16651_ _19047_/Q _16673_/B vssd1 vssd1 vccd1 vccd1 _16651_/Y sky130_fd_sc_hd__nand2_1
X_13863_ _19193_/Q vssd1 vssd1 vccd1 vccd1 _13863_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17171__S _17535_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12814_ _19231_/Q _13532_/A _12810_/Y _18807_/Q _12813_/X vssd1 vssd1 vccd1 vccd1
+ _12833_/A sky130_fd_sc_hd__o221a_1
X_15602_ _15602_/A _15602_/B vssd1 vssd1 vccd1 vccd1 _15602_/Y sky130_fd_sc_hd__nor2_1
XFILLER_74_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_138_HCLK_A clkbuf_4_3_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19370_ _19971_/CLK _19370_/D repeater241/X vssd1 vssd1 vccd1 vccd1 _19370_/Q sky130_fd_sc_hd__dfrtp_4
X_16582_ _16582_/A _16583_/B vssd1 vssd1 vccd1 vccd1 _16582_/Y sky130_fd_sc_hd__nor2_1
X_13794_ _18718_/Q vssd1 vssd1 vccd1 vccd1 _13911_/B sky130_fd_sc_hd__inv_2
XFILLER_188_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18321_ _19637_/CLK _18321_/D vssd1 vssd1 vccd1 vccd1 _18321_/Q sky130_fd_sc_hd__dfxtp_1
X_12745_ _19245_/Q _13545_/A _12741_/Y _18827_/Q _12744_/X vssd1 vssd1 vccd1 vccd1
+ _12758_/B sky130_fd_sc_hd__o221a_1
X_15533_ _18577_/Q vssd1 vssd1 vccd1 vccd1 _15533_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_repeater177_A _17518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12008__B1 _09027_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15464_ _15467_/B _15463_/Y _15459_/X vssd1 vssd1 vccd1 vccd1 _15464_/X sky130_fd_sc_hd__o21a_1
X_18252_ _18268_/CLK _18252_/D vssd1 vssd1 vccd1 vccd1 _18252_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12676_ _18982_/Q _12670_/X hold298/X _12671_/X vssd1 vssd1 vccd1 vccd1 _18982_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_179_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17203_ _15963_/X _09559_/Y _17534_/S vssd1 vssd1 vccd1 vccd1 _17203_/X sky130_fd_sc_hd__mux2_1
XPHY_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14415_ hold325/X vssd1 vssd1 vccd1 vccd1 _14415_/X sky130_fd_sc_hd__buf_2
XPHY_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11627_ _19557_/Q _11626_/Y _11588_/A _11571_/B vssd1 vssd1 vccd1 vccd1 _19557_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15395_ _18530_/Q _13217_/B _13218_/B vssd1 vssd1 vccd1 vccd1 _15395_/X sky130_fd_sc_hd__a21bo_1
X_18183_ _18198_/CLK _18183_/D vssd1 vssd1 vccd1 vccd1 _18183_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14346_ _18426_/Q _14337_/A _14314_/X _14338_/A vssd1 vssd1 vccd1 vccd1 _18426_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17134_ _17133_/X _09723_/Y _17413_/S vssd1 vssd1 vccd1 vccd1 _17134_/X sky130_fd_sc_hd__mux2_1
X_11558_ _11582_/A _11581_/A _11584_/A _11583_/A vssd1 vssd1 vccd1 vccd1 _11559_/C
+ sky130_fd_sc_hd__or4_4
XFILLER_144_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10509_ _15270_/A _17609_/X vssd1 vssd1 vccd1 vccd1 _11653_/A sky130_fd_sc_hd__or2b_1
XFILLER_195_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17065_ _17064_/X _19959_/Q _17518_/S vssd1 vssd1 vccd1 vccd1 _17065_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14277_ _14277_/A vssd1 vssd1 vccd1 vccd1 _14277_/X sky130_fd_sc_hd__buf_2
XFILLER_155_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11489_ _11489_/A vssd1 vssd1 vccd1 vccd1 _11489_/Y sky130_fd_sc_hd__inv_2
X_16016_ _18012_/Q vssd1 vssd1 vccd1 vccd1 _16016_/Y sky130_fd_sc_hd__inv_2
X_13228_ _18541_/Q _13228_/B vssd1 vssd1 vccd1 vccd1 _13231_/A sky130_fd_sc_hd__or2_2
XFILLER_170_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17346__S _17564_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13159_ _13159_/A _13159_/B _13159_/C _13159_/D vssd1 vssd1 vccd1 vccd1 _13160_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_111_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19176__RESET_B repeater212/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17967_ _19842_/CLK _17967_/D vssd1 vssd1 vccd1 vccd1 _17967_/Q sky130_fd_sc_hd__dfxtp_1
X_19706_ _19720_/CLK _19706_/D repeater202/X vssd1 vssd1 vccd1 vccd1 _19706_/Q sky130_fd_sc_hd__dfstp_1
X_16918_ _16917_/X _09431_/Y _17529_/S vssd1 vssd1 vccd1 vccd1 _16918_/X sky130_fd_sc_hd__mux2_1
XFILLER_214_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12495__B1 _12382_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17898_ _15952_/Y _15953_/Y _15954_/Y _15955_/Y _17908_/S0 _18759_/Q vssd1 vssd1
+ vccd1 vccd1 _17898_/X sky130_fd_sc_hd__mux4_2
XFILLER_226_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19637_ _19637_/CLK _19637_/D repeater258/X vssd1 vssd1 vccd1 vccd1 _19637_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_226_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16849_ _16848_/X _14057_/Y _17490_/S vssd1 vssd1 vccd1 vccd1 _16849_/X sky130_fd_sc_hd__mux2_2
XFILLER_65_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17081__S _17524_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_214_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19568_ _19576_/CLK _19568_/D repeater282/X vssd1 vssd1 vccd1 vccd1 _19568_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_206_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09321_ _18654_/Q _09317_/X _18654_/Q _09317_/X vssd1 vssd1 vccd1 vccd1 _09322_/A
+ sky130_fd_sc_hd__o2bb2a_1
X_18519_ _19814_/CLK _18519_/D repeater223/X vssd1 vssd1 vccd1 vccd1 _18519_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_222_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19499_ _20036_/CLK _19499_/D repeater194/X vssd1 vssd1 vccd1 vccd1 _19499_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_230_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12519__A _12528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09252_ _20059_/Q _20060_/Q _09253_/S vssd1 vssd1 vccd1 vccd1 _20060_/D sky130_fd_sc_hd__mux2_1
XFILLER_21_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_221_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09183_ _14711_/A vssd1 vssd1 vccd1 vccd1 _09183_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__10039__A _10039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09415__B2 _09414_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19946__RESET_B repeater244/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17256__S _17318_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08967_ _10324_/A _18778_/Q _19858_/Q _08966_/Y vssd1 vssd1 vccd1 vccd1 _08967_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_248_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12486__B1 _12241_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold172_A HADDR[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18899__RESET_B repeater188/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_216_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18828__RESET_B repeater239/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_216_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10860_ _19706_/Q _10855_/X _10451_/X _10857_/X vssd1 vssd1 vccd1 vccd1 _19706_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_204_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09519_ _09490_/A _19320_/Q _20015_/Q _09518_/Y vssd1 vssd1 vccd1 vccd1 _09519_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_25_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10791_ _10791_/A _13766_/D vssd1 vssd1 vccd1 vccd1 _10794_/B sky130_fd_sc_hd__or2_1
XFILLER_24_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11333__A _18977_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12530_ _19067_/Q _12528_/X _12299_/X _12529_/X vssd1 vssd1 vccd1 vccd1 _19067_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_235_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_240_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12461_ _19112_/Q _12457_/X _12406_/X _12458_/X vssd1 vssd1 vccd1 vccd1 _19112_/D
+ sky130_fd_sc_hd__a22o_1
X_14200_ _19105_/Q vssd1 vssd1 vccd1 vccd1 _14200_/Y sky130_fd_sc_hd__inv_2
XFILLER_184_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11412_ _11412_/A _11412_/B _11412_/C _11412_/D vssd1 vssd1 vccd1 vccd1 _11457_/B
+ sky130_fd_sc_hd__and4_1
X_15180_ _17937_/Q _15171_/A _09255_/X _15172_/A vssd1 vssd1 vccd1 vccd1 _17937_/D
+ sky130_fd_sc_hd__a22o_1
X_12392_ hold308/X vssd1 vssd1 vccd1 vccd1 _12392_/X sky130_fd_sc_hd__buf_2
X_14131_ _14014_/A _14131_/A2 _14129_/Y _14118_/X vssd1 vssd1 vccd1 vccd1 _18684_/D
+ sky130_fd_sc_hd__a211oi_2
X_11343_ _19604_/Q _11341_/Y _11459_/A _18960_/Q _11342_/X vssd1 vssd1 vccd1 vccd1
+ _11347_/C sky130_fd_sc_hd__o221a_1
XFILLER_152_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14062_ _14061_/Y _18698_/Q _19072_/Q _14013_/A vssd1 vssd1 vccd1 vccd1 _14062_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09709__A2 _19421_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_180_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11274_ _19602_/Q vssd1 vssd1 vccd1 vccd1 _11482_/A sky130_fd_sc_hd__inv_2
XFILLER_153_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17166__S _17536_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13013_ _13006_/A _13006_/B _13011_/Y _12986_/A vssd1 vssd1 vccd1 vccd1 _18927_/D
+ sky130_fd_sc_hd__a211oi_2
X_10225_ _19656_/Q vssd1 vssd1 vccd1 vccd1 _10956_/D sky130_fd_sc_hd__inv_2
XFILLER_152_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18870_ _20036_/CLK _18870_/D repeater199/X vssd1 vssd1 vccd1 vccd1 _18870_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__10724__B1 _10448_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17821_ _18190_/Q _18182_/Q _18174_/Q _18158_/Q _17918_/S0 _18750_/Q vssd1 vssd1
+ vccd1 vccd1 _17821_/X sky130_fd_sc_hd__mux4_1
X_10156_ _10156_/A vssd1 vssd1 vccd1 vccd1 _10156_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_output144_A _19671_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17752_ _15296_/Y _12058_/A _17756_/S vssd1 vssd1 vccd1 vccd1 _17752_/X sky130_fd_sc_hd__mux2_2
XANTENNA__12477__B1 _12296_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10087_ _10087_/A _10091_/A vssd1 vssd1 vccd1 vccd1 _10088_/B sky130_fd_sc_hd__or2_4
X_14964_ _14965_/A vssd1 vssd1 vccd1 vccd1 _14964_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_59_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09342__A0 _09255_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20103__RESET_B repeater233/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17404__A1 _17874_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16703_ _16827_/X _16637_/X _16841_/X _16638_/X vssd1 vssd1 vccd1 vccd1 _16703_/X
+ sky130_fd_sc_hd__o22a_1
X_13915_ _13830_/B _13829_/A _13914_/X _13830_/A vssd1 vssd1 vccd1 vccd1 _13916_/C
+ sky130_fd_sc_hd__o31a_1
XANTENNA__18569__RESET_B repeater272/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17683_ _15500_/X _19452_/Q _17683_/S vssd1 vssd1 vccd1 vccd1 _18569_/D sky130_fd_sc_hd__mux2_1
X_14895_ _15109_/A _15145_/B _15121_/C vssd1 vssd1 vccd1 vccd1 _14897_/A sky130_fd_sc_hd__or3_4
XFILLER_47_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19422_ _19997_/CLK _19422_/D repeater271/X vssd1 vssd1 vccd1 vccd1 _19422_/Q sky130_fd_sc_hd__dfrtp_2
X_16634_ _16634_/A vssd1 vssd1 vccd1 vccd1 _16634_/X sky130_fd_sc_hd__clkbuf_2
X_13846_ _19194_/Q vssd1 vssd1 vccd1 vccd1 _13846_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17168__A0 _17473_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19353_ _19968_/CLK _19353_/D hold371/X vssd1 vssd1 vccd1 vccd1 _19353_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_204_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16565_ _17116_/X _16563_/X _17169_/X _15908_/X _16564_/X vssd1 vssd1 vccd1 vccd1
+ _16565_/X sky130_fd_sc_hd__o221a_1
X_13777_ _18736_/Q _13202_/X _13776_/Y vssd1 vssd1 vccd1 vccd1 _18736_/D sky130_fd_sc_hd__o21a_1
X_10989_ _10989_/A vssd1 vssd1 vccd1 vccd1 _10989_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_62_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18304_ _18416_/CLK _18304_/D vssd1 vssd1 vccd1 vccd1 _18304_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15516_ _15535_/A _15516_/B vssd1 vssd1 vccd1 vccd1 _15516_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__16915__A0 _17473_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12728_ _18953_/Q vssd1 vssd1 vccd1 vccd1 _14816_/A sky130_fd_sc_hd__clkbuf_2
X_19284_ _19288_/CLK _19284_/D repeater211/X vssd1 vssd1 vccd1 vccd1 _19284_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_148_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16496_ _17218_/X _15896_/X _17221_/X _16493_/X _16495_/X vssd1 vssd1 vccd1 vccd1
+ _16496_/X sky130_fd_sc_hd__o221a_2
XFILLER_176_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18235_ _20076_/CLK _18235_/D vssd1 vssd1 vccd1 vccd1 _18235_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_230_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12659_ _12659_/A _12659_/B vssd1 vssd1 vccd1 vccd1 _12698_/A sky130_fd_sc_hd__or2_4
X_15447_ _15479_/A _15447_/B vssd1 vssd1 vccd1 vccd1 _17683_/S sky130_fd_sc_hd__nor2_8
XANTENNA__16391__A1 _17326_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18166_ _18169_/CLK _18166_/D vssd1 vssd1 vccd1 vccd1 _18166_/Q sky130_fd_sc_hd__dfxtp_1
X_15378_ _19794_/Q _10654_/B _10655_/B vssd1 vssd1 vccd1 vccd1 _15378_/X sky130_fd_sc_hd__a21bo_1
XFILLER_172_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17117_ _16544_/Y _19276_/Q _17541_/S vssd1 vssd1 vccd1 vccd1 _17117_/X sky130_fd_sc_hd__mux2_1
X_14329_ _14727_/A vssd1 vssd1 vccd1 vccd1 _14329_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__19357__RESET_B hold371/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18097_ _20090_/CLK _18097_/D vssd1 vssd1 vccd1 vccd1 _18097_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12074__A hold291/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16143__B2 _15915_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17048_ _17047_/X _13859_/Y _17545_/S vssd1 vssd1 vccd1 vccd1 _17048_/X sky130_fd_sc_hd__mux2_1
XFILLER_131_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17076__S _17548_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09870_ _09870_/A _09963_/A vssd1 vssd1 vccd1 vccd1 _09871_/B sky130_fd_sc_hd__or2_2
XANTENNA__16446__A2 _15830_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18999_ _19137_/CLK _18999_/D repeater249/X vssd1 vssd1 vccd1 vccd1 _18999_/Q sky130_fd_sc_hd__dfrtp_1
Xrepeater200 repeater206/X vssd1 vssd1 vccd1 vccd1 repeater200/X sky130_fd_sc_hd__buf_6
XFILLER_97_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater211 repeater212/X vssd1 vssd1 vccd1 vccd1 repeater211/X sky130_fd_sc_hd__buf_8
Xrepeater222 repeater225/X vssd1 vssd1 vccd1 vccd1 repeater222/X sky130_fd_sc_hd__buf_8
Xrepeater233 repeater234/X vssd1 vssd1 vccd1 vccd1 repeater233/X sky130_fd_sc_hd__buf_8
XANTENNA__12468__B1 hold281/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater244 repeater245/X vssd1 vssd1 vccd1 vccd1 repeater244/X sky130_fd_sc_hd__buf_8
XFILLER_238_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater255 repeater266/X vssd1 vssd1 vccd1 vccd1 repeater255/X sky130_fd_sc_hd__buf_8
XFILLER_66_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater266 repeater267/X vssd1 vssd1 vccd1 vccd1 repeater266/X sky130_fd_sc_hd__buf_4
XFILLER_54_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater277 hold362/A vssd1 vssd1 vccd1 vccd1 hold345/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__14209__A1 _19113_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17159__A0 _15963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_20_HCLK clkbuf_4_3_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20059_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_clkbuf_leaf_121_HCLK_A clkbuf_opt_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09304_ _09304_/A vssd1 vssd1 vccd1 vccd1 _09305_/B sky130_fd_sc_hd__inv_2
XANTENNA__11153__A _19627_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12640__B1 _12028_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09235_ _19881_/Q _15709_/A vssd1 vssd1 vccd1 vccd1 _09235_/Y sky130_fd_sc_hd__nand2_1
XFILLER_166_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_194_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09166_ _14699_/A _09163_/X hold344/X _09165_/X vssd1 vssd1 vccd1 vccd1 _20081_/D
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_162_HCLK clkbuf_4_0_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19510_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_107_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_175_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19098__RESET_B repeater252/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09097_ _14793_/A vssd1 vssd1 vccd1 vccd1 _12234_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_134_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19027__RESET_B repeater269/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17925__D _19672_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15295__A _15318_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10010_ _19935_/Q vssd1 vssd1 vccd1 vccd1 _10022_/C sky130_fd_sc_hd__inv_2
XFILLER_95_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09999_ _19942_/Q _09998_/Y _09968_/A _09852_/B vssd1 vssd1 vccd1 vccd1 _19942_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_130_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17714__S _18546_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12459__B1 _12401_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_185_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11961_ _19383_/Q _11955_/X _09051_/X _11956_/X vssd1 vssd1 vccd1 vccd1 _19383_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18662__RESET_B repeater204/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10912_ _19682_/Q _19681_/Q _10912_/C vssd1 vssd1 vccd1 vccd1 _10914_/A sky130_fd_sc_hd__or3_1
X_13700_ _13700_/A _14641_/B vssd1 vssd1 vccd1 vccd1 _13700_/Y sky130_fd_sc_hd__nor2_1
X_14680_ _14680_/A _14680_/B vssd1 vssd1 vccd1 vccd1 _15196_/A sky130_fd_sc_hd__or2_4
X_11892_ _11892_/A vssd1 vssd1 vccd1 vccd1 _11892_/X sky130_fd_sc_hd__buf_1
XFILLER_205_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13631_ _11869_/A _13641_/B _19873_/Q _13630_/B vssd1 vssd1 vccd1 vccd1 _13637_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_44_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10843_ _10844_/A vssd1 vssd1 vccd1 vccd1 _10843_/X sky130_fd_sc_hd__buf_1
XFILLER_198_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13562_ _13557_/A _13557_/B _13597_/A _13558_/Y vssd1 vssd1 vccd1 vccd1 _18834_/D
+ sky130_fd_sc_hd__a211oi_2
X_16350_ _17975_/Q vssd1 vssd1 vccd1 vccd1 _16350_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12631__B1 _12401_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10774_ _10774_/A vssd1 vssd1 vccd1 vccd1 _10774_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_9_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17796__S1 _19646_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12513_ _12529_/A vssd1 vssd1 vccd1 vccd1 _12513_/X sky130_fd_sc_hd__buf_1
X_15301_ _19884_/Q vssd1 vssd1 vccd1 vccd1 _15301_/Y sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_43_HCLK_A clkbuf_opt_2_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_212_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11998__A _11998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16281_ _18239_/Q vssd1 vssd1 vccd1 vccd1 _16281_/Y sky130_fd_sc_hd__inv_2
X_13493_ _13493_/A vssd1 vssd1 vccd1 vccd1 _15319_/B sky130_fd_sc_hd__inv_2
X_18020_ _18142_/CLK _18020_/D vssd1 vssd1 vccd1 vccd1 _18020_/Q sky130_fd_sc_hd__dfxtp_1
X_12444_ _12458_/A vssd1 vssd1 vccd1 vccd1 _12444_/X sky130_fd_sc_hd__buf_1
X_15232_ _15232_/A _15232_/B _15232_/C vssd1 vssd1 vccd1 vccd1 _15232_/X sky130_fd_sc_hd__and3_1
XFILLER_154_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12934__A1 _19266_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15163_ _17950_/Q _15158_/X _14705_/A _15160_/X vssd1 vssd1 vccd1 vccd1 _17950_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_3_0_0_HCLK_A clkbuf_3_1_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12375_ hold284/X vssd1 vssd1 vccd1 vccd1 _12375_/X sky130_fd_sc_hd__buf_2
XANTENNA__19450__RESET_B repeater271/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14114_ _14024_/A _14114_/A2 _14111_/Y _14135_/B vssd1 vssd1 vccd1 vccd1 _18694_/D
+ sky130_fd_sc_hd__a211oi_2
X_11326_ _19606_/Q _11325_/Y _11486_/A _18988_/Q vssd1 vssd1 vccd1 vccd1 _11326_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_4_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19971_ _19971_/CLK _19971_/D repeater241/X vssd1 vssd1 vccd1 vccd1 _19971_/Q sky130_fd_sc_hd__dfrtp_1
X_15094_ _15094_/A _15094_/B _15094_/C vssd1 vssd1 vccd1 vccd1 _15096_/A sky130_fd_sc_hd__or3_4
X_14045_ _14042_/Y _18699_/Q _19075_/Q _14016_/A _14044_/Y vssd1 vssd1 vccd1 vccd1
+ _14045_/X sky130_fd_sc_hd__o221a_1
XFILLER_107_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18922_ _19290_/CLK _18922_/D repeater211/X vssd1 vssd1 vccd1 vccd1 _18922_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_141_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_180_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11257_ _19586_/Q _19000_/Q _11467_/A _16466_/A vssd1 vssd1 vccd1 vccd1 _11261_/C
+ sky130_fd_sc_hd__o22a_1
XFILLER_68_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10208_ _19840_/Q _19667_/Q _10206_/Y _10967_/A vssd1 vssd1 vccd1 vccd1 _10209_/D
+ sky130_fd_sc_hd__o22a_1
X_18853_ _18866_/CLK _18853_/D repeater231/X vssd1 vssd1 vccd1 vccd1 _18853_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_95_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11188_ _17712_/X _11184_/X _19619_/Q _11185_/X vssd1 vssd1 vccd1 vccd1 _19619_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_94_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17804_ _17800_/X _17801_/X _17802_/X _17803_/X _18751_/Q _18752_/Q vssd1 vssd1 vccd1
+ vccd1 _17804_/X sky130_fd_sc_hd__mux4_2
XFILLER_94_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10139_ _16986_/X _10136_/X _19903_/Q _10138_/X vssd1 vssd1 vccd1 vccd1 _19903_/D
+ sky130_fd_sc_hd__o22a_1
X_18784_ _19157_/CLK _18784_/D repeater267/X vssd1 vssd1 vccd1 vccd1 _18784_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_227_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15996_ _17482_/X _16512_/A _17479_/X _16513_/A _15995_/X vssd1 vssd1 vccd1 vccd1
+ _15996_/X sky130_fd_sc_hd__o221a_1
XFILLER_208_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_43_HCLK clkbuf_opt_2_HCLK/A vssd1 vssd1 vccd1 vccd1 _19545_/CLK sky130_fd_sc_hd__clkbuf_16
X_17735_ _15374_/X _19710_/Q _18508_/D vssd1 vssd1 vccd1 vccd1 _17735_/X sky130_fd_sc_hd__mux2_1
X_14947_ _18084_/Q _14940_/A _14933_/X _14941_/A vssd1 vssd1 vccd1 vccd1 _18084_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_36_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17666_ _15571_/Y _19469_/Q _17683_/S vssd1 vssd1 vccd1 vccd1 _18586_/D sky130_fd_sc_hd__mux2_1
XFILLER_208_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14878_ _18125_/Q _14871_/X _14709_/X _14873_/X vssd1 vssd1 vccd1 vccd1 _18125_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19405_ _19984_/CLK _19405_/D repeater243/X vssd1 vssd1 vccd1 vccd1 _19405_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_23_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16617_ _16617_/A _16621_/B vssd1 vssd1 vccd1 vccd1 _16617_/Y sky130_fd_sc_hd__nor2_1
X_13829_ _13829_/A _13829_/B vssd1 vssd1 vccd1 vccd1 _13917_/A sky130_fd_sc_hd__or2_1
X_17597_ _15342_/X _19706_/Q _17600_/S vssd1 vssd1 vccd1 vccd1 _17597_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12069__A hold284/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_211_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19336_ _20013_/CLK _19336_/D repeater242/X vssd1 vssd1 vccd1 vccd1 _19336_/Q sky130_fd_sc_hd__dfrtp_1
X_16548_ _16548_/A _16583_/B vssd1 vssd1 vccd1 vccd1 _16548_/Y sky130_fd_sc_hd__nor2_1
XFILLER_149_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17787__S1 _19646_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19538__RESET_B repeater221/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19267_ _19283_/CLK _19267_/D repeater212/X vssd1 vssd1 vccd1 vccd1 _19267_/Q sky130_fd_sc_hd__dfrtp_1
X_16479_ _17026_/X _16555_/A _17028_/X _16556_/A vssd1 vssd1 vccd1 vccd1 _16479_/Y
+ sky130_fd_sc_hd__a22oi_4
X_09020_ _20122_/Q _09015_/X _09016_/X _09019_/X vssd1 vssd1 vccd1 vccd1 _20122_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_148_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14375__B1 _14329_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18218_ _18268_/CLK _18218_/D vssd1 vssd1 vccd1 vccd1 _18218_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__19778__CLK _19780_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19198_ _19222_/CLK _19198_/D hold365/X vssd1 vssd1 vccd1 vccd1 _19198_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__09809__C _09813_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18149_ _18165_/CLK _18149_/D vssd1 vssd1 vccd1 vccd1 _18149_/Q sky130_fd_sc_hd__dfxtp_1
Xhold202 input12/X vssd1 vssd1 vccd1 vccd1 hold202/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold213 hold213/A vssd1 vssd1 vccd1 vccd1 hold213/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold224 hold224/A vssd1 vssd1 vccd1 vccd1 hold224/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold235 HWDATA[15] vssd1 vssd1 vccd1 vccd1 input44/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold246 HWDATA[5] vssd1 vssd1 vccd1 vccd1 input65/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20096__RESET_B repeater233/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold257 input42/X vssd1 vssd1 vccd1 vccd1 hold257/X sky130_fd_sc_hd__dlygate4sd3_1
X_20111_ _20122_/CLK _20111_/D repeater217/X vssd1 vssd1 vccd1 vccd1 _20111_/Q sky130_fd_sc_hd__dfrtp_2
Xhold268 input69/X vssd1 vssd1 vccd1 vccd1 hold268/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold279 input58/X vssd1 vssd1 vccd1 vccd1 hold279/X sky130_fd_sc_hd__dlygate4sd3_1
X_09922_ _09872_/A _19356_/Q _09858_/A _19342_/Q vssd1 vssd1 vccd1 vccd1 _09922_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_236_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12689__B1 _12030_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12532__A hold326/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09853_ _09853_/A _09995_/A vssd1 vssd1 vccd1 vccd1 _09854_/B sky130_fd_sc_hd__or2_2
X_20042_ _20066_/CLK _20042_/D repeater209/X vssd1 vssd1 vccd1 vccd1 _20042_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_59_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17534__S _17534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09784_ _09784_/A vssd1 vssd1 vccd1 vccd1 _09784_/Y sky130_fd_sc_hd__inv_2
XFILLER_105_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18182__CLK _18198_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19961__RESET_B hold371/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17778__S1 _19646_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19279__RESET_B repeater212/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09218_ _18649_/Q _09212_/B _09213_/A vssd1 vssd1 vccd1 vccd1 _15714_/A sky130_fd_sc_hd__o21ai_1
XFILLER_210_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10490_ _19538_/Q _19537_/Q _11654_/A vssd1 vssd1 vccd1 vccd1 _10492_/C sky130_fd_sc_hd__or3_1
XANTENNA_hold302_A HWDATA[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17709__S _18546_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09149_ _09149_/A vssd1 vssd1 vccd1 vccd1 _09156_/A sky130_fd_sc_hd__buf_1
XFILLER_151_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12160_ _19277_/Q _12157_/X _12026_/X _12158_/X vssd1 vssd1 vccd1 vccd1 _19277_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_100_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11111_ _11110_/Y _17754_/S _19637_/Q _11091_/X vssd1 vssd1 vccd1 vccd1 _11116_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_107_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12091_ _19317_/Q _12082_/X _12090_/X _12084_/X vssd1 vssd1 vccd1 vccd1 _19317_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_146_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12442__A _12478_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11042_ _17752_/X _10268_/B _10263_/X vssd1 vssd1 vccd1 vccd1 _11043_/B sky130_fd_sc_hd__a21oi_1
XFILLER_89_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_66_HCLK clkbuf_opt_3_HCLK/A vssd1 vssd1 vccd1 vccd1 _20107_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_77_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18843__RESET_B repeater233/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17444__S _17517_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15850_ _15850_/A _15850_/B vssd1 vssd1 vccd1 vccd1 _15850_/X sky130_fd_sc_hd__or2_1
XFILLER_130_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_237_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input20_A HADDR[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14801_ _14803_/A vssd1 vssd1 vccd1 vccd1 _14801_/X sky130_fd_sc_hd__clkbuf_2
X_15781_ _19870_/Q _19438_/Q vssd1 vssd1 vccd1 vccd1 _15781_/X sky130_fd_sc_hd__and2_4
X_12993_ _12877_/A _12877_/B _12991_/Y _12986_/X vssd1 vssd1 vccd1 vccd1 _18935_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_29_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17520_ _17519_/X _10004_/Y _17548_/S vssd1 vssd1 vccd1 vccd1 _17520_/X sky130_fd_sc_hd__mux2_1
XFILLER_245_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14732_ _14733_/A vssd1 vssd1 vccd1 vccd1 _14732_/X sky130_fd_sc_hd__clkbuf_2
X_11944_ _19396_/Q _11939_/X _09021_/X _11942_/X vssd1 vssd1 vccd1 vccd1 _19396_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_55_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17451_ _17450_/X _13530_/A _17536_/S vssd1 vssd1 vccd1 vccd1 _17451_/X sky130_fd_sc_hd__mux2_4
XFILLER_45_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14663_ _18245_/Q _14656_/X _14580_/X _14658_/X vssd1 vssd1 vccd1 vccd1 _18245_/D
+ sky130_fd_sc_hd__a22o_1
X_11875_ _11891_/A vssd1 vssd1 vccd1 vccd1 _11875_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_output107_A _16397_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16402_ _17993_/Q vssd1 vssd1 vccd1 vccd1 _16402_/Y sky130_fd_sc_hd__inv_2
X_10826_ _10451_/A _17750_/X _17750_/S _10823_/Y _19722_/Q vssd1 vssd1 vccd1 vccd1
+ _19722_/D sky130_fd_sc_hd__a32o_1
X_13614_ _13620_/A vssd1 vssd1 vccd1 vccd1 _17762_/S sky130_fd_sc_hd__inv_2
XFILLER_220_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12604__B1 _12533_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17382_ _17381_/X _19943_/Q _17414_/S vssd1 vssd1 vccd1 vccd1 _17382_/X sky130_fd_sc_hd__mux2_2
X_14594_ _18285_/Q _14587_/X _14580_/X _14589_/X vssd1 vssd1 vccd1 vccd1 _18285_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19920__CLK _19920_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19121_ _19609_/CLK _19121_/D hold357/X vssd1 vssd1 vccd1 vccd1 _19121_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17769__S1 _19648_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16333_ _18072_/Q vssd1 vssd1 vccd1 vccd1 _16333_/Y sky130_fd_sc_hd__inv_2
X_10757_ _19755_/Q _10754_/Y _17985_/Q _10754_/A _15389_/B vssd1 vssd1 vccd1 vccd1
+ _19755_/D sky130_fd_sc_hd__o221a_1
X_13545_ _13545_/A _13545_/B vssd1 vssd1 vccd1 vccd1 _13580_/A sky130_fd_sc_hd__or2_1
XANTENNA__15149__A2 _15146_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19631__RESET_B repeater258/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_repeater257_A repeater258/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19052_ _19157_/CLK _19052_/D repeater268/X vssd1 vssd1 vccd1 vccd1 _19052_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_118_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13476_ _13476_/A vssd1 vssd1 vccd1 vccd1 _13476_/Y sky130_fd_sc_hd__inv_2
X_16264_ _18343_/Q vssd1 vssd1 vccd1 vccd1 _16264_/Y sky130_fd_sc_hd__inv_2
X_10688_ _11935_/B vssd1 vssd1 vccd1 vccd1 _11830_/B sky130_fd_sc_hd__inv_2
XFILLER_139_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18003_ _19847_/CLK _18003_/D vssd1 vssd1 vccd1 vccd1 _18003_/Q sky130_fd_sc_hd__dfxtp_1
X_15215_ _15224_/A _15215_/B vssd1 vssd1 vccd1 vccd1 _15388_/A sky130_fd_sc_hd__or2_2
X_12427_ _12427_/A vssd1 vssd1 vccd1 vccd1 _12427_/X sky130_fd_sc_hd__clkbuf_2
X_16195_ _18745_/Q _15819_/Y _13749_/Y _17962_/Q vssd1 vssd1 vccd1 vccd1 _16195_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_154_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12358_ _19167_/Q _12352_/X _12223_/X _12354_/X vssd1 vssd1 vccd1 vccd1 _19167_/D
+ sky130_fd_sc_hd__a22o_1
X_15146_ _15147_/A vssd1 vssd1 vccd1 vccd1 _15146_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__20008__CLK _20013_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11309_ _11467_/A _18968_/Q _11475_/A _18977_/Q vssd1 vssd1 vccd1 vccd1 _11309_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15077_ _18006_/Q _15071_/X _14791_/X _15073_/X vssd1 vssd1 vccd1 vccd1 _18006_/D
+ sky130_fd_sc_hd__a22o_1
X_19954_ _19956_/CLK _19954_/D repeater245/X vssd1 vssd1 vccd1 vccd1 _19954_/Q sky130_fd_sc_hd__dfrtp_1
X_12289_ _19205_/Q _12283_/X _12032_/X _12284_/X vssd1 vssd1 vccd1 vccd1 _19205_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_114_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19300__CLK _20013_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14028_ _14028_/A _14028_/B vssd1 vssd1 vccd1 vccd1 _14104_/A sky130_fd_sc_hd__or2_1
X_18905_ _18908_/CLK _18905_/D repeater188/X vssd1 vssd1 vccd1 vccd1 _18905_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_113_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19885_ _20050_/CLK _19885_/D repeater200/X vssd1 vssd1 vccd1 vccd1 _19885_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18584__RESET_B repeater274/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17354__S _17534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18836_ _19900_/CLK _18836_/D repeater196/X vssd1 vssd1 vccd1 vccd1 _18836_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_68_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11894__A1 _19421_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18767_ _20058_/CLK _18767_/D repeater271/X vssd1 vssd1 vccd1 vccd1 _18767_/Q sky130_fd_sc_hd__dfrtp_1
X_15979_ _15967_/Y _15864_/B _15969_/X _15978_/X vssd1 vssd1 vccd1 vccd1 _15979_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_48_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14279__A _14279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17718_ _15422_/X _19523_/Q _18546_/D vssd1 vssd1 vccd1 vccd1 _17718_/X sky130_fd_sc_hd__mux2_1
XFILLER_222_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18698_ _18701_/CLK _18698_/D hold359/X vssd1 vssd1 vccd1 vccd1 _18698_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_36_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17649_ _15638_/X _19040_/Q _17655_/S vssd1 vssd1 vccd1 vccd1 _18603_/D sky130_fd_sc_hd__mux2_1
XFILLER_91_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_223_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14596__B1 _14567_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_223_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_220_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19319_ _19320_/CLK _19319_/D repeater213/X vssd1 vssd1 vccd1 vccd1 _19319_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_188_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17534__A0 _17533_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19372__RESET_B repeater241/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09003_ _10686_/C vssd1 vssd1 vccd1 vccd1 _10186_/A sky130_fd_sc_hd__buf_1
XANTENNA__17529__S _17529_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_89_HCLK clkbuf_4_12_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19952_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_105_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09905_ _19359_/Q vssd1 vssd1 vccd1 vccd1 _09905_/Y sky130_fd_sc_hd__inv_2
XANTENNA__10137__A1 _17919_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18548__CLK _19780_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17264__S _17534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20025_ _20091_/CLK _20025_/D repeater238/X vssd1 vssd1 vccd1 vccd1 _20025_/Q sky130_fd_sc_hd__dfrtp_1
X_09836_ _19950_/Q vssd1 vssd1 vccd1 vccd1 _09858_/A sky130_fd_sc_hd__inv_2
XFILLER_219_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09767_ _09767_/A vssd1 vssd1 vccd1 vccd1 _09767_/X sky130_fd_sc_hd__buf_2
XANTENNA__13093__A _19166_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold252_A HWDATA[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09698_ _09792_/A _19409_/Q _09792_/A _19409_/Q vssd1 vssd1 vccd1 vccd1 _09698_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_132_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrebuffer50 _18730_/Q vssd1 vssd1 vccd1 vccd1 _13873_/B2 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_4047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19943__CLK _19984_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrebuffer61 _14009_/B vssd1 vssd1 vccd1 vccd1 _14143_/B1 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_215_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer72 _11461_/B vssd1 vssd1 vccd1 vccd1 _11542_/C1 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_42_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrebuffer83 _13066_/B vssd1 vssd1 vccd1 vccd1 _13206_/A2 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer94 _13537_/C vssd1 vssd1 vccd1 vccd1 _13598_/A sky130_fd_sc_hd__dlygate4sd1_1
XPHY_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_230_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11660_ _15389_/A _18520_/Q vssd1 vssd1 vccd1 vccd1 _11660_/Y sky130_fd_sc_hd__nor2_1
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10611_ _19811_/Q _10606_/A _10613_/A _10609_/X vssd1 vssd1 vccd1 vccd1 _19811_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11591_ _19573_/Q _19572_/Q _11591_/C vssd1 vssd1 vccd1 vccd1 _11591_/X sky130_fd_sc_hd__and3_1
XPHY_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12437__A _12487_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13330_ _18845_/Q vssd1 vssd1 vccd1 vccd1 _13468_/A sky130_fd_sc_hd__inv_2
XANTENNA__10073__B1 _10079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14339__B1 _14273_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11341__A _18986_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10542_ _10595_/A vssd1 vssd1 vccd1 vccd1 _10583_/A sky130_fd_sc_hd__clkbuf_2
XPHY_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17439__S _17512_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13261_ _13723_/A vssd1 vssd1 vccd1 vccd1 _15082_/A sky130_fd_sc_hd__clkbuf_2
X_10473_ _17697_/X _10471_/X _19822_/Q _10472_/X vssd1 vssd1 vccd1 vccd1 _19822_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_183_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12212_ _12228_/A vssd1 vssd1 vccd1 vccd1 _12212_/X sky130_fd_sc_hd__clkbuf_2
X_15000_ _18956_/Q vssd1 vssd1 vccd1 vccd1 _15000_/X sky130_fd_sc_hd__buf_2
XFILLER_136_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13192_ _13073_/A _13192_/A2 _13190_/Y _13182_/X vssd1 vssd1 vccd1 vccd1 _18901_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_135_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17923__S1 _19646_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12143_ _12150_/A vssd1 vssd1 vccd1 vccd1 _12143_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_150_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16951_ _17769_/X _18789_/Q _16957_/S vssd1 vssd1 vccd1 vccd1 _16951_/X sky130_fd_sc_hd__mux2_1
X_12074_ hold291/X vssd1 vssd1 vccd1 vccd1 _12074_/X sky130_fd_sc_hd__buf_2
XFILLER_49_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11025_ _19649_/Q _11025_/B vssd1 vssd1 vccd1 vccd1 _11026_/A sky130_fd_sc_hd__nand2_1
XANTENNA__15483__A _15512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15902_ _15902_/A vssd1 vssd1 vccd1 vccd1 _16494_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__17174__S _17541_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19670_ _19812_/CLK _19670_/D repeater225/X vssd1 vssd1 vccd1 vccd1 _19670_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_237_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16882_ _17473_/A0 _09943_/Y _17522_/S vssd1 vssd1 vccd1 vccd1 _16882_/X sky130_fd_sc_hd__mux2_1
X_18621_ _19867_/CLK hold212/X repeater262/X vssd1 vssd1 vccd1 vccd1 _18621_/Q sky130_fd_sc_hd__dfrtp_1
X_15833_ _15822_/Y _15864_/B _15825_/Y _15828_/X _15832_/X vssd1 vssd1 vccd1 vccd1
+ _15833_/X sky130_fd_sc_hd__o221a_1
XFILLER_64_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18552_ _19810_/CLK _18552_/D repeater224/X vssd1 vssd1 vccd1 vccd1 _18552_/Q sky130_fd_sc_hd__dfrtp_1
X_15764_ _18880_/Q vssd1 vssd1 vccd1 vccd1 _15764_/Y sky130_fd_sc_hd__inv_2
X_12976_ _12887_/A _12975_/A _18944_/Q _12975_/Y _12958_/X vssd1 vssd1 vccd1 vccd1
+ _18944_/D sky130_fd_sc_hd__o221a_1
XFILLER_18_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17503_ _17502_/X _17899_/X _17568_/S vssd1 vssd1 vccd1 vccd1 _17503_/X sky130_fd_sc_hd__mux2_2
XFILLER_33_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14715_ _18218_/Q _14700_/A _14626_/X _14701_/A vssd1 vssd1 vccd1 vccd1 _18218_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19812__RESET_B repeater222/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18483_ _19545_/CLK _18483_/D repeater225/X vssd1 vssd1 vccd1 vccd1 _18483_/Q sky130_fd_sc_hd__dfrtp_1
X_11927_ _19401_/Q _11891_/A _11926_/X _11892_/A vssd1 vssd1 vccd1 vccd1 _19401_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16567__A1 _17146_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15695_ _15702_/A _15695_/B vssd1 vssd1 vccd1 vccd1 _15695_/Y sky130_fd_sc_hd__nor2_1
XPHY_4570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17434_ _16096_/Y _16095_/Y _17564_/S vssd1 vssd1 vccd1 vccd1 _17434_/X sky130_fd_sc_hd__mux2_1
XFILLER_220_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14646_ _18257_/Q _14643_/X _09168_/X _14645_/X vssd1 vssd1 vccd1 vccd1 _18257_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_205_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11858_ _13641_/A _19329_/Q vssd1 vssd1 vccd1 vccd1 _12058_/B sky130_fd_sc_hd__or2_2
XFILLER_82_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10809_ _10809_/A vssd1 vssd1 vccd1 vccd1 _10810_/A sky130_fd_sc_hd__inv_2
X_17365_ _17364_/X _13891_/Y _17545_/S vssd1 vssd1 vccd1 vccd1 _17365_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13250__B1 _12541_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14577_ _18295_/Q _14572_/X _14537_/X _14574_/X vssd1 vssd1 vccd1 vccd1 _18295_/D
+ sky130_fd_sc_hd__a22o_1
X_11789_ _19469_/Q _11784_/X _09021_/X _11787_/X vssd1 vssd1 vccd1 vccd1 _19469_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_13_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19104_ _19109_/CLK _19104_/D hold361/X vssd1 vssd1 vccd1 vccd1 _19104_/Q sky130_fd_sc_hd__dfrtp_4
X_16316_ _19820_/Q vssd1 vssd1 vccd1 vccd1 _16316_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13528_ _13528_/A _13528_/B vssd1 vssd1 vccd1 vccd1 _13610_/A sky130_fd_sc_hd__or2_1
X_17296_ _17295_/X _13069_/A _17542_/S vssd1 vssd1 vccd1 vccd1 _17296_/X sky130_fd_sc_hd__mux2_1
XFILLER_185_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12066__B _12187_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19035_ _19157_/CLK _19035_/D repeater267/X vssd1 vssd1 vccd1 vccd1 _19035_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17349__S _17517_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16247_ _16509_/A vssd1 vssd1 vccd1 vccd1 _16595_/A sky130_fd_sc_hd__inv_2
X_13459_ _13459_/A vssd1 vssd1 vccd1 vccd1 _13459_/Y sky130_fd_sc_hd__inv_2
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput104 _16151_/Y vssd1 vssd1 vccd1 vccd1 HRDATA[3] sky130_fd_sc_hd__clkbuf_2
XANTENNA__14750__B1 _14749_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput115 _16755_/LO vssd1 vssd1 vccd1 vccd1 IRQ[12] sky130_fd_sc_hd__clkbuf_2
X_16178_ _18094_/Q vssd1 vssd1 vccd1 vccd1 _16178_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18765__RESET_B repeater196/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput126 _15778_/X vssd1 vssd1 vccd1 vccd1 IRQ[8] sky130_fd_sc_hd__clkbuf_2
Xoutput137 _18671_/Q vssd1 vssd1 vccd1 vccd1 pwm_S7 sky130_fd_sc_hd__clkbuf_2
XANTENNA__17914__S1 _19634_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15129_ _17972_/Q _15122_/X _14931_/X _15124_/X vssd1 vssd1 vccd1 vccd1 _17972_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_126_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19937_ _19937_/CLK _19937_/D repeater189/X vssd1 vssd1 vccd1 vccd1 _19937_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__15393__A _15419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17084__S _17546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19868_ _20059_/CLK _19868_/D repeater199/X vssd1 vssd1 vccd1 vccd1 _19868_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_229_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19966__CLK _19976_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09621_ _10029_/B vssd1 vssd1 vccd1 vccd1 _10079_/A sky130_fd_sc_hd__clkbuf_4
X_18819_ _18827_/CLK _18819_/D repeater231/X vssd1 vssd1 vccd1 vccd1 _18819_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_28_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19799_ _19808_/CLK _19799_/D repeater222/X vssd1 vssd1 vccd1 vccd1 _19799_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_244_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_237_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09552_ _19321_/Q vssd1 vssd1 vccd1 vccd1 _09552_/Y sky130_fd_sc_hd__inv_2
XFILLER_102_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09483_ _09483_/A _09589_/A vssd1 vssd1 vccd1 vccd1 _09484_/B sky130_fd_sc_hd__or2_2
XANTENNA__19553__RESET_B repeater274/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16558__A1 _17163_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17850__S0 _17913_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15230__A1 _15205_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12257__A _12257_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16671__B _16718_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17259__S _17493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14741__B1 _14691_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17905__S1 _18759_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_219_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20008_ _20013_/CLK _20008_/D repeater241/X vssd1 vssd1 vccd1 vccd1 _20008_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_47_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09819_ _19967_/Q vssd1 vssd1 vccd1 vccd1 _09875_/A sky130_fd_sc_hd__inv_2
XFILLER_247_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12830_ _18828_/Q vssd1 vssd1 vccd1 vccd1 _13551_/A sky130_fd_sc_hd__inv_2
XFILLER_46_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09279__A2 _09270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12761_ _19240_/Q vssd1 vssd1 vccd1 vccd1 _12761_/Y sky130_fd_sc_hd__inv_2
XPHY_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14500_ _18339_/Q _14492_/A _12731_/X _14493_/A vssd1 vssd1 vccd1 vccd1 _18339_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11712_ _15858_/A _11708_/X _16925_/X _16950_/S vssd1 vssd1 vccd1 vccd1 hold219/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_202_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17841__S0 _17913_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12692_ _12699_/A vssd1 vssd1 vccd1 vccd1 _12692_/X sky130_fd_sc_hd__clkbuf_2
X_15480_ _18565_/Q vssd1 vssd1 vccd1 vccd1 _15480_/Y sky130_fd_sc_hd__inv_2
XFILLER_199_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14431_ _18381_/Q _14424_/X _14417_/X _14426_/X vssd1 vssd1 vccd1 vccd1 _18381_/D
+ sky130_fd_sc_hd__a22o_1
X_11643_ _11548_/B _11642_/A _19548_/Q _11645_/A _11588_/X vssd1 vssd1 vccd1 vccd1
+ _19548_/D sky130_fd_sc_hd__o221a_1
XPHY_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17150_ _15963_/X _09514_/Y _17534_/S vssd1 vssd1 vccd1 vccd1 _17150_/X sky130_fd_sc_hd__mux2_1
XPHY_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14362_ _18421_/Q _14349_/X _14326_/X _14353_/X vssd1 vssd1 vccd1 vccd1 _18421_/D
+ sky130_fd_sc_hd__a22o_1
X_11574_ _11574_/A _11612_/A vssd1 vssd1 vccd1 vccd1 _11575_/B sky130_fd_sc_hd__or2_2
XANTENNA__14980__B1 hold247/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16581__B _16581_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput17 HADDR[24] vssd1 vssd1 vccd1 vccd1 input17/X sky130_fd_sc_hd__buf_1
XFILLER_6_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput28 input28/A vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__buf_1
XPHY_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16101_ _18269_/Q vssd1 vssd1 vccd1 vccd1 _16101_/Y sky130_fd_sc_hd__inv_2
X_10525_ _10734_/A _10525_/B _19535_/Q _10525_/D vssd1 vssd1 vccd1 vccd1 _11652_/B
+ sky130_fd_sc_hd__nor4_2
X_13313_ _18852_/Q vssd1 vssd1 vccd1 vccd1 _13430_/A sky130_fd_sc_hd__clkinvlp_4
Xinput39 input39/A vssd1 vssd1 vccd1 vccd1 input39/X sky130_fd_sc_hd__buf_1
XANTENNA__17169__S _17318_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14293_ _18455_/Q _14288_/X _14279_/X _14290_/X vssd1 vssd1 vccd1 vccd1 _18455_/D
+ sky130_fd_sc_hd__a22o_1
X_17081_ _17080_/X _15475_/A _17524_/S vssd1 vssd1 vccd1 vccd1 _17081_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_183_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13244_ _15419_/A _13241_/X _12596_/X _13243_/X vssd1 vssd1 vccd1 vccd1 _18879_/D
+ sky130_fd_sc_hd__a22o_1
X_16032_ _18236_/Q vssd1 vssd1 vccd1 vccd1 _16032_/Y sky130_fd_sc_hd__inv_2
X_10456_ _19828_/Q _10450_/X _10423_/X _10452_/X vssd1 vssd1 vccd1 vccd1 _19828_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_6_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_14_0_HCLK_A clkbuf_3_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13175_ _13175_/A vssd1 vssd1 vccd1 vccd1 _13175_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16801__S _17534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10387_ _19852_/Q _10335_/B _10319_/A _08964_/X vssd1 vssd1 vccd1 vccd1 _19852_/D
+ sky130_fd_sc_hd__o22a_1
XANTENNA__18863__CLK _18866_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19989__CLK _19992_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12126_ _19297_/Q _12121_/X _11920_/X _12122_/X vssd1 vssd1 vccd1 vccd1 _19297_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_69_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17983_ _20124_/CLK _17983_/D vssd1 vssd1 vccd1 vccd1 _17983_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_238_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19722_ _19795_/CLK _19722_/D repeater219/X vssd1 vssd1 vccd1 vccd1 _19722_/Q sky130_fd_sc_hd__dfrtp_1
X_12057_ _13641_/A _12056_/A _11853_/A _12056_/Y vssd1 vssd1 vccd1 vccd1 _19330_/D
+ sky130_fd_sc_hd__a22o_1
X_16934_ _19478_/Q hold186/X _16946_/S vssd1 vssd1 vccd1 vccd1 _16934_/X sky130_fd_sc_hd__mux2_1
XFILLER_78_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11008_ _11008_/A vssd1 vssd1 vccd1 vccd1 _19658_/D sky130_fd_sc_hd__inv_2
X_19653_ _19855_/CLK _19653_/D repeater264/X vssd1 vssd1 vccd1 vccd1 _19653_/Q sky130_fd_sc_hd__dfrtp_4
X_16865_ _16864_/X _09697_/Y _17523_/S vssd1 vssd1 vccd1 vccd1 _16865_/X sky130_fd_sc_hd__mux2_1
XFILLER_226_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11864__A4 _10954_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18604_ _19041_/CLK _18604_/D repeater266/X vssd1 vssd1 vccd1 vccd1 _18604_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_219_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15816_ _18098_/Q vssd1 vssd1 vccd1 vccd1 _15816_/Y sky130_fd_sc_hd__inv_2
X_19584_ _19591_/CLK _19584_/D hold361/X vssd1 vssd1 vccd1 vccd1 _19584_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__10150__A _12257_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16796_ _15963_/X _12774_/Y _17534_/S vssd1 vssd1 vccd1 vccd1 _16796_/X sky130_fd_sc_hd__mux2_1
XFILLER_92_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15996__C1 _15995_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18535_ _19822_/CLK _18535_/D repeater228/X vssd1 vssd1 vccd1 vccd1 _18535_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_93_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15747_ _19671_/Q _19670_/Q _15747_/C vssd1 vssd1 vccd1 vccd1 _15747_/X sky130_fd_sc_hd__and3_1
XFILLER_34_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12959_ _18950_/Q _12892_/Y _12893_/Y _12892_/A _12958_/X vssd1 vssd1 vccd1 vccd1
+ _18950_/D sky130_fd_sc_hd__o221a_1
XANTENNA__18243__CLK _19847_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17832__S0 _17918_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18466_ _19630_/CLK _18466_/D vssd1 vssd1 vccd1 vccd1 _18466_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15678_ _18612_/Q _15678_/B vssd1 vssd1 vccd1 vccd1 _15678_/X sky130_fd_sc_hd__and2_1
XFILLER_21_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17417_ _17416_/X _13531_/A _17536_/S vssd1 vssd1 vccd1 vccd1 _17417_/X sky130_fd_sc_hd__mux2_2
X_14629_ _14857_/A _14629_/B _15157_/C vssd1 vssd1 vccd1 vccd1 _14631_/A sky130_fd_sc_hd__or3_4
X_18397_ _18416_/CLK _18397_/D vssd1 vssd1 vccd1 vccd1 _18397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_193_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17348_ _17347_/X _15598_/A _17474_/S vssd1 vssd1 vccd1 vccd1 _17348_/X sky130_fd_sc_hd__mux2_1
XANTENNA__14971__B1 _14812_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17079__S _17542_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17279_ _17278_/X _15622_/A _17318_/S vssd1 vssd1 vccd1 vccd1 _17279_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19018_ _19115_/CLK _19018_/D hold353/X vssd1 vssd1 vccd1 vccd1 _19018_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_228_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17899__S0 _18760_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08983_ _10132_/B _08983_/B vssd1 vssd1 vccd1 vccd1 _08983_/X sky130_fd_sc_hd__or2_1
XFILLER_244_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12540__A hold336/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_8_HCLK_A clkbuf_4_2_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_119_HCLK clkbuf_opt_0_HCLK/A vssd1 vssd1 vccd1 vccd1 _19591_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_28_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19734__RESET_B repeater207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09604_ _09604_/A _09604_/B _09604_/C vssd1 vssd1 vccd1 vccd1 _20014_/D sky130_fd_sc_hd__nor3_1
XANTENNA__17542__S _17542_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16666__B _16668_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09535_ _19317_/Q vssd1 vssd1 vccd1 vccd1 _09535_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17728__A0 _17936_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09466_ _09466_/A _09618_/A vssd1 vssd1 vccd1 vccd1 _09467_/B sky130_fd_sc_hd__or2_2
XPHY_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17823__S0 _17918_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_240_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09397_ _19913_/Q _19373_/Q _10085_/A _09396_/Y vssd1 vssd1 vccd1 vccd1 _09397_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16682__A _16682_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_240_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09969__B1 _09968_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09433__A2 _09431_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18687__RESET_B hold359/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16703__A1 _16827_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10310_ _18615_/Q _18614_/Q _10310_/C _15678_/B vssd1 vssd1 vccd1 vccd1 _15693_/A
+ sky130_fd_sc_hd__or4_4
XANTENNA__13517__A1 _18759_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11290_ _11473_/A _19007_/Q _11480_/A _19014_/Q vssd1 vssd1 vccd1 vccd1 _11290_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_3_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17717__S _18546_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10241_ _19655_/Q vssd1 vssd1 vccd1 vccd1 _10956_/C sky130_fd_sc_hd__inv_2
XFILLER_106_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10172_ _19884_/Q _10166_/X _09086_/X _10168_/X vssd1 vssd1 vccd1 vccd1 _19884_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_121_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10751__A1 _19756_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12450__A _12457_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14980_ _18065_/Q _14976_/X hold247/X _14979_/X vssd1 vssd1 vccd1 vccd1 _18065_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_120_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13931_ _13909_/B _13823_/B _13929_/Y _13927_/X vssd1 vssd1 vccd1 vccd1 _18724_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_87_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_208_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11700__B1 _10870_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11066__A _19633_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17452__S _17522_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16650_ _19461_/Q _16673_/B vssd1 vssd1 vccd1 vccd1 _16650_/Y sky130_fd_sc_hd__nand2_1
XFILLER_74_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13862_ _13858_/Y _18706_/Q _13859_/Y _18731_/Q _13861_/X vssd1 vssd1 vccd1 vccd1
+ _13867_/C sky130_fd_sc_hd__o221a_1
XFILLER_234_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15601_ _15601_/A vssd1 vssd1 vccd1 vccd1 _15606_/B sky130_fd_sc_hd__inv_2
X_12813_ _19239_/Q _13539_/A _19247_/Q _13547_/A vssd1 vssd1 vccd1 vccd1 _12813_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_90_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16581_ _16572_/X _16581_/B _16581_/C vssd1 vssd1 vccd1 vccd1 _16581_/Y sky130_fd_sc_hd__nand3b_4
XFILLER_16_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_234_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13793_ _18719_/Q vssd1 vssd1 vccd1 vccd1 _13911_/A sky130_fd_sc_hd__inv_2
XFILLER_43_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18320_ _18431_/CLK _18320_/D vssd1 vssd1 vccd1 vccd1 _18320_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15532_ _15535_/A _15532_/B vssd1 vssd1 vccd1 vccd1 _15532_/Y sky130_fd_sc_hd__nor2_1
X_12744_ _19246_/Q _13546_/A _16546_/A _18818_/Q vssd1 vssd1 vccd1 vccd1 _12744_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_15_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17814__S0 _18751_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12609__B _15863_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18251_ _18268_/CLK _18251_/D vssd1 vssd1 vccd1 vccd1 _18251_/Q sky130_fd_sc_hd__dfxtp_1
X_15463_ _15463_/A _15463_/B vssd1 vssd1 vccd1 vccd1 _15463_/Y sky130_fd_sc_hd__nor2_1
XPHY_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12675_ _18983_/Q _12670_/X hold296/X _12671_/X vssd1 vssd1 vccd1 vccd1 _18983_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17202_ _17201_/X _13543_/A _17536_/S vssd1 vssd1 vccd1 vccd1 _17202_/X sky130_fd_sc_hd__mux2_1
XPHY_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14414_ _18391_/Q _14409_/X _14359_/X _14411_/X vssd1 vssd1 vccd1 vccd1 _18391_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11626_ _11626_/A _11626_/B vssd1 vssd1 vccd1 vccd1 _11626_/Y sky130_fd_sc_hd__nor2_1
X_18182_ _18198_/CLK _18182_/D vssd1 vssd1 vccd1 vccd1 _18182_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15394_ _15402_/A _17583_/X vssd1 vssd1 vccd1 vccd1 _18529_/D sky130_fd_sc_hd__and2_1
XPHY_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17133_ _17486_/A0 _09897_/Y _17543_/S vssd1 vssd1 vccd1 vccd1 _17133_/X sky130_fd_sc_hd__mux2_1
X_14345_ _18427_/Q _14337_/A _14312_/X _14338_/A vssd1 vssd1 vccd1 vccd1 _18427_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_128_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11557_ _19570_/Q vssd1 vssd1 vccd1 vccd1 _11583_/A sky130_fd_sc_hd__inv_2
XPHY_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10508_ _10508_/A _10508_/B _10508_/C _10514_/D vssd1 vssd1 vccd1 vccd1 _15270_/A
+ sky130_fd_sc_hd__nor4_2
XFILLER_6_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17064_ _16621_/Y _19421_/Q _17541_/S vssd1 vssd1 vccd1 vccd1 _17064_/X sky130_fd_sc_hd__mux2_1
X_11488_ _11488_/A _11488_/B vssd1 vssd1 vccd1 vccd1 _11489_/A sky130_fd_sc_hd__or2_1
XANTENNA_output99_A _16715_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14276_ _18465_/Q _14272_/X _14273_/X _14275_/X vssd1 vssd1 vccd1 vccd1 _18465_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_195_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16015_ _18164_/Q vssd1 vssd1 vccd1 vccd1 _16015_/Y sky130_fd_sc_hd__inv_2
X_13227_ _18540_/Q _13227_/B vssd1 vssd1 vccd1 vccd1 _13228_/B sky130_fd_sc_hd__or2_1
X_10439_ _19838_/Q _10433_/X _09067_/X _10435_/X vssd1 vssd1 vccd1 vccd1 _19838_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_170_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13158_ _13156_/Y _18888_/Q _19174_/Q _13075_/A _13157_/X vssd1 vssd1 vccd1 vccd1
+ _13159_/D sky130_fd_sc_hd__o221a_1
X_12109_ _19310_/Q _12106_/X _12107_/X _12108_/X vssd1 vssd1 vccd1 vccd1 _19310_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_69_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17966_ _19842_/CLK _17966_/D vssd1 vssd1 vccd1 vccd1 _17966_/Q sky130_fd_sc_hd__dfxtp_1
X_13089_ _13089_/A _13089_/B vssd1 vssd1 vccd1 vccd1 _13090_/A sky130_fd_sc_hd__or2_4
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16917_ _15963_/X _09529_/Y _17534_/S vssd1 vssd1 vccd1 vccd1 _16917_/X sky130_fd_sc_hd__mux2_1
X_19705_ _19720_/CLK _19705_/D repeater202/X vssd1 vssd1 vccd1 vccd1 _19705_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_77_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17897_ _15948_/Y _15949_/Y _15950_/Y _15951_/Y _17908_/S0 _18759_/Q vssd1 vssd1
+ vccd1 vccd1 _17897_/X sky130_fd_sc_hd__mux4_1
XANTENNA__17362__S _17488_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16848_ _15768_/Y _14172_/Y _17546_/S vssd1 vssd1 vccd1 vccd1 _16848_/X sky130_fd_sc_hd__mux2_1
X_19636_ _19851_/CLK _19636_/D repeater258/X vssd1 vssd1 vccd1 vccd1 _19636_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_226_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19567_ _19576_/CLK _19567_/D repeater282/X vssd1 vssd1 vccd1 vccd1 _19567_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18759__CLK _20123_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16779_ _16722_/Y _15565_/Y _17513_/S vssd1 vssd1 vccd1 vccd1 _16779_/X sky130_fd_sc_hd__mux2_1
XFILLER_241_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09320_ _20044_/Q vssd1 vssd1 vccd1 vccd1 _09320_/Y sky130_fd_sc_hd__inv_2
X_18518_ _20049_/CLK _18518_/D repeater208/X vssd1 vssd1 vccd1 vccd1 _18518_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17805__S0 _17918_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_230_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19498_ _20036_/CLK _19498_/D repeater194/X vssd1 vssd1 vccd1 vccd1 _19498_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_61_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09251_ _20060_/Q _20061_/Q _09253_/S vssd1 vssd1 vccd1 vccd1 _20061_/D sky130_fd_sc_hd__mux2_1
X_18449_ _19855_/CLK _18449_/D vssd1 vssd1 vccd1 vccd1 _18449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_222_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09182_ _20075_/Q vssd1 vssd1 vccd1 vccd1 _14713_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__18641__SET_B repeater204/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12535__A hold332/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15846__A _15846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17537__S _17537_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19986__RESET_B repeater193/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_144_HCLK_A clkbuf_4_1_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17110__A1 _12905_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08966_ _18778_/Q vssd1 vssd1 vccd1 vccd1 _08966_/Y sky130_fd_sc_hd__inv_2
XFILLER_102_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13683__B1 _13682_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12486__B2 _12458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17272__S _17488_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_216_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19684__CLK _19780_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_231_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09518_ _19305_/Q vssd1 vssd1 vccd1 vccd1 _09518_/Y sky130_fd_sc_hd__inv_2
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10790_ _19739_/Q _18653_/Q _10786_/Y _10788_/Y _10789_/Y vssd1 vssd1 vccd1 vccd1
+ _19739_/D sky130_fd_sc_hd__a32o_1
XFILLER_140_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18868__RESET_B repeater217/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15188__B1 _10715_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09449_ _19371_/Q vssd1 vssd1 vccd1 vccd1 _09449_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12460_ _19113_/Q _12457_/X _12404_/X _12458_/X vssd1 vssd1 vccd1 vccd1 _19113_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_130_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11411_ _11549_/A _19126_/Q _11574_/A _19141_/Q _11410_/X vssd1 vssd1 vccd1 vccd1
+ _11412_/D sky130_fd_sc_hd__o221a_1
X_12391_ _19152_/Q _12388_/X _12389_/X _12390_/X vssd1 vssd1 vccd1 vccd1 _19152_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09738__B _09813_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09811__C1 _09759_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11342_ _11483_/A _18985_/Q _11469_/A _18971_/Q vssd1 vssd1 vccd1 vccd1 _11342_/X
+ sky130_fd_sc_hd__o22a_1
X_14130_ _18685_/Q _14129_/Y _14116_/X _14130_/C1 vssd1 vssd1 vccd1 vccd1 _18685_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_125_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17447__S _17529_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11273_ _11469_/A _19003_/Q _19592_/Q _16542_/A _11272_/X vssd1 vssd1 vccd1 vccd1
+ _11299_/C sky130_fd_sc_hd__o221a_1
X_14061_ _19087_/Q vssd1 vssd1 vccd1 vccd1 _14061_/Y sky130_fd_sc_hd__inv_2
XFILLER_140_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12174__B1 _11981_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13012_ _18928_/Q _13011_/Y _13008_/B _12980_/X vssd1 vssd1 vccd1 vccd1 _18928_/D
+ sky130_fd_sc_hd__o211a_1
X_10224_ _10956_/A vssd1 vssd1 vccd1 vccd1 _10224_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__19656__RESET_B repeater270/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20041__CLK _20051_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10724__A1 _19771_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11921__B1 _11920_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17820_ _18334_/Q _18214_/Q _18206_/Q _18198_/Q _17918_/S0 _18750_/Q vssd1 vssd1
+ vccd1 vccd1 _17820_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10155_ _10155_/A vssd1 vssd1 vccd1 vccd1 _10156_/A sky130_fd_sc_hd__inv_2
XANTENNA__12180__A _12313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16860__A0 _17473_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17751_ _18482_/Q _15298_/X _18508_/Q vssd1 vssd1 vccd1 vccd1 _17751_/X sky130_fd_sc_hd__mux2_1
XFILLER_121_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_66_HCLK_A clkbuf_opt_3_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10086_ _10086_/A _10086_/B vssd1 vssd1 vccd1 vccd1 _10091_/A sky130_fd_sc_hd__or2_1
X_14963_ _14990_/A _14963_/B _15058_/C vssd1 vssd1 vccd1 vccd1 _14965_/A sky130_fd_sc_hd__or3_4
XANTENNA_output137_A _18671_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17182__S _17546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16702_ _17048_/X _16683_/X _16806_/X _16684_/X _16701_/X vssd1 vssd1 vccd1 vccd1
+ _16705_/B sky130_fd_sc_hd__o221a_4
XANTENNA__09342__A1 _20036_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13914_ _13914_/A _13914_/B _13914_/C _13913_/X vssd1 vssd1 vccd1 vccd1 _13914_/X
+ sky130_fd_sc_hd__or4b_4
XFILLER_208_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17682_ _15503_/Y _19453_/Q _17683_/S vssd1 vssd1 vccd1 vccd1 _18570_/D sky130_fd_sc_hd__mux2_1
XFILLER_235_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14894_ _15145_/A vssd1 vssd1 vccd1 vccd1 _15109_/A sky130_fd_sc_hd__buf_1
XANTENNA__09893__A2 _19360_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19421_ _19997_/CLK _19421_/D repeater185/X vssd1 vssd1 vccd1 vccd1 _19421_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_90_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16633_ _16633_/A vssd1 vssd1 vccd1 vccd1 _16633_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_74_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13845_ _19203_/Q vssd1 vssd1 vccd1 vccd1 _13845_/Y sky130_fd_sc_hd__inv_2
XFILLER_223_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19352_ _19352_/CLK _19352_/D hold373/X vssd1 vssd1 vccd1 vccd1 _19352_/Q sky130_fd_sc_hd__dfrtp_1
X_16564_ _17193_/X _16687_/A _17184_/X _16683_/A vssd1 vssd1 vccd1 vccd1 _16564_/X
+ sky130_fd_sc_hd__o22a_1
X_13776_ _19190_/Q vssd1 vssd1 vccd1 vccd1 _13776_/Y sky130_fd_sc_hd__inv_2
XFILLER_200_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10988_ _19663_/Q _10988_/B vssd1 vssd1 vccd1 vccd1 _10988_/Y sky130_fd_sc_hd__nor2_1
XFILLER_204_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18303_ _18431_/CLK _18303_/D vssd1 vssd1 vccd1 vccd1 _18303_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15515_ _18573_/Q _15518_/C _15514_/Y _15510_/Y vssd1 vssd1 vccd1 vccd1 _15516_/B
+ sky130_fd_sc_hd__o22a_1
X_12727_ _14814_/A _12710_/A _12726_/X _12711_/A vssd1 vssd1 vccd1 vccd1 _18954_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__15179__B1 _09339_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19283_ _19283_/CLK _19283_/D repeater212/X vssd1 vssd1 vccd1 vccd1 _19283_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_176_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16495_ _17233_/X _16687_/A _17225_/X _16683_/A vssd1 vssd1 vccd1 vccd1 _16495_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_204_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18234_ _20076_/CLK _18234_/D vssd1 vssd1 vccd1 vccd1 _18234_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15446_ _15479_/A _18556_/Q vssd1 vssd1 vccd1 vccd1 _15446_/Y sky130_fd_sc_hd__nor2_1
XPHY_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12658_ _18992_/Q _12629_/A _12543_/X _12630_/A vssd1 vssd1 vccd1 vccd1 _18992_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11609_ _11609_/A vssd1 vssd1 vccd1 vccd1 _11609_/Y sky130_fd_sc_hd__inv_2
X_18165_ _18165_/CLK _18165_/D vssd1 vssd1 vccd1 vccd1 _18165_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__19407__CLK _19984_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15377_ _19793_/Q _10653_/B _10654_/B vssd1 vssd1 vccd1 vccd1 _15377_/X sky130_fd_sc_hd__a21bo_1
X_12589_ _19037_/Q _12583_/X hold270/X _12584_/X vssd1 vssd1 vccd1 vccd1 _19037_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17116_ _17115_/X _15504_/Y _17513_/S vssd1 vssd1 vccd1 vccd1 _17116_/X sky130_fd_sc_hd__mux2_1
XFILLER_172_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14328_ hold264/X vssd1 vssd1 vccd1 vccd1 _14727_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_116_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_opt_1_HCLK clkbuf_opt_1_HCLK/A vssd1 vssd1 vccd1 vccd1 _18642_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_156_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18096_ _20090_/CLK _18096_/D vssd1 vssd1 vccd1 vccd1 _18096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17357__S _17534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17047_ _17046_/X _14042_/Y _17490_/S vssd1 vssd1 vccd1 vccd1 _17047_/X sky130_fd_sc_hd__mux2_2
X_14259_ _14259_/A vssd1 vssd1 vccd1 vccd1 _14260_/A sky130_fd_sc_hd__inv_2
XFILLER_143_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11912__B1 _11911_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12090__A hold296/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19326__RESET_B repeater241/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18998_ _19208_/CLK _18998_/D repeater249/X vssd1 vssd1 vccd1 vccd1 _18998_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_140_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16851__A0 _15963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater201 repeater202/X vssd1 vssd1 vccd1 vccd1 repeater201/X sky130_fd_sc_hd__clkbuf_8
Xrepeater212 repeater216/X vssd1 vssd1 vccd1 vccd1 repeater212/X sky130_fd_sc_hd__buf_8
Xrepeater223 repeater225/X vssd1 vssd1 vccd1 vccd1 repeater223/X sky130_fd_sc_hd__buf_6
XFILLER_245_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17949_ _18137_/CLK _17949_/D vssd1 vssd1 vccd1 vccd1 _17949_/Q sky130_fd_sc_hd__dfxtp_1
Xrepeater234 repeater235/X vssd1 vssd1 vccd1 vccd1 repeater234/X sky130_fd_sc_hd__buf_8
XANTENNA__17092__S _17488_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrepeater245 hold373/A vssd1 vssd1 vccd1 vccd1 repeater245/X sky130_fd_sc_hd__clkbuf_8
XFILLER_226_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater256 repeater260/X vssd1 vssd1 vccd1 vccd1 repeater256/X sky130_fd_sc_hd__buf_6
XFILLER_238_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater267 repeater268/X vssd1 vssd1 vccd1 vccd1 repeater267/X sky130_fd_sc_hd__buf_6
Xrepeater278 hold343/X vssd1 vssd1 vccd1 vccd1 hold346/A sky130_fd_sc_hd__buf_6
XFILLER_93_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19619_ _19927_/CLK _19619_/D repeater230/X vssd1 vssd1 vccd1 vccd1 _19619_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_38_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09303_ _18659_/Q _09303_/B vssd1 vssd1 vccd1 vccd1 _09304_/A sky130_fd_sc_hd__nand2_1
XFILLER_61_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09234_ _15711_/A vssd1 vssd1 vccd1 vccd1 _09234_/Y sky130_fd_sc_hd__inv_2
XFILLER_166_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09165_ _09165_/A vssd1 vssd1 vccd1 vccd1 _09165_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_181_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09096_ hold332/X vssd1 vssd1 vccd1 vccd1 _14793_/A sky130_fd_sc_hd__buf_4
XANTENNA__17331__A1 _12933_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17267__S _17543_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12156__B1 _12104_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15893__A1 _17536_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15893__B2 _15845_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17095__A0 _17094_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11903__B1 _09064_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09998_ _09998_/A vssd1 vssd1 vccd1 vccd1 _09998_/Y sky130_fd_sc_hd__inv_2
XFILLER_237_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16842__A0 _15768_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12459__A1 _19114_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08949_ _10327_/A _18781_/Q _19852_/Q _08945_/Y _08948_/X vssd1 vssd1 vccd1 vccd1
+ _08969_/A sky130_fd_sc_hd__o221a_1
XFILLER_69_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11960_ _19384_/Q _11955_/X _09049_/X _11956_/X vssd1 vssd1 vccd1 vccd1 _19384_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_57_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10911_ _18511_/Q vssd1 vssd1 vccd1 vccd1 _10912_/C sky130_fd_sc_hd__inv_2
XFILLER_44_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_233_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11891_ _11891_/A vssd1 vssd1 vccd1 vccd1 _11891_/X sky130_fd_sc_hd__buf_1
XFILLER_72_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17730__S _18508_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13630_ _13630_/A _13630_/B vssd1 vssd1 vccd1 vccd1 _13630_/X sky130_fd_sc_hd__or2_1
XANTENNA__09088__B1 _09086_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10842_ _10842_/A _14245_/D vssd1 vssd1 vccd1 vccd1 _10844_/A sky130_fd_sc_hd__or2_4
XANTENNA__10890__B1 _10868_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_232_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13561_ _18835_/Q _13558_/Y _12829_/Y _13558_/A _13560_/X vssd1 vssd1 vccd1 vccd1
+ _18835_/D sky130_fd_sc_hd__o221a_1
XANTENNA__12631__A1 _19013_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10773_ _10773_/A vssd1 vssd1 vccd1 vccd1 _10774_/A sky130_fd_sc_hd__inv_2
XFILLER_201_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15300_ _20046_/Q vssd1 vssd1 vccd1 vccd1 _15300_/Y sky130_fd_sc_hd__inv_2
X_12512_ _12528_/A vssd1 vssd1 vccd1 vccd1 _12512_/X sky130_fd_sc_hd__buf_1
XFILLER_201_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11998__B _15769_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16280_ _18255_/Q vssd1 vssd1 vccd1 vccd1 _16280_/Y sky130_fd_sc_hd__inv_2
XFILLER_197_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13492_ _15858_/A _15858_/B _15190_/A _15909_/A vssd1 vssd1 vccd1 vccd1 _15195_/A
+ sky130_fd_sc_hd__or4_4
XANTENNA__17570__A1 _19773_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15231_ _15231_/A vssd1 vssd1 vccd1 vccd1 _18640_/D sky130_fd_sc_hd__inv_2
X_12443_ _12479_/A vssd1 vssd1 vccd1 vccd1 _12458_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_8_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11198__B2 _11192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12395__B1 _12394_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15162_ _17951_/Q _15158_/X _14703_/A _15160_/X vssd1 vssd1 vccd1 vccd1 _17951_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12374_ _12400_/A vssd1 vssd1 vccd1 vccd1 _12374_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__19837__RESET_B repeater272/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14113_ _18695_/Q _14111_/Y _14113_/B1 _14112_/X vssd1 vssd1 vccd1 vccd1 _18695_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__17177__S _17541_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11325_ _18988_/Q vssd1 vssd1 vccd1 vccd1 _11325_/Y sky130_fd_sc_hd__inv_2
X_15093_ _17994_/Q _15084_/A _09255_/X _15085_/A vssd1 vssd1 vccd1 vccd1 _17994_/D
+ sky130_fd_sc_hd__a22o_1
X_19970_ _19970_/CLK _19970_/D hold370/X vssd1 vssd1 vccd1 vccd1 _19970_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_4_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12147__B1 _12088_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14044_ _14043_/Y _18701_/Q _19085_/Q _14026_/A vssd1 vssd1 vccd1 vccd1 _14044_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_4_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11256_ _19000_/Q vssd1 vssd1 vccd1 vccd1 _16466_/A sky130_fd_sc_hd__inv_2
X_18921_ _18947_/CLK _18921_/D repeater211/X vssd1 vssd1 vccd1 vccd1 _18921_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__19490__RESET_B repeater260/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10207_ _19667_/Q vssd1 vssd1 vccd1 vccd1 _10967_/A sky130_fd_sc_hd__inv_2
XFILLER_68_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18852_ _18852_/CLK _18852_/D repeater232/X vssd1 vssd1 vccd1 vccd1 _18852_/Q sky130_fd_sc_hd__dfrtp_2
X_11187_ _17711_/X _11184_/X _19620_/Q _11185_/X vssd1 vssd1 vccd1 vccd1 _19620_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_repeater202_A repeater203/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11370__B2 _19143_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17803_ _18474_/Q _18450_/Q _18458_/Q _18058_/Q _17918_/S0 _18750_/Q vssd1 vssd1
+ vccd1 vccd1 _17803_/X sky130_fd_sc_hd__mux4_1
X_10138_ _10138_/A vssd1 vssd1 vccd1 vccd1 _10138_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_227_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18783_ _19865_/CLK _18783_/D repeater265/X vssd1 vssd1 vccd1 vccd1 _18783_/Q sky130_fd_sc_hd__dfrtp_1
X_15995_ _17508_/X _15901_/A _17474_/X _15908_/A vssd1 vssd1 vccd1 vccd1 _15995_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_83_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17734_ _15375_/X _19711_/Q _18508_/D vssd1 vssd1 vccd1 vccd1 _17734_/X sky130_fd_sc_hd__mux2_1
X_10069_ _19925_/Q _10068_/Y _10057_/X _10042_/B vssd1 vssd1 vccd1 vccd1 _19925_/D
+ sky130_fd_sc_hd__o211a_1
X_14946_ _18085_/Q _14939_/X _14931_/X _14941_/X vssd1 vssd1 vccd1 vccd1 _18085_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_48_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17665_ _15574_/X _19470_/Q _17683_/S vssd1 vssd1 vccd1 vccd1 _18587_/D sky130_fd_sc_hd__mux2_1
X_14877_ _18126_/Q _14871_/X _14707_/X _14873_/X vssd1 vssd1 vccd1 vccd1 _18126_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18719__RESET_B repeater253/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17640__S _17655_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16616_ _16616_/A vssd1 vssd1 vccd1 vccd1 _16621_/B sky130_fd_sc_hd__buf_4
X_19404_ _19984_/CLK _19404_/D repeater243/X vssd1 vssd1 vccd1 vccd1 _19404_/Q sky130_fd_sc_hd__dfrtp_2
X_13828_ _13914_/A _13921_/A vssd1 vssd1 vccd1 vccd1 _13829_/B sky130_fd_sc_hd__or2_2
XFILLER_211_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17596_ _15344_/X _19707_/Q _17600_/S vssd1 vssd1 vccd1 vccd1 _17596_/X sky130_fd_sc_hd__mux2_1
XFILLER_223_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16547_ _16547_/A _16583_/B vssd1 vssd1 vccd1 vccd1 _16547_/Y sky130_fd_sc_hd__nor2_1
X_19335_ _20013_/CLK _19335_/D repeater242/X vssd1 vssd1 vccd1 vccd1 _19335_/Q sky130_fd_sc_hd__dfrtp_4
X_13759_ _18748_/Q _13758_/X _18748_/Q _13758_/X vssd1 vssd1 vccd1 vccd1 _18748_/D
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16483__C _17564_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19266_ _20035_/CLK _19266_/D repeater212/X vssd1 vssd1 vccd1 vccd1 _19266_/Q sky130_fd_sc_hd__dfrtp_2
X_16478_ _16905_/X _16597_/A _16903_/X _16598_/A vssd1 vssd1 vccd1 vccd1 _16481_/B
+ sky130_fd_sc_hd__a22oi_4
XANTENNA__17561__A1 _08945_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18217_ _19630_/CLK _18217_/D vssd1 vssd1 vccd1 vccd1 _18217_/Q sky130_fd_sc_hd__dfxtp_1
X_15429_ _19620_/Q _11165_/B _11166_/B vssd1 vssd1 vccd1 vccd1 _15429_/X sky130_fd_sc_hd__a21bo_1
XFILLER_164_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19197_ _19221_/CLK _19197_/D hold365/X vssd1 vssd1 vccd1 vccd1 _19197_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_117_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18148_ _19849_/CLK _18148_/D vssd1 vssd1 vccd1 vccd1 _18148_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_116_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold203 HADDR[1] vssd1 vssd1 vccd1 vccd1 input12/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17087__S _17546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold214 hold214/A vssd1 vssd1 vccd1 vccd1 hold214/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold225 hold225/A vssd1 vssd1 vccd1 vccd1 hold225/X sky130_fd_sc_hd__dlygate4sd3_1
X_18079_ _20124_/CLK _18079_/D vssd1 vssd1 vccd1 vccd1 _18079_/Q sky130_fd_sc_hd__dfxtp_1
Xhold236 hold236/A vssd1 vssd1 vccd1 vccd1 hold236/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 hold247/A vssd1 vssd1 vccd1 vccd1 hold247/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12436__D_N _19500_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12138__B1 _12069_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20110_ _20122_/CLK _20110_/D repeater217/X vssd1 vssd1 vccd1 vccd1 _20110_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_172_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold258 HWDATA[13] vssd1 vssd1 vccd1 vccd1 input42/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_236_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold269 HWDATA[9] vssd1 vssd1 vccd1 vccd1 input69/A sky130_fd_sc_hd__dlygate4sd3_1
X_09921_ _19357_/Q vssd1 vssd1 vccd1 vccd1 _09921_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12689__A1 _18973_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17077__A0 _17486_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20041_ _20051_/CLK _20041_/D repeater209/X vssd1 vssd1 vccd1 vccd1 _20041_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__19160__RESET_B hold370/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09852_ _09852_/A _09852_/B vssd1 vssd1 vccd1 vccd1 _09995_/A sky130_fd_sc_hd__or2_1
XFILLER_112_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10164__A2 _10155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09783_ _09742_/A _09742_/B _09734_/A _09781_/Y vssd1 vssd1 vccd1 vccd1 _19986_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_86_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_241_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18477__CLK _19780_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09217_ _19886_/Q vssd1 vssd1 vccd1 vccd1 _09217_/Y sky130_fd_sc_hd__inv_2
XFILLER_148_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09148_ _09151_/A vssd1 vssd1 vccd1 vccd1 _09156_/B sky130_fd_sc_hd__buf_1
XFILLER_136_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09079_ hold260/X vssd1 vssd1 vccd1 vccd1 _09079_/X sky130_fd_sc_hd__buf_6
XFILLER_163_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12129__B1 _11926_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11110_ _19637_/Q vssd1 vssd1 vccd1 vccd1 _11110_/Y sky130_fd_sc_hd__inv_2
XFILLER_135_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12090_ hold296/X vssd1 vssd1 vccd1 vccd1 _12090_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_146_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11041_ _19648_/Q _11040_/A _10267_/Y _11043_/A vssd1 vssd1 vccd1 vccd1 _19648_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_104_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16815__A0 _16814_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15753__B _15753_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13629__B1 _17614_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14800_ _15058_/A _15034_/B _15094_/C vssd1 vssd1 vccd1 vccd1 _14803_/A sky130_fd_sc_hd__or3_4
XFILLER_162_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15780_ _19905_/Q _19400_/Q vssd1 vssd1 vccd1 vccd1 _15780_/X sky130_fd_sc_hd__and2_2
X_12992_ _18936_/Q _12991_/Y _12879_/B _12980_/X vssd1 vssd1 vccd1 vccd1 _18936_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__11104__A1 _11093_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12301__B1 _12299_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14731_ _14743_/A _14731_/B _14784_/C vssd1 vssd1 vccd1 vccd1 _14733_/A sky130_fd_sc_hd__or3_4
X_11943_ _19397_/Q _11939_/X _09016_/X _11942_/X vssd1 vssd1 vccd1 vccd1 _19397_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_245_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17460__S _17548_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17450_ _17449_/X _13374_/Y _17535_/S vssd1 vssd1 vccd1 vccd1 _17450_/X sky130_fd_sc_hd__mux2_1
XFILLER_55_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14662_ _18246_/Q _14656_/X _14578_/X _14658_/X vssd1 vssd1 vccd1 vccd1 _18246_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_33_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11874_ _11914_/A vssd1 vssd1 vccd1 vccd1 _11891_/A sky130_fd_sc_hd__buf_2
XFILLER_45_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16401_ _18121_/Q vssd1 vssd1 vccd1 vccd1 _16401_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13613_ _18801_/Q vssd1 vssd1 vccd1 vccd1 _13613_/Y sky130_fd_sc_hd__inv_2
X_10825_ _10448_/A _17750_/X _17750_/S _10823_/Y _19723_/Q vssd1 vssd1 vccd1 vccd1
+ _19723_/D sky130_fd_sc_hd__a32o_1
X_17381_ _16215_/Y _19405_/Q _17517_/S vssd1 vssd1 vccd1 vccd1 _17381_/X sky130_fd_sc_hd__mux2_1
X_14593_ _18286_/Q _14587_/X _14578_/X _14589_/X vssd1 vssd1 vccd1 vccd1 _18286_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_232_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19120_ _19609_/CLK _19120_/D hold357/X vssd1 vssd1 vccd1 vccd1 _19120_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_198_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16332_ _17992_/Q vssd1 vssd1 vccd1 vccd1 _16332_/Y sky130_fd_sc_hd__inv_2
X_13544_ _13544_/A _13583_/A vssd1 vssd1 vccd1 vccd1 _13545_/B sky130_fd_sc_hd__or2_2
XFILLER_13_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10756_ _15283_/A vssd1 vssd1 vccd1 vccd1 _15389_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_201_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19051_ _19576_/CLK _19051_/D repeater255/X vssd1 vssd1 vccd1 vccd1 _19051_/Q sky130_fd_sc_hd__dfrtp_1
X_16263_ _18351_/Q vssd1 vssd1 vccd1 vccd1 _16263_/Y sky130_fd_sc_hd__inv_2
X_13475_ _13468_/A _13468_/B _13473_/Y _13437_/X vssd1 vssd1 vccd1 vccd1 _18845_/D
+ sky130_fd_sc_hd__a211oi_2
XANTENNA_repeater152_A _17385_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10687_ _15839_/A vssd1 vssd1 vccd1 vccd1 _15854_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__16804__S _17543_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10418__A _12232_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18002_ _18412_/CLK _18002_/D vssd1 vssd1 vccd1 vccd1 _18002_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12368__B1 _12238_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15214_ _15211_/A _15204_/X _15213_/X vssd1 vssd1 vccd1 vccd1 _18639_/D sky130_fd_sc_hd__o21ai_1
XFILLER_139_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12426_ _19133_/Q _12420_/X _12296_/X _12421_/X vssd1 vssd1 vccd1 vccd1 _19133_/D
+ sky130_fd_sc_hd__a22o_1
X_16194_ _18110_/Q vssd1 vssd1 vccd1 vccd1 _16194_/Y sky130_fd_sc_hd__inv_2
XFILLER_154_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15145_ _15145_/A _15145_/B _15145_/C vssd1 vssd1 vccd1 vccd1 _15147_/A sky130_fd_sc_hd__or3_4
X_12357_ _19168_/Q _12352_/X _12356_/X _12354_/X vssd1 vssd1 vccd1 vccd1 _19168_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_181_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output81_A _16524_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11308_ _18969_/Q vssd1 vssd1 vccd1 vccd1 _11308_/Y sky130_fd_sc_hd__inv_2
X_15076_ _18007_/Q _15071_/X hold244/X _15073_/X vssd1 vssd1 vccd1 vccd1 _18007_/D
+ sky130_fd_sc_hd__a22o_1
X_19953_ _19956_/CLK _19953_/D repeater245/X vssd1 vssd1 vccd1 vccd1 _19953_/Q sky130_fd_sc_hd__dfrtp_4
X_12288_ _19206_/Q _12283_/X _12030_/X _12284_/X vssd1 vssd1 vccd1 vccd1 _19206_/D
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_10_HCLK clkbuf_4_2_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20076_/CLK sky130_fd_sc_hd__clkbuf_16
X_14027_ _14027_/A _14108_/A vssd1 vssd1 vccd1 vccd1 _14028_/B sky130_fd_sc_hd__or2_2
XFILLER_113_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18904_ _19352_/CLK _18904_/D repeater212/X vssd1 vssd1 vccd1 vccd1 _18904_/Q sky130_fd_sc_hd__dfrtp_1
X_11239_ _19608_/Q vssd1 vssd1 vccd1 vccd1 _11488_/A sky130_fd_sc_hd__inv_2
X_19884_ _20050_/CLK _19884_/D repeater200/X vssd1 vssd1 vccd1 vccd1 _19884_/Q sky130_fd_sc_hd__dfrtp_1
X_18835_ _19255_/CLK _18835_/D repeater239/X vssd1 vssd1 vccd1 vccd1 _18835_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_209_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15978_ _15970_/Y _15971_/X _15972_/Y _15973_/X _15977_/X vssd1 vssd1 vccd1 vccd1
+ _15978_/X sky130_fd_sc_hd__o221a_1
XFILLER_36_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18766_ _19855_/CLK _18766_/D repeater264/X vssd1 vssd1 vccd1 vccd1 _18766_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__14293__B1 _14279_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_152_HCLK clkbuf_4_1_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19647_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_48_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17717_ _15423_/X _19524_/Q _18546_/D vssd1 vssd1 vccd1 vccd1 _17717_/X sky130_fd_sc_hd__mux2_1
X_14929_ _20078_/Q vssd1 vssd1 vccd1 vccd1 _14929_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_64_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18697_ _18701_/CLK _18697_/D hold351/X vssd1 vssd1 vccd1 vccd1 _18697_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__17231__A0 _15768_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17370__S _19498_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17648_ _15644_/X _19041_/Q _17655_/S vssd1 vssd1 vccd1 vccd1 _18604_/D sky130_fd_sc_hd__mux2_1
XANTENNA__19745__CLK _20070_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_223_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17579_ _15401_/X _19528_/Q _17584_/S vssd1 vssd1 vccd1 vccd1 _17579_/X sky130_fd_sc_hd__mux2_1
X_19318_ _19325_/CLK _19318_/D repeater213/X vssd1 vssd1 vccd1 vccd1 _19318_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_188_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19249_ _19324_/CLK _19249_/D repeater237/X vssd1 vssd1 vccd1 vccd1 _19249_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12359__B1 _12225_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09002_ _15749_/A _15821_/B vssd1 vssd1 vccd1 vccd1 _10686_/C sky130_fd_sc_hd__or2_1
XFILLER_118_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19341__RESET_B repeater245/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12543__A _14405_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17545__S _17545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09904_ _19331_/Q vssd1 vssd1 vccd1 vccd1 _09904_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12531__B1 _12302_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20024_ _20091_/CLK _20024_/D repeater236/X vssd1 vssd1 vccd1 vccd1 _20024_/Q sky130_fd_sc_hd__dfrtp_1
X_09835_ _19951_/Q vssd1 vssd1 vccd1 vccd1 _09859_/A sky130_fd_sc_hd__inv_2
XFILLER_100_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09766_ _09753_/A _09765_/A _19997_/Q _09765_/Y _09759_/X vssd1 vssd1 vccd1 vccd1
+ _19997_/D sky130_fd_sc_hd__o221a_1
XFILLER_101_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14284__B1 _13680_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_227_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_227_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09697_ _19420_/Q vssd1 vssd1 vccd1 vccd1 _09697_/Y sky130_fd_sc_hd__inv_2
XPHY_4026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrebuffer40 _17055_/A1 vssd1 vssd1 vccd1 vccd1 _12147_/A1 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_4037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17280__S _17534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrebuffer51 _09859_/B vssd1 vssd1 vccd1 vccd1 _09985_/C1 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_4048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer62 _13539_/B vssd1 vssd1 vccd1 vccd1 _13595_/C1 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrebuffer73 _11461_/B vssd1 vssd1 vccd1 vccd1 _11540_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14036__B1 _19078_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_215_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrebuffer84 _11463_/B vssd1 vssd1 vccd1 vccd1 _11539_/C1 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_82_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrebuffer95 _13537_/C vssd1 vssd1 vccd1 vccd1 _13599_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10610_ _19812_/Q _10606_/X _10615_/A _10609_/X vssd1 vssd1 vccd1 vccd1 _19812_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11590_ _11590_/A _11590_/B vssd1 vssd1 vccd1 vccd1 _11591_/C sky130_fd_sc_hd__nor2_1
XPHY_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12437__B _15863_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10541_ _19813_/Q vssd1 vssd1 vccd1 vccd1 _10595_/A sky130_fd_sc_hd__clkbuf_2
XPHY_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13260_ _18756_/Q vssd1 vssd1 vccd1 vccd1 _13723_/A sky130_fd_sc_hd__inv_2
XFILLER_210_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10472_ _10472_/A vssd1 vssd1 vccd1 vccd1 _10472_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_33_HCLK _18641_/CLK vssd1 vssd1 vccd1 vccd1 _18137_/CLK sky130_fd_sc_hd__clkbuf_16
X_12211_ _19244_/Q _12205_/X _12104_/X _12206_/X vssd1 vssd1 vccd1 vccd1 _19244_/D
+ sky130_fd_sc_hd__a22o_1
X_13191_ _18902_/Q _13190_/Y _13180_/X _13191_/C1 vssd1 vssd1 vccd1 vccd1 _18902_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_151_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_191_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12142_ _19289_/Q _12134_/X _12080_/X _12137_/X vssd1 vssd1 vccd1 vccd1 _19289_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_135_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17455__S _17546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12073_ _19325_/Q _12068_/X _12069_/X _12072_/X vssd1 vssd1 vccd1 vccd1 _19325_/D
+ sky130_fd_sc_hd__a22o_1
X_16950_ _19494_/Q hold139/X _16950_/S vssd1 vssd1 vccd1 vccd1 _16950_/X sky130_fd_sc_hd__mux2_1
XFILLER_151_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12522__B1 _12356_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11024_ _11023_/Y _17753_/S _19650_/Q _11029_/A vssd1 vssd1 vccd1 vccd1 _11025_/B
+ sky130_fd_sc_hd__o22a_1
X_15901_ _15901_/A vssd1 vssd1 vccd1 vccd1 _16506_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_103_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16881_ _16880_/X _09496_/Y _17414_/S vssd1 vssd1 vccd1 vccd1 _16881_/X sky130_fd_sc_hd__mux2_1
XFILLER_38_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15832_ _15832_/A _15850_/B vssd1 vssd1 vccd1 vccd1 _15832_/X sky130_fd_sc_hd__or2_1
X_18620_ _18623_/CLK hold230/X hold351/X vssd1 vssd1 vccd1 vccd1 _18620_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_49_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18642__CLK _18642_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15763_ _18521_/Q _18522_/Q _18523_/Q vssd1 vssd1 vccd1 vccd1 _18521_/D sky130_fd_sc_hd__o21ba_1
X_18551_ _19780_/CLK _18551_/D repeater227/X vssd1 vssd1 vccd1 vccd1 _18551_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_46_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12825__A1 _19235_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12975_ _12975_/A vssd1 vssd1 vccd1 vccd1 _12975_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17190__S _17545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17502_ _17501_/X _13254_/Y _17567_/S vssd1 vssd1 vccd1 vccd1 _17502_/X sky130_fd_sc_hd__mux2_1
X_14714_ _18219_/Q _14700_/A _14713_/X _14701_/A vssd1 vssd1 vccd1 vccd1 _18219_/D
+ sky130_fd_sc_hd__a22o_1
X_18482_ _19545_/CLK _18482_/D repeater225/X vssd1 vssd1 vccd1 vccd1 _18482_/Q sky130_fd_sc_hd__dfrtp_1
X_11926_ _11926_/A vssd1 vssd1 vccd1 vccd1 _11926_/X sky130_fd_sc_hd__buf_4
XFILLER_206_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15694_ _18616_/Q _15693_/A _15692_/Y _15693_/Y vssd1 vssd1 vccd1 vccd1 _15695_/B
+ sky130_fd_sc_hd__o22a_1
XPHY_4560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17433_ _17432_/X _17879_/X _17568_/S vssd1 vssd1 vccd1 vccd1 _17433_/X sky130_fd_sc_hd__mux2_2
XPHY_4582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14645_ _14645_/A vssd1 vssd1 vccd1 vccd1 _14645_/X sky130_fd_sc_hd__clkbuf_2
XPHY_4593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11857_ _19330_/Q vssd1 vssd1 vccd1 vccd1 _13641_/A sky130_fd_sc_hd__buf_1
XFILLER_220_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12589__B1 hold270/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10808_ _10809_/A vssd1 vssd1 vccd1 vccd1 _10808_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_14_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17364_ _17363_/X _14068_/Y _17544_/S vssd1 vssd1 vccd1 vccd1 _17364_/X sky130_fd_sc_hd__mux2_1
XPHY_3892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14576_ _18296_/Q _14572_/X _14535_/X _14574_/X vssd1 vssd1 vccd1 vccd1 _18296_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_220_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11788_ _19470_/Q _11784_/X _09016_/X _11787_/X vssd1 vssd1 vccd1 vccd1 _19470_/D
+ sky130_fd_sc_hd__a22o_1
X_16315_ _18877_/Q vssd1 vssd1 vccd1 vccd1 _16315_/Y sky130_fd_sc_hd__inv_2
X_19103_ _19109_/CLK _19103_/D hold361/X vssd1 vssd1 vccd1 vccd1 _19103_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_186_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13527_ _13491_/Y _17759_/X _13499_/X _13526_/X vssd1 vssd1 vccd1 vccd1 _18836_/D
+ sky130_fd_sc_hd__o22ai_1
X_10739_ _19764_/Q _10738_/X _17757_/X vssd1 vssd1 vccd1 vccd1 _19764_/D sky130_fd_sc_hd__mux2_1
XFILLER_201_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17295_ _17294_/X _16500_/Y _17541_/S vssd1 vssd1 vccd1 vccd1 _17295_/X sky130_fd_sc_hd__mux2_1
XFILLER_185_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19034_ _19577_/CLK _19034_/D repeater267/X vssd1 vssd1 vccd1 vccd1 _19034_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_185_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16246_ _17388_/X _16597_/A _17392_/X _16594_/A vssd1 vssd1 vccd1 vccd1 _16246_/Y
+ sky130_fd_sc_hd__a22oi_4
XFILLER_118_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13458_ _13430_/B _13338_/B _13456_/Y _13445_/X vssd1 vssd1 vccd1 vccd1 _18851_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_173_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12409_ _19144_/Q _12400_/X _12408_/X _12402_/X vssd1 vssd1 vccd1 vccd1 _19144_/D
+ sky130_fd_sc_hd__a22o_1
X_16177_ _18126_/Q vssd1 vssd1 vccd1 vccd1 _16177_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13389_ _20101_/Q _13470_/A _20113_/Q _13431_/D _13388_/X vssd1 vssd1 vccd1 vccd1
+ _13389_/X sky130_fd_sc_hd__a221o_1
Xoutput105 _16251_/Y vssd1 vssd1 vccd1 vccd1 HRDATA[4] sky130_fd_sc_hd__clkbuf_2
XFILLER_115_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput116 _16756_/LO vssd1 vssd1 vccd1 vccd1 IRQ[13] sky130_fd_sc_hd__clkbuf_2
XFILLER_142_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput127 _15779_/X vssd1 vssd1 vccd1 vccd1 IRQ[9] sky130_fd_sc_hd__clkbuf_2
XFILLER_127_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput138 _16759_/LO vssd1 vssd1 vccd1 vccd1 scl_o_S4 sky130_fd_sc_hd__clkbuf_2
X_15128_ _17973_/Q _15122_/X _14929_/X _15124_/X vssd1 vssd1 vccd1 vccd1 _17973_/D
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_3_3_0_HCLK clkbuf_3_3_0_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_7_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__18172__CLK _18198_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19298__CLK _20013_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17365__S _17545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19936_ _19937_/CLK _19936_/D repeater236/X vssd1 vssd1 vccd1 vccd1 _19936_/Q sky130_fd_sc_hd__dfrtp_1
X_15059_ _15060_/A vssd1 vssd1 vccd1 vccd1 _15059_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_99_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19867_ _19867_/CLK _19867_/D repeater263/X vssd1 vssd1 vccd1 vccd1 _19867_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_110_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17452__A0 _17486_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09620_ _09620_/A vssd1 vssd1 vccd1 vccd1 _10029_/B sky130_fd_sc_hd__clkinv_1
X_18818_ _18856_/CLK _18818_/D repeater231/X vssd1 vssd1 vccd1 vccd1 _18818_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_244_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19798_ _19808_/CLK _19798_/D repeater222/X vssd1 vssd1 vccd1 vccd1 _19798_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_209_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09551_ _19295_/Q vssd1 vssd1 vccd1 vccd1 _09551_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18749_ _19900_/CLK _18749_/D repeater199/X vssd1 vssd1 vccd1 vccd1 _18749_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_237_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09482_ _09482_/A _09482_/B vssd1 vssd1 vccd1 vccd1 _09589_/A sky130_fd_sc_hd__or2_1
XANTENNA__17755__A1 _11059_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_212_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17850__S1 _19632_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12538__A _13678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17507__A1 _12058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_56_HCLK clkbuf_4_9_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20049_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_149_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15849__A _19756_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_180_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_180_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20080__RESET_B repeater204/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17275__S _17548_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12504__B1 _12398_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17443__A0 _17486_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20007_ _20013_/CLK _20007_/D repeater241/X vssd1 vssd1 vccd1 vccd1 _20007_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__11617__A _11617_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09818_ _19968_/Q vssd1 vssd1 vccd1 vccd1 _09876_/A sky130_fd_sc_hd__inv_2
XFILLER_246_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09749_ _09749_/A _09772_/A vssd1 vssd1 vccd1 vccd1 _09750_/B sky130_fd_sc_hd__or2_2
XFILLER_15_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12760_ _19229_/Q vssd1 vssd1 vccd1 vccd1 _12760_/Y sky130_fd_sc_hd__inv_2
XPHY_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17746__A1 _11153_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ _11731_/A vssd1 vssd1 vccd1 vccd1 _16950_/S sky130_fd_sc_hd__buf_6
XFILLER_242_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12691_ _12698_/A vssd1 vssd1 vccd1 vccd1 _12691_/X sky130_fd_sc_hd__clkbuf_2
XPHY_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17841__S1 _19632_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_202_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14430_ _18382_/Q _14424_/X _14415_/X _14426_/X vssd1 vssd1 vccd1 vccd1 _18382_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_14_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11642_ _11642_/A vssd1 vssd1 vccd1 vccd1 _11645_/A sky130_fd_sc_hd__inv_2
XPHY_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13232__B2 _17584_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14361_ _18422_/Q _14349_/X hold324/X _14353_/X vssd1 vssd1 vccd1 vccd1 _18422_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11573_ _11573_/A _11573_/B vssd1 vssd1 vccd1 vccd1 _11612_/A sky130_fd_sc_hd__or2_1
XPHY_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19263__RESET_B repeater212/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput18 HADDR[25] vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__buf_1
XPHY_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16100_ _17972_/Q vssd1 vssd1 vccd1 vccd1 _16100_/Y sky130_fd_sc_hd__inv_2
X_13312_ _18853_/Q vssd1 vssd1 vccd1 vccd1 _13429_/D sky130_fd_sc_hd__inv_2
XFILLER_10_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10524_ _19536_/Q vssd1 vssd1 vccd1 vccd1 _10525_/B sky130_fd_sc_hd__inv_2
XFILLER_167_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput29 input29/A vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__buf_1
X_17080_ _17486_/A0 _16438_/Y _17517_/S vssd1 vssd1 vccd1 vccd1 _17080_/X sky130_fd_sc_hd__mux2_1
X_14292_ _18456_/Q _14288_/X _14277_/X _14290_/X vssd1 vssd1 vccd1 vccd1 _18456_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16031_ _18252_/Q vssd1 vssd1 vccd1 vccd1 _16031_/Y sky130_fd_sc_hd__inv_2
X_13243_ _13243_/A vssd1 vssd1 vccd1 vccd1 _13243_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__13279__A _19518_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10455_ _19829_/Q _10450_/X _10421_/X _10452_/X vssd1 vssd1 vccd1 vccd1 _19829_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12183__A _12187_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13174_ _13083_/A _13174_/A2 _13172_/Y _13199_/B vssd1 vssd1 vccd1 vccd1 _18911_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_163_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10386_ _10345_/X _08921_/X _10368_/X _10385_/X vssd1 vssd1 vccd1 vccd1 _19853_/D
+ sky130_fd_sc_hd__o22ai_1
XANTENNA__10415__B _15826_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17185__S _17546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15494__A _15571_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12125_ _19298_/Q _12121_/X _11918_/X _12122_/X vssd1 vssd1 vccd1 vccd1 _19298_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_124_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17982_ _20124_/CLK _17982_/D vssd1 vssd1 vccd1 vccd1 _17982_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19721_ _19795_/CLK _19721_/D repeater226/X vssd1 vssd1 vccd1 vccd1 _19721_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_238_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12056_ _12056_/A vssd1 vssd1 vccd1 vccd1 _12056_/Y sky130_fd_sc_hd__inv_2
X_16933_ _19477_/Q hold190/X _16946_/S vssd1 vssd1 vccd1 vccd1 _16933_/X sky130_fd_sc_hd__mux2_1
XFILLER_120_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11007_ _11002_/B _11006_/Y _10973_/B _10989_/X _10958_/A vssd1 vssd1 vccd1 vccd1
+ _11008_/A sky130_fd_sc_hd__o32a_1
X_19652_ _19873_/CLK _19652_/D repeater265/X vssd1 vssd1 vccd1 vccd1 _19652_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_226_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16864_ _17473_/A0 _09884_/Y _17522_/S vssd1 vssd1 vccd1 vccd1 _16864_/X sky130_fd_sc_hd__mux2_1
XFILLER_203_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18603_ _19041_/CLK _18603_/D repeater263/X vssd1 vssd1 vccd1 vccd1 _18603_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_93_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15815_ _18082_/Q vssd1 vssd1 vccd1 vccd1 _15815_/Y sky130_fd_sc_hd__inv_2
X_19583_ _19591_/CLK _19583_/D hold363/X vssd1 vssd1 vccd1 vccd1 _19583_/Q sky130_fd_sc_hd__dfrtp_4
X_16795_ _16794_/X _19222_/Q _17545_/S vssd1 vssd1 vccd1 vccd1 _16795_/X sky130_fd_sc_hd__mux2_1
XFILLER_219_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10150__B _15883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_234_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15746_ _18664_/Q vssd1 vssd1 vccd1 vccd1 _15746_/Y sky130_fd_sc_hd__inv_2
X_18534_ _19822_/CLK _18534_/D repeater228/X vssd1 vssd1 vccd1 vccd1 _18534_/Q sky130_fd_sc_hd__dfrtp_1
X_12958_ _13060_/B vssd1 vssd1 vccd1 vccd1 _12958_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_93_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_79_HCLK clkbuf_4_13_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _18947_/CLK sky130_fd_sc_hd__clkbuf_16
X_11909_ hold268/X vssd1 vssd1 vccd1 vccd1 _11909_/X sky130_fd_sc_hd__clkbuf_4
X_15677_ _15681_/B vssd1 vssd1 vccd1 vccd1 _15683_/B sky130_fd_sc_hd__inv_2
X_18465_ _18465_/CLK _18465_/D vssd1 vssd1 vccd1 vccd1 _18465_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_178_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17832__S1 _18750_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12889_ _12889_/A vssd1 vssd1 vccd1 vccd1 _12890_/B sky130_fd_sc_hd__inv_2
XPHY_4390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17416_ _17415_/X _13397_/Y _17529_/S vssd1 vssd1 vccd1 vccd1 _17416_/X sky130_fd_sc_hd__mux2_1
X_14628_ _14628_/A _14628_/B _15195_/B vssd1 vssd1 vccd1 vccd1 _15157_/C sky130_fd_sc_hd__or3_4
X_18396_ _18416_/CLK _18396_/D vssd1 vssd1 vccd1 vccd1 _18396_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14420__B1 _14419_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17347_ _17473_/A0 _16300_/Y _17473_/S vssd1 vssd1 vccd1 vccd1 _17347_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14559_ _14559_/A vssd1 vssd1 vccd1 vccd1 _14560_/A sky130_fd_sc_hd__inv_2
XFILLER_159_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17278_ _17473_/A0 _16518_/Y _17547_/S vssd1 vssd1 vccd1 vccd1 _17278_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16229_ _19525_/Q vssd1 vssd1 vccd1 vccd1 _16229_/Y sky130_fd_sc_hd__inv_2
XFILLER_146_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19017_ _19115_/CLK _19017_/D hold353/X vssd1 vssd1 vccd1 vccd1 _19017_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_162_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17899__S1 _18761_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17095__S _17545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12821__A _19233_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08982_ _08982_/A _08982_/B vssd1 vssd1 vccd1 vccd1 _08983_/B sky130_fd_sc_hd__or2_1
XFILLER_130_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19919_ _19927_/CLK _19919_/D repeater230/X vssd1 vssd1 vccd1 vccd1 _19919_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_69_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_244_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09603_ _09474_/B _09605_/A _09474_/A vssd1 vssd1 vccd1 vccd1 _09604_/C sky130_fd_sc_hd__o21a_1
XFILLER_84_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18068__CLK _19851_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09534_ _19297_/Q vssd1 vssd1 vccd1 vccd1 _09534_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17728__A1 _19685_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_224_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09465_ _09465_/A _09465_/B vssd1 vssd1 vccd1 vccd1 _09618_/A sky130_fd_sc_hd__or2_2
XFILLER_52_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17823__S1 _18750_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_104_HCLK_A clkbuf_4_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_240_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09396_ _19373_/Q vssd1 vssd1 vccd1 vccd1 _09396_/Y sky130_fd_sc_hd__inv_2
XFILLER_178_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11776__A1 hold202/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16902__S _17385_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10240_ _19828_/Q vssd1 vssd1 vccd1 vccd1 _10240_/Y sky130_fd_sc_hd__inv_2
XFILLER_79_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18656__RESET_B repeater210/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10171_ _19885_/Q _10166_/X _09082_/X _10168_/X vssd1 vssd1 vccd1 vccd1 _19885_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_78_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17733__S _18508_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13930_ _18725_/Q _13929_/Y _13907_/X _13825_/B vssd1 vssd1 vccd1 vccd1 _18725_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_47_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_208_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13861_ _13844_/Y _18720_/Q _13860_/Y _18725_/Q vssd1 vssd1 vccd1 vccd1 _13861_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_170_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15600_ _18594_/Q vssd1 vssd1 vccd1 vccd1 _15602_/A sky130_fd_sc_hd__inv_2
XFILLER_75_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_216_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12812_ _18824_/Q vssd1 vssd1 vccd1 vccd1 _13547_/A sky130_fd_sc_hd__inv_2
XFILLER_170_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16580_ _17143_/X _16577_/X _17256_/X _16578_/X _16579_/X vssd1 vssd1 vccd1 vccd1
+ _16581_/C sky130_fd_sc_hd__o221a_1
XFILLER_27_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13792_ _18720_/Q vssd1 vssd1 vccd1 vccd1 _13910_/D sky130_fd_sc_hd__inv_2
XFILLER_103_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15531_ _15530_/A _15530_/B _15530_/Y vssd1 vssd1 vccd1 vccd1 _15532_/B sky130_fd_sc_hd__a21oi_1
X_12743_ _19241_/Q vssd1 vssd1 vccd1 vccd1 _16546_/A sky130_fd_sc_hd__inv_2
XANTENNA__17814__S1 _18752_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_230_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18250_ _18268_/CLK _18250_/D vssd1 vssd1 vccd1 vccd1 _18250_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15462_ _15462_/A vssd1 vssd1 vccd1 vccd1 _15467_/B sky130_fd_sc_hd__inv_2
XFILLER_188_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12674_ _18984_/Q _12670_/X hold306/X _12671_/X vssd1 vssd1 vccd1 vccd1 _18984_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_43_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14402__B1 _14329_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17201_ _17200_/X _13369_/Y _17535_/S vssd1 vssd1 vccd1 vccd1 _17201_/X sky130_fd_sc_hd__mux2_1
XPHY_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14413_ _18392_/Q _14409_/X _14356_/X _14411_/X vssd1 vssd1 vccd1 vccd1 _18392_/D
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_8_HCLK clkbuf_4_2_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _18473_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11625_ _11625_/A _11629_/A vssd1 vssd1 vccd1 vccd1 _11626_/B sky130_fd_sc_hd__or2_2
X_18181_ _18216_/CLK _18181_/D vssd1 vssd1 vccd1 vccd1 _18181_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15393_ _15419_/A vssd1 vssd1 vccd1 vccd1 _15402_/A sky130_fd_sc_hd__buf_1
XPHY_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_26_HCLK_A clkbuf_4_9_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17132_ _16551_/Y _15632_/Y _17318_/S vssd1 vssd1 vccd1 vccd1 _17132_/X sky130_fd_sc_hd__mux2_2
XPHY_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14344_ _18428_/Q _14337_/A _14329_/X _14338_/A vssd1 vssd1 vccd1 vccd1 _18428_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11556_ _11574_/A _11573_/A _11556_/C _11556_/D vssd1 vssd1 vccd1 vccd1 _11559_/B
+ sky130_fd_sc_hd__or4_4
XPHY_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_89_HCLK_A clkbuf_4_12_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10507_ _19545_/Q _19534_/Q vssd1 vssd1 vccd1 vccd1 _10508_/B sky130_fd_sc_hd__or2_1
XFILLER_144_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17063_ _17062_/X _11408_/Y _17548_/S vssd1 vssd1 vccd1 vccd1 _17063_/X sky130_fd_sc_hd__mux2_1
XANTENNA_repeater232_A repeater233/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14275_ _14275_/A vssd1 vssd1 vccd1 vccd1 _14275_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_171_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11487_ _11487_/A _11494_/A vssd1 vssd1 vccd1 vccd1 _11488_/B sky130_fd_sc_hd__or2_1
XANTENNA__16812__S _17545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16014_ _18052_/Q vssd1 vssd1 vccd1 vccd1 _16014_/Y sky130_fd_sc_hd__inv_2
X_13226_ _18539_/Q _13226_/B vssd1 vssd1 vccd1 vccd1 _13227_/B sky130_fd_sc_hd__or2_1
XFILLER_170_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10438_ _19839_/Q _10433_/X _09064_/X _10435_/X vssd1 vssd1 vccd1 vccd1 _19839_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_170_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13157_ _19189_/Q _13091_/Y _19182_/Q _13083_/A vssd1 vssd1 vccd1 vccd1 _13157_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_112_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10369_ _10364_/B _10367_/Y _10368_/X _10354_/X _10324_/A vssd1 vssd1 vccd1 vccd1
+ _10370_/A sky130_fd_sc_hd__o32a_1
XANTENNA__14469__B1 _14415_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12108_ _12122_/A vssd1 vssd1 vccd1 vccd1 _12108_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_111_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17965_ _19842_/CLK _17965_/D vssd1 vssd1 vccd1 vccd1 _17965_/Q sky130_fd_sc_hd__dfxtp_1
X_13088_ _13088_/A _13166_/A vssd1 vssd1 vccd1 vccd1 _13089_/B sky130_fd_sc_hd__or2_2
XFILLER_100_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17407__A0 _17486_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19704_ _20057_/CLK _19704_/D repeater202/X vssd1 vssd1 vccd1 vccd1 _19704_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__17643__S _17655_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16916_ _16915_/X _15533_/Y _17474_/S vssd1 vssd1 vccd1 vccd1 _16916_/X sky130_fd_sc_hd__mux2_1
X_12039_ _19341_/Q _12034_/X _12038_/X _12036_/X vssd1 vssd1 vccd1 vccd1 _19341_/D
+ sky130_fd_sc_hd__a22o_1
X_17896_ _15944_/Y _15945_/Y _15946_/Y _15947_/Y _17908_/S0 _18759_/Q vssd1 vssd1
+ vccd1 vccd1 _17896_/X sky130_fd_sc_hd__mux4_2
XANTENNA__19336__CLK _20013_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19635_ _19637_/CLK _19635_/D repeater258/X vssd1 vssd1 vccd1 vccd1 _19635_/Q sky130_fd_sc_hd__dfrtp_4
X_16847_ _16846_/X _13087_/A _17488_/S vssd1 vssd1 vccd1 vccd1 _16847_/X sky130_fd_sc_hd__mux2_1
XFILLER_226_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19566_ _19566_/CLK _19566_/D repeater255/X vssd1 vssd1 vccd1 vccd1 _19566_/Q sky130_fd_sc_hd__dfrtp_1
X_16778_ _16723_/Y _15696_/Y _17474_/S vssd1 vssd1 vccd1 vccd1 _16778_/X sky130_fd_sc_hd__mux2_1
XFILLER_46_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18517_ _19822_/CLK _18517_/D repeater227/X vssd1 vssd1 vccd1 vccd1 _18517_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_80_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_234_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15729_ _20041_/Q vssd1 vssd1 vccd1 vccd1 _15729_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19486__CLK _19510_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12088__A hold306/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17805__S1 _18750_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19497_ _20036_/CLK _19497_/D repeater198/X vssd1 vssd1 vccd1 vccd1 _19497_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_178_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09250_ _20061_/Q _20062_/Q _09250_/S vssd1 vssd1 vccd1 vccd1 _20062_/D sky130_fd_sc_hd__mux2_1
XFILLER_222_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18448_ _19668_/CLK _18448_/D vssd1 vssd1 vccd1 vccd1 _18448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_221_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09181_ _14711_/A _09164_/A _09180_/X _09165_/A vssd1 vssd1 vccd1 vccd1 _20076_/D
+ sky130_fd_sc_hd__a22o_1
X_18379_ _19515_/CLK _18379_/D vssd1 vssd1 vccd1 vccd1 _18379_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16146__B1 _17433_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08965_ _19858_/Q vssd1 vssd1 vccd1 vccd1 _10324_/A sky130_fd_sc_hd__inv_2
XFILLER_248_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15862__A _19024_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12486__A2 _12457_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19955__RESET_B repeater245/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_229_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11694__B1 _10882_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09517_ _19324_/Q vssd1 vssd1 vccd1 vccd1 _09517_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09448_ _19923_/Q vssd1 vssd1 vccd1 vccd1 _10039_/A sky130_fd_sc_hd__inv_2
XFILLER_13_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18853__CLK _18866_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19979__CLK _19992_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_200_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09379_ _19932_/Q _09374_/Y _19926_/Q _09375_/Y _09378_/X vssd1 vssd1 vccd1 vccd1
+ _09379_/X sky130_fd_sc_hd__a221o_1
XFILLER_12_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11410_ _19577_/Q _11408_/Y _19569_/Q _11409_/Y vssd1 vssd1 vccd1 vccd1 _11410_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_184_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12390_ _12402_/A vssd1 vssd1 vccd1 vccd1 _12390_/X sky130_fd_sc_hd__buf_1
XFILLER_123_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18837__RESET_B repeater231/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09100__A hold264/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11341_ _18986_/Q vssd1 vssd1 vccd1 vccd1 _11341_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14060_ _19091_/Q vssd1 vssd1 vccd1 vccd1 _14060_/Y sky130_fd_sc_hd__inv_2
X_11272_ _11479_/A _19013_/Q _19595_/Q _16582_/A vssd1 vssd1 vccd1 vccd1 _11272_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_3_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13371__B1 _20101_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13011_ _13011_/A vssd1 vssd1 vccd1 vccd1 _13011_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10223_ _19654_/Q vssd1 vssd1 vccd1 vccd1 _10956_/A sky130_fd_sc_hd__inv_2
XFILLER_106_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10185__B1 _19876_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10154_ _10155_/A vssd1 vssd1 vccd1 vccd1 _10154_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_121_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15772__A _15772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17463__S _17564_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17750_ _15735_/B _19700_/Q _17750_/S vssd1 vssd1 vccd1 vccd1 _17750_/X sky130_fd_sc_hd__mux2_2
X_14962_ _18074_/Q _14953_/A _14949_/X _14954_/A vssd1 vssd1 vccd1 vccd1 _18074_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_248_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10085_ _10085_/A _10094_/A vssd1 vssd1 vccd1 vccd1 _10086_/B sky130_fd_sc_hd__or2_1
XFILLER_87_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_248_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16587__B _16615_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16701_ _16809_/X _16633_/X _16824_/X _16634_/X vssd1 vssd1 vccd1 vccd1 _16701_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_235_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13913_ _19125_/Q _13927_/A vssd1 vssd1 vccd1 vccd1 _13913_/X sky130_fd_sc_hd__or2_1
XFILLER_208_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14893_ _18114_/Q _14884_/A _14842_/X _14885_/A vssd1 vssd1 vccd1 vccd1 _18114_/D
+ sky130_fd_sc_hd__a22o_1
X_17681_ _15507_/X _19454_/Q _17683_/S vssd1 vssd1 vccd1 vccd1 _18571_/D sky130_fd_sc_hd__mux2_1
XFILLER_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16612__A1 _16866_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19420_ _19997_/CLK _19420_/D repeater192/X vssd1 vssd1 vccd1 vccd1 _19420_/Q sky130_fd_sc_hd__dfrtp_1
X_16632_ _19046_/Q vssd1 vssd1 vccd1 vccd1 _16632_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16612__B2 _15887_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13844_ _19209_/Q vssd1 vssd1 vccd1 vccd1 _13844_/Y sky130_fd_sc_hd__inv_2
XFILLER_223_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19351_ _19352_/CLK _19351_/D repeater245/X vssd1 vssd1 vccd1 vccd1 _19351_/Q sky130_fd_sc_hd__dfrtp_1
X_16563_ _16638_/A vssd1 vssd1 vccd1 vccd1 _16563_/X sky130_fd_sc_hd__clkbuf_4
X_13775_ _18662_/Q _18737_/Q _13775_/S vssd1 vssd1 vccd1 vccd1 _18737_/D sky130_fd_sc_hd__mux2_1
XANTENNA__16807__S _17534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10987_ _10987_/A vssd1 vssd1 vccd1 vccd1 _10988_/B sky130_fd_sc_hd__inv_2
XFILLER_90_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_188_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17799__S0 _19647_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_231_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18302_ _18431_/CLK _18302_/D vssd1 vssd1 vccd1 vccd1 _18302_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_200_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15514_ _18573_/Q vssd1 vssd1 vccd1 vccd1 _15514_/Y sky130_fd_sc_hd__inv_2
X_12726_ _14812_/A vssd1 vssd1 vccd1 vccd1 _12726_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_204_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16494_ _16494_/A vssd1 vssd1 vccd1 vccd1 _16687_/A sky130_fd_sc_hd__buf_2
X_19282_ _19282_/CLK _19282_/D repeater216/X vssd1 vssd1 vccd1 vccd1 _19282_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_31_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18233_ _18412_/CLK _18233_/D vssd1 vssd1 vccd1 vccd1 _18233_/Q sky130_fd_sc_hd__dfxtp_1
X_15445_ _15571_/A vssd1 vssd1 vccd1 vccd1 _15479_/A sky130_fd_sc_hd__buf_4
X_12657_ _18993_/Q _12629_/A _12541_/X _12630_/A vssd1 vssd1 vccd1 vccd1 _18993_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12636__A _12650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_150_HCLK_A clkbuf_4_1_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20112__RESET_B repeater217/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11608_ _11577_/A _11577_/B _11569_/A _11606_/Y vssd1 vssd1 vccd1 vccd1 _19564_/D
+ sky130_fd_sc_hd__a211oi_2
X_15376_ _19792_/Q _10652_/B _10653_/B vssd1 vssd1 vccd1 vccd1 _15376_/X sky130_fd_sc_hd__a21bo_1
XFILLER_168_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18164_ _18165_/CLK _18164_/D vssd1 vssd1 vccd1 vccd1 _18164_/Q sky130_fd_sc_hd__dfxtp_1
X_12588_ _19038_/Q _12583_/X hold256/X _12584_/X vssd1 vssd1 vccd1 vccd1 _19038_/D
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_109_HCLK clkbuf_4_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19585_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__18578__RESET_B repeater269/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17638__S _17655_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14327_ _18437_/Q _14318_/X _14326_/X _14320_/X vssd1 vssd1 vccd1 vccd1 _18437_/D
+ sky130_fd_sc_hd__a22o_1
X_17115_ _17473_/A0 _16560_/Y _17512_/S vssd1 vssd1 vccd1 vccd1 _17115_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18095_ _20090_/CLK _18095_/D vssd1 vssd1 vccd1 vccd1 _18095_/Q sky130_fd_sc_hd__dfxtp_1
X_11539_ _19581_/Q _11538_/Y _11521_/X _11539_/C1 vssd1 vssd1 vccd1 vccd1 _19581_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__18507__RESET_B repeater222/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17046_ _15768_/Y _14187_/Y _17546_/S vssd1 vssd1 vccd1 vccd1 _17046_/X sky130_fd_sc_hd__mux2_1
XANTENNA__14154__A2 _18701_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14258_ _14259_/A vssd1 vssd1 vccd1 vccd1 _14258_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_99_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13209_ _13064_/A _13209_/A2 _13207_/Y _13202_/X vssd1 vssd1 vccd1 vccd1 _18891_/D
+ sky130_fd_sc_hd__a211oi_2
X_14189_ _19116_/Q vssd1 vssd1 vccd1 vccd1 _14189_/Y sky130_fd_sc_hd__inv_2
XANTENNA__10176__B1 _09094_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11912__A1 _19409_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18997_ _19137_/CLK _18997_/D repeater249/X vssd1 vssd1 vccd1 vccd1 _18997_/Q sky130_fd_sc_hd__dfrtp_4
Xrepeater202 repeater203/X vssd1 vssd1 vccd1 vccd1 repeater202/X sky130_fd_sc_hd__buf_8
XANTENNA__17373__S _17568_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater213 repeater214/X vssd1 vssd1 vccd1 vccd1 repeater213/X sky130_fd_sc_hd__buf_8
XFILLER_100_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17948_ _18765_/CLK _17948_/D vssd1 vssd1 vccd1 vccd1 _17948_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_227_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater224 repeater225/X vssd1 vssd1 vccd1 vccd1 repeater224/X sky130_fd_sc_hd__buf_4
Xrepeater235 repeater236/X vssd1 vssd1 vccd1 vccd1 repeater235/X sky130_fd_sc_hd__buf_6
XFILLER_39_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrepeater246 hold372/A vssd1 vssd1 vccd1 vccd1 hold373/A sky130_fd_sc_hd__buf_4
Xrepeater257 repeater258/X vssd1 vssd1 vccd1 vccd1 repeater257/X sky130_fd_sc_hd__buf_8
Xrepeater268 repeater269/X vssd1 vssd1 vccd1 vccd1 repeater268/X sky130_fd_sc_hd__buf_6
X_17879_ _17875_/X _17876_/X _17877_/X _17878_/X _18760_/Q _18761_/Q vssd1 vssd1 vccd1
+ vccd1 _17879_/X sky130_fd_sc_hd__mux4_2
XFILLER_238_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater279 hold360/A vssd1 vssd1 vccd1 vccd1 hold362/A sky130_fd_sc_hd__buf_8
XFILLER_26_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19618_ _19937_/CLK _19618_/D repeater230/X vssd1 vssd1 vccd1 vccd1 _19618_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__16603__B2 _15898_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19549_ _19561_/CLK _19549_/D repeater269/X vssd1 vssd1 vccd1 vccd1 _19549_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_53_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09302_ _09302_/A vssd1 vssd1 vccd1 vccd1 _09303_/B sky130_fd_sc_hd__inv_2
XFILLER_80_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09233_ _19883_/Q vssd1 vssd1 vccd1 vccd1 _09233_/Y sky130_fd_sc_hd__inv_2
XFILLER_221_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09164_ _09164_/A vssd1 vssd1 vccd1 vccd1 _09165_/A sky130_fd_sc_hd__inv_2
XFILLER_119_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17548__S _17548_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09095_ _20095_/Q _09084_/X _09094_/X _09087_/X vssd1 vssd1 vccd1 vccd1 _20095_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_72_HCLK_A clkbuf_opt_4_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19501__CLK _19510_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15893__A2 _16493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09997_ _09852_/A _09852_/B _09995_/Y _09990_/X vssd1 vssd1 vccd1 vccd1 _19943_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_131_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16688__A _16688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17283__S _17473_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08948_ _19853_/Q _08946_/Y _19861_/Q _08947_/Y vssd1 vssd1 vccd1 vccd1 _08948_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA_hold275_A sda_i_S4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10910_ _19684_/Q _10908_/Y _17936_/Q _10908_/A _15384_/A vssd1 vssd1 vccd1 vccd1
+ _19684_/D sky130_fd_sc_hd__o221a_1
XANTENNA__19036__RESET_B repeater267/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14001__A _18673_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11890_ _19423_/Q _11884_/X _09039_/X _11885_/X vssd1 vssd1 vccd1 vccd1 _19423_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_217_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14605__B1 _14604_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10841_ _10841_/A vssd1 vssd1 vccd1 vccd1 _14245_/D sky130_fd_sc_hd__buf_2
X_13560_ _13591_/A vssd1 vssd1 vccd1 vccd1 _13560_/X sky130_fd_sc_hd__buf_2
XFILLER_240_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10772_ _10773_/A vssd1 vssd1 vccd1 vccd1 _10772_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_44_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12511_ _19078_/Q _12505_/X _12410_/X _12506_/X vssd1 vssd1 vccd1 vccd1 _19078_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_201_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13491_ _18836_/Q vssd1 vssd1 vccd1 vccd1 _13491_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15030__B1 _15002_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15230_ _15205_/Y _15334_/B _15386_/A _15208_/A _15204_/X vssd1 vssd1 vccd1 vccd1
+ _15231_/A sky130_fd_sc_hd__o32a_1
XFILLER_200_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12442_ _12478_/A vssd1 vssd1 vccd1 vccd1 _12479_/A sky130_fd_sc_hd__inv_2
XANTENNA__11198__A2 _11191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18671__RESET_B repeater252/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15161_ _17952_/Q _15158_/X _14699_/A _15160_/X vssd1 vssd1 vccd1 vccd1 _17952_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17458__S _17546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12373_ _12427_/A vssd1 vssd1 vccd1 vccd1 _12400_/A sky130_fd_sc_hd__buf_2
X_14112_ _14112_/A vssd1 vssd1 vccd1 vccd1 _14112_/X sky130_fd_sc_hd__buf_2
X_11324_ _18960_/Q vssd1 vssd1 vccd1 vccd1 _11324_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15092_ _17995_/Q _15084_/A _09339_/X _15085_/A vssd1 vssd1 vccd1 vccd1 _17995_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18749__CLK _19900_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14043_ _19090_/Q vssd1 vssd1 vccd1 vccd1 _14043_/Y sky130_fd_sc_hd__inv_2
X_18920_ _19290_/CLK _18920_/D repeater211/X vssd1 vssd1 vccd1 vccd1 _18920_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_141_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11255_ _19586_/Q vssd1 vssd1 vccd1 vccd1 _11467_/A sky130_fd_sc_hd__inv_2
XFILLER_69_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10158__B1 _09086_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_192_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10206_ _19840_/Q vssd1 vssd1 vccd1 vccd1 _10206_/Y sky130_fd_sc_hd__inv_2
X_18851_ _18866_/CLK _18851_/D repeater232/X vssd1 vssd1 vccd1 vccd1 _18851_/Q sky130_fd_sc_hd__dfrtp_4
X_11186_ _17710_/X _11184_/X _19621_/Q _11185_/X vssd1 vssd1 vccd1 vccd1 _19621_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_68_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11370__A2 _19130_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17193__S _17548_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17802_ _18354_/Q _17994_/Q _18410_/Q _18394_/Q _17918_/S0 _18750_/Q vssd1 vssd1
+ vccd1 vccd1 _17802_/X sky130_fd_sc_hd__mux4_2
X_10137_ _17919_/X _08917_/A _10138_/A _19904_/Q _10136_/X vssd1 vssd1 vccd1 vccd1
+ _19904_/D sky130_fd_sc_hd__a32o_1
XFILLER_122_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18782_ _19855_/CLK _18782_/D repeater265/X vssd1 vssd1 vccd1 vccd1 _18782_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_209_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15994_ _16637_/A vssd1 vssd1 vccd1 vccd1 _16513_/A sky130_fd_sc_hd__buf_2
XFILLER_248_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17733_ _15376_/X _19712_/Q _18508_/D vssd1 vssd1 vccd1 vccd1 _17733_/X sky130_fd_sc_hd__mux2_1
X_10068_ _10068_/A vssd1 vssd1 vccd1 vccd1 _10068_/Y sky130_fd_sc_hd__inv_2
X_14945_ _18086_/Q _14939_/X _14929_/X _14941_/X vssd1 vssd1 vccd1 vccd1 _18086_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_235_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_235_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17664_ _15577_/Y _19025_/Q _17664_/S vssd1 vssd1 vccd1 vccd1 _18588_/D sky130_fd_sc_hd__mux2_1
XFILLER_75_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14876_ _18127_/Q _14871_/X _14705_/X _14873_/X vssd1 vssd1 vccd1 vccd1 _18127_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_211_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19403_ _19984_/CLK _19403_/D repeater243/X vssd1 vssd1 vccd1 vccd1 _19403_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_235_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16615_ _16615_/A _16615_/B vssd1 vssd1 vccd1 vccd1 _16615_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09005__A _19500_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13827_ _13914_/B _13827_/B vssd1 vssd1 vccd1 vccd1 _13921_/A sky130_fd_sc_hd__or2_1
X_17595_ _15346_/X _19708_/Q _17600_/S vssd1 vssd1 vccd1 vccd1 _17595_/X sky130_fd_sc_hd__mux2_1
XFILLER_90_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19334_ _19952_/CLK _19334_/D repeater244/X vssd1 vssd1 vccd1 vccd1 _19334_/Q sky130_fd_sc_hd__dfrtp_1
X_16546_ _16546_/A _16583_/B vssd1 vssd1 vccd1 vccd1 _16546_/Y sky130_fd_sc_hd__nor2_1
X_13758_ _13745_/Y _13760_/B _13757_/A _17763_/S _13757_/Y vssd1 vssd1 vccd1 vccd1
+ _13758_/X sky130_fd_sc_hd__a32o_1
XFILLER_62_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_188_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18759__RESET_B repeater195/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12709_ _12710_/A vssd1 vssd1 vccd1 vccd1 _12709_/X sky130_fd_sc_hd__clkbuf_2
X_19265_ _19952_/CLK _19265_/D repeater245/X vssd1 vssd1 vccd1 vccd1 _19265_/Q sky130_fd_sc_hd__dfrtp_4
X_16477_ _17103_/X _16594_/A _17105_/X _16595_/A vssd1 vssd1 vccd1 vccd1 _16481_/A
+ sky130_fd_sc_hd__a22oi_1
X_13689_ _18769_/Q _13685_/X _13678_/X _13686_/Y vssd1 vssd1 vccd1 vccd1 _18769_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18279__CLK _19847_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15021__B1 _15020_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18216_ _18216_/CLK _18216_/D vssd1 vssd1 vccd1 vccd1 _18216_/Q sky130_fd_sc_hd__dfxtp_1
X_15428_ _19619_/Q _11164_/B _11165_/B vssd1 vssd1 vccd1 vccd1 _15428_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__14375__A2 _14368_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19196_ _19222_/CLK _19196_/D repeater188/X vssd1 vssd1 vccd1 vccd1 _19196_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_163_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17368__S _17548_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15359_ _18501_/Q _14231_/B _14232_/B vssd1 vssd1 vccd1 vccd1 _15359_/X sky130_fd_sc_hd__a21bo_1
X_18147_ _18165_/CLK _18147_/D vssd1 vssd1 vccd1 vccd1 _18147_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold204 hold204/A vssd1 vssd1 vccd1 vccd1 hold204/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold215 hold215/A vssd1 vssd1 vccd1 vccd1 hold215/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold226 hold226/A vssd1 vssd1 vccd1 vccd1 hold226/X sky130_fd_sc_hd__dlygate4sd3_1
X_18078_ _18137_/CLK _18078_/D vssd1 vssd1 vccd1 vccd1 _18078_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_171_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold237 input66/X vssd1 vssd1 vccd1 vccd1 hold237/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold248 input67/X vssd1 vssd1 vccd1 vccd1 hold248/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09920_ _09853_/A _19336_/Q _19942_/Q _09917_/Y _09919_/X vssd1 vssd1 vccd1 vccd1
+ _09928_/B sky130_fd_sc_hd__o221a_1
X_17029_ _16666_/Y _19085_/Q _17490_/S vssd1 vssd1 vccd1 vccd1 _17029_/X sky130_fd_sc_hd__mux2_1
Xhold259 hold259/A vssd1 vssd1 vccd1 vccd1 hold259/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11346__C1 _11345_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20040_ _20051_/CLK _20040_/D repeater209/X vssd1 vssd1 vccd1 vccd1 _20040_/Q sky130_fd_sc_hd__dfrtp_1
X_09851_ _09851_/A _09998_/A vssd1 vssd1 vccd1 vccd1 _09852_/B sky130_fd_sc_hd__or2_2
XANTENNA__11897__B1 _09051_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15088__B1 hold244/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09782_ _19987_/Q _09781_/Y _09731_/A _09744_/B vssd1 vssd1 vccd1 vccd1 _19987_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__14835__B1 _14802_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_227_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11445__A _19155_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20031__CLK _20115_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09216_ _19887_/Q _15715_/A _19887_/Q _15715_/A vssd1 vssd1 vccd1 vccd1 _09242_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_10_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17278__S _17547_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09147_ _13494_/A _15321_/B hold344/X _09146_/Y vssd1 vssd1 vccd1 vccd1 _09151_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_108_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09078_ _20100_/Q _09069_/X _09077_/X _09072_/X vssd1 vssd1 vccd1 vccd1 _20100_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_151_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16910__S _17522_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19970__RESET_B hold370/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11040_ _11040_/A vssd1 vssd1 vccd1 vccd1 _11043_/A sky130_fd_sc_hd__inv_2
XFILLER_1_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11888__B1 hold305/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15079__B1 hold263/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_190_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14826__B1 _14791_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12991_ _12991_/A vssd1 vssd1 vccd1 vccd1 _12991_/Y sky130_fd_sc_hd__inv_2
XFILLER_217_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17741__S _18508_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11355__A _18980_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11942_ _11956_/A vssd1 vssd1 vccd1 vccd1 _11942_/X sky130_fd_sc_hd__buf_1
X_14730_ _18210_/Q _14718_/A _14693_/X _14719_/A vssd1 vssd1 vccd1 vccd1 _18210_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_245_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_217_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14661_ _18247_/Q _14656_/X _14606_/X _14658_/X vssd1 vssd1 vccd1 vccd1 _18247_/D
+ sky130_fd_sc_hd__a22o_1
X_11873_ _15772_/A _11998_/A vssd1 vssd1 vccd1 vccd1 _11914_/A sky130_fd_sc_hd__or2_2
XFILLER_189_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13612_ _18804_/Q _13445_/A _13591_/A _13610_/A vssd1 vssd1 vccd1 vccd1 _18804_/D
+ sky130_fd_sc_hd__o211a_1
X_16400_ _18033_/Q vssd1 vssd1 vccd1 vccd1 _16400_/Y sky130_fd_sc_hd__inv_2
X_10824_ _10446_/A _17750_/X _17750_/S _19724_/Q _10823_/Y vssd1 vssd1 vccd1 vccd1
+ _19724_/D sky130_fd_sc_hd__a32o_1
X_14592_ _18287_/Q _14587_/X _14537_/X _14589_/X vssd1 vssd1 vccd1 vccd1 _18287_/D
+ sky130_fd_sc_hd__a22o_1
X_17380_ _16216_/Y _15463_/A _17518_/S vssd1 vssd1 vccd1 vccd1 _17380_/X sky130_fd_sc_hd__mux2_1
XFILLER_220_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18852__RESET_B repeater232/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13543_ _13543_/A _13543_/B vssd1 vssd1 vccd1 vccd1 _13583_/A sky130_fd_sc_hd__or2_1
X_16331_ _18120_/Q vssd1 vssd1 vccd1 vccd1 _16331_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10755_ _11648_/A vssd1 vssd1 vccd1 vccd1 _15283_/A sky130_fd_sc_hd__inv_2
XANTENNA__11812__B1 _09064_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_198_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15003__B1 _15002_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11090__A _15318_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19050_ _19576_/CLK _19050_/D repeater255/X vssd1 vssd1 vccd1 vccd1 _19050_/Q sky130_fd_sc_hd__dfrtp_1
X_16262_ _18151_/Q vssd1 vssd1 vccd1 vccd1 _16262_/Y sky130_fd_sc_hd__inv_2
X_13474_ _18846_/Q _13473_/Y _13470_/B _13443_/X vssd1 vssd1 vccd1 vccd1 _18846_/D
+ sky130_fd_sc_hd__o211a_1
X_10686_ _15858_/C _15829_/B _10686_/C vssd1 vssd1 vccd1 vccd1 _15839_/A sky130_fd_sc_hd__or3_4
X_15213_ _15213_/A _15213_/B vssd1 vssd1 vccd1 vccd1 _15213_/X sky130_fd_sc_hd__or2_1
XFILLER_145_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18001_ _18412_/CLK _18001_/D vssd1 vssd1 vccd1 vccd1 _18001_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13565__B1 _13597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17188__S _17546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12425_ _19134_/Q _12420_/X _12225_/X _12421_/X vssd1 vssd1 vccd1 vccd1 _19134_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12368__B2 _12335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16193_ _18102_/Q vssd1 vssd1 vccd1 vccd1 _16193_/Y sky130_fd_sc_hd__inv_2
X_15144_ _17961_/Q _15135_/A _09255_/X _15136_/A vssd1 vssd1 vccd1 vccd1 _17961_/D
+ sky130_fd_sc_hd__a22o_1
X_12356_ hold251/X vssd1 vssd1 vccd1 vccd1 _12356_/X sky130_fd_sc_hd__clkbuf_4
X_11307_ _19596_/Q _11304_/Y _11481_/A _18983_/Q _11306_/X vssd1 vssd1 vccd1 vccd1
+ _11315_/B sky130_fd_sc_hd__o221a_1
X_15075_ _18008_/Q _15071_/X hold236/X _15073_/X vssd1 vssd1 vccd1 vccd1 _18008_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_113_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19952_ _19952_/CLK _19952_/D repeater244/X vssd1 vssd1 vccd1 vccd1 _19952_/Q sky130_fd_sc_hd__dfrtp_1
X_12287_ _19207_/Q _12283_/X _12028_/X _12284_/X vssd1 vssd1 vccd1 vccd1 _19207_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16820__S _17541_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_206_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17059__A1 _20115_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14026_ _14026_/A _14026_/B vssd1 vssd1 vccd1 vccd1 _14108_/A sky130_fd_sc_hd__or2_1
X_18903_ _18908_/CLK _18903_/D hold372/X vssd1 vssd1 vccd1 vccd1 _18903_/Q sky130_fd_sc_hd__dfrtp_1
X_11238_ _19014_/Q vssd1 vssd1 vccd1 vccd1 _16643_/A sky130_fd_sc_hd__inv_2
XFILLER_68_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11879__B1 _09016_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19883_ _20050_/CLK _19883_/D repeater200/X vssd1 vssd1 vccd1 vccd1 _19883_/Q sky130_fd_sc_hd__dfrtp_1
X_18834_ _19255_/CLK _18834_/D repeater239/X vssd1 vssd1 vccd1 vccd1 _18834_/Q sky130_fd_sc_hd__dfrtp_1
X_11169_ _19624_/Q _11169_/B vssd1 vssd1 vccd1 vccd1 _11170_/B sky130_fd_sc_hd__or2_1
XFILLER_68_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18765_ _18765_/CLK _18765_/D repeater196/X vssd1 vssd1 vccd1 vccd1 _18765_/Q sky130_fd_sc_hd__dfrtp_1
X_15977_ _15974_/Y _15831_/A _15975_/Y _15976_/X vssd1 vssd1 vccd1 vccd1 _15977_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_209_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17651__S _17655_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17716_ _15424_/X _19525_/Q _18546_/D vssd1 vssd1 vccd1 vccd1 _17716_/X sky130_fd_sc_hd__mux2_1
X_14928_ _18095_/Q _14920_/X _14927_/X _14923_/X vssd1 vssd1 vccd1 vccd1 _18095_/D
+ sky130_fd_sc_hd__a22o_1
X_18696_ _18701_/CLK _18696_/D hold351/X vssd1 vssd1 vccd1 vccd1 _18696_/Q sky130_fd_sc_hd__dfrtp_1
X_17647_ _15647_/Y _19042_/Q _17655_/S vssd1 vssd1 vccd1 vccd1 _18605_/D sky130_fd_sc_hd__mux2_1
X_14859_ _14859_/A vssd1 vssd1 vccd1 vccd1 _14860_/A sky130_fd_sc_hd__inv_2
XFILLER_51_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17578_ _15403_/X _19765_/Q _17584_/S vssd1 vssd1 vccd1 vccd1 _17578_/X sky130_fd_sc_hd__mux2_1
X_19317_ _19324_/CLK _19317_/D repeater214/X vssd1 vssd1 vccd1 vccd1 _19317_/Q sky130_fd_sc_hd__dfrtp_2
X_16529_ _17137_/X _16508_/X _17126_/X _16235_/X _16528_/X vssd1 vssd1 vccd1 vccd1
+ _16529_/X sky130_fd_sc_hd__o221a_1
XANTENNA__11803__B1 hold300/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19248_ _19320_/CLK _19248_/D repeater214/X vssd1 vssd1 vccd1 vccd1 _19248_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_192_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12359__A1 _19166_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09001_ _19497_/Q vssd1 vssd1 vccd1 vccd1 _15821_/B sky130_fd_sc_hd__inv_2
XFILLER_164_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17098__S _17518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19179_ _19288_/CLK _19179_/D repeater212/X vssd1 vssd1 vccd1 vccd1 _19179_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__19799__RESET_B repeater222/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17917__S0 _17918_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_191_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19728__RESET_B repeater207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09903_ _09877_/A _19361_/Q _19969_/Q _09900_/Y _09902_/X vssd1 vssd1 vccd1 vccd1
+ _09911_/B sky130_fd_sc_hd__o221a_1
XFILLER_132_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19381__RESET_B repeater230/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20023_ _20091_/CLK _20023_/D repeater236/X vssd1 vssd1 vccd1 vccd1 _20023_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__13655__A _15199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09834_ _19952_/Q vssd1 vssd1 vccd1 vccd1 _09860_/A sky130_fd_sc_hd__inv_2
XFILLER_112_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_246_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09765_ _09765_/A vssd1 vssd1 vccd1 vccd1 _09765_/Y sky130_fd_sc_hd__inv_2
XFILLER_246_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17561__S _17566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12295__B1 _12225_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_227_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09696_ _09793_/A _19410_/Q _19981_/Q _09694_/Y _09695_/X vssd1 vssd1 vccd1 vccd1
+ _09703_/B sky130_fd_sc_hd__o221a_1
XPHY_4016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer30 _13069_/C vssd1 vssd1 vccd1 vccd1 _13200_/A sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_242_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer41 _14013_/B vssd1 vssd1 vccd1 vccd1 _14132_/A sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_227_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrebuffer52 _09859_/B vssd1 vssd1 vccd1 vccd1 _09983_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_4049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer63 _13539_/B vssd1 vssd1 vccd1 vccd1 _13593_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14036__A1 _19069_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrebuffer74 _13073_/B vssd1 vssd1 vccd1 vccd1 _13194_/C1 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrebuffer85 _11463_/B vssd1 vssd1 vccd1 vccd1 _11537_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_230_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13390__A _20111_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer96 _13537_/C vssd1 vssd1 vccd1 vccd1 _13596_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12047__B1 _11918_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold140_A HADDR[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_hold238_A HWDATA[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16905__S _17542_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10540_ _10933_/A vssd1 vssd1 vccd1 vccd1 _10909_/A sky130_fd_sc_hd__buf_2
XPHY_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrebuffer120 _14031_/B vssd1 vssd1 vccd1 vccd1 _14101_/A sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_6_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10471_ _10471_/A vssd1 vssd1 vccd1 vccd1 _10471_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__17908__S0 _17908_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12210_ _19245_/Q _12205_/X _12102_/X _12206_/X vssd1 vssd1 vccd1 vccd1 _19245_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17289__A1 _09424_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16743__A_N _16682_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13190_ _13190_/A vssd1 vssd1 vccd1 vccd1 _13190_/Y sky130_fd_sc_hd__inv_2
XFILLER_203_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19469__RESET_B repeater274/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_191_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17736__S _18508_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12141_ _19290_/Q _12134_/X _12078_/X _12137_/X vssd1 vssd1 vccd1 vccd1 _19290_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_163_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12072_ _12096_/A vssd1 vssd1 vccd1 vccd1 _12072_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_150_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11023_ _19650_/Q vssd1 vssd1 vccd1 vccd1 _11023_/Y sky130_fd_sc_hd__inv_2
X_15900_ _15900_/A vssd1 vssd1 vccd1 vccd1 _15901_/A sky130_fd_sc_hd__clkbuf_2
X_16880_ _16879_/X _09426_/Y _17413_/S vssd1 vssd1 vccd1 vccd1 _16880_/X sky130_fd_sc_hd__mux2_1
X_15831_ _15831_/A vssd1 vssd1 vccd1 vccd1 _15850_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_66_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17471__S _17567_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18550_ _19825_/CLK _18550_/D repeater223/X vssd1 vssd1 vccd1 vccd1 _18550_/Q sky130_fd_sc_hd__dfrtp_1
X_15762_ _15765_/C _15762_/B _18527_/Q vssd1 vssd1 vccd1 vccd1 _18523_/D sky130_fd_sc_hd__nor3_1
XFILLER_18_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12286__B1 _12026_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12974_ _18945_/Q _12970_/C _12962_/X _12972_/A vssd1 vssd1 vccd1 vccd1 _18945_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_57_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17501_ _17500_/X _08946_/Y _17566_/S vssd1 vssd1 vccd1 vccd1 _17501_/X sky130_fd_sc_hd__mux2_1
X_14713_ _14713_/A vssd1 vssd1 vccd1 vccd1 _14713_/X sky130_fd_sc_hd__clkbuf_2
X_18481_ _19545_/CLK _18481_/D repeater225/X vssd1 vssd1 vccd1 vccd1 _18481_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_61_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11925_ _19402_/Q _11891_/A _11924_/X _11892_/A vssd1 vssd1 vccd1 vccd1 _19402_/D
+ sky130_fd_sc_hd__a22o_1
X_15693_ _15693_/A vssd1 vssd1 vccd1 vccd1 _15693_/Y sky130_fd_sc_hd__inv_2
XANTENNA_output112_A _16747_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17432_ _17431_/X _15194_/Y _17567_/S vssd1 vssd1 vccd1 vccd1 _17432_/X sky130_fd_sc_hd__mux2_1
XPHY_4583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16972__A0 _15963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11856_ _11856_/A _15201_/B vssd1 vssd1 vccd1 vccd1 _11856_/Y sky130_fd_sc_hd__nor2_1
X_14644_ _14644_/A vssd1 vssd1 vccd1 vccd1 _14645_/A sky130_fd_sc_hd__inv_2
XPHY_4594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10807_ _10807_/A _17621_/S vssd1 vssd1 vccd1 vccd1 _10809_/A sky130_fd_sc_hd__nand2_2
XFILLER_220_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14575_ _18297_/Q _14572_/X _14531_/X _14574_/X vssd1 vssd1 vccd1 vccd1 _18297_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17363_ _15768_/Y _14204_/Y _17546_/S vssd1 vssd1 vccd1 vccd1 _17363_/X sky130_fd_sc_hd__mux2_1
XPHY_3893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09444__A2_N _19380_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11787_ _11801_/A vssd1 vssd1 vccd1 vccd1 _11787_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__16815__S _17545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19102_ _19585_/CLK _19102_/D hold361/X vssd1 vssd1 vccd1 vccd1 _19102_/Q sky130_fd_sc_hd__dfrtp_1
X_16314_ _19770_/Q vssd1 vssd1 vccd1 vccd1 _16314_/Y sky130_fd_sc_hd__inv_2
XFILLER_158_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10738_ _18550_/Q _15270_/C _11648_/A _15271_/D vssd1 vssd1 vccd1 vccd1 _10738_/X
+ sky130_fd_sc_hd__a211o_1
X_13526_ _13500_/Y _13509_/X _13513_/Y _13518_/Y _13525_/X vssd1 vssd1 vccd1 vccd1
+ _13526_/X sky130_fd_sc_hd__a2111o_1
XANTENNA__15939__B _16344_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17294_ _17486_/A0 _13123_/Y _17543_/S vssd1 vssd1 vccd1 vccd1 _17294_/X sky130_fd_sc_hd__mux2_1
XFILLER_158_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10148__B _19515_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_185_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19033_ _19577_/CLK _19033_/D repeater267/X vssd1 vssd1 vccd1 vccd1 _19033_/Q sky130_fd_sc_hd__dfrtp_1
X_13457_ _18852_/Q _13456_/Y _13340_/B _13443_/X vssd1 vssd1 vccd1 vccd1 _18852_/D
+ sky130_fd_sc_hd__o211a_1
X_16245_ _16494_/A vssd1 vssd1 vccd1 vccd1 _16594_/A sky130_fd_sc_hd__inv_2
X_10669_ _10676_/A vssd1 vssd1 vccd1 vccd1 _10669_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_opt_0_HCLK_A clkbuf_opt_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19892__RESET_B repeater205/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12644__A _12651_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12408_ hold310/X vssd1 vssd1 vccd1 vccd1 _12408_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__12210__B1 _12102_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13388_ _20095_/Q _13464_/A _20119_/Q _13387_/Y vssd1 vssd1 vccd1 vccd1 _13388_/X
+ sky130_fd_sc_hd__a22o_1
X_16176_ _18246_/Q _16344_/B vssd1 vssd1 vccd1 vccd1 _16176_/Y sky130_fd_sc_hd__nand2_1
XFILLER_127_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput106 _16327_/Y vssd1 vssd1 vccd1 vccd1 HRDATA[5] sky130_fd_sc_hd__clkbuf_2
Xoutput117 _16757_/LO vssd1 vssd1 vccd1 vccd1 IRQ[14] sky130_fd_sc_hd__clkbuf_2
XANTENNA__17646__S _17655_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput128 _19749_/Q vssd1 vssd1 vccd1 vccd1 MSO_S2 sky130_fd_sc_hd__clkbuf_2
X_15127_ _17974_/Q _15122_/X _14927_/X _15124_/X vssd1 vssd1 vccd1 vccd1 _17974_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_5_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12339_ _19176_/Q _12334_/X _12102_/X _12335_/X vssd1 vssd1 vccd1 vccd1 _19176_/D
+ sky130_fd_sc_hd__a22o_1
Xoutput139 _16760_/LO vssd1 vssd1 vccd1 vccd1 scl_o_S5 sky130_fd_sc_hd__clkbuf_2
XFILLER_142_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19139__RESET_B repeater274/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19935_ _19937_/CLK _19935_/D repeater189/X vssd1 vssd1 vccd1 vccd1 _19935_/Q sky130_fd_sc_hd__dfrtp_1
X_15058_ _15058_/A _19850_/Q _15058_/C vssd1 vssd1 vccd1 vccd1 _15060_/A sky130_fd_sc_hd__or3_4
XFILLER_142_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14009_ _14009_/A _14009_/B vssd1 vssd1 vccd1 vccd1 _14139_/A sky130_fd_sc_hd__or2_1
X_19866_ _19867_/CLK _19866_/D repeater263/X vssd1 vssd1 vccd1 vccd1 _19866_/Q sky130_fd_sc_hd__dfrtp_1
X_18817_ _18856_/CLK _18817_/D repeater231/X vssd1 vssd1 vccd1 vccd1 _18817_/Q sky130_fd_sc_hd__dfrtp_1
X_19797_ _19808_/CLK _19797_/D repeater224/X vssd1 vssd1 vccd1 vccd1 _19797_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_244_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17381__S _17517_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09550_ _20008_/Q _16212_/A _09468_/A _19297_/Q _09549_/X vssd1 vssd1 vccd1 vccd1
+ _09564_/A sky130_fd_sc_hd__o221a_1
XFILLER_209_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18748_ _20036_/CLK _18748_/D repeater198/X vssd1 vssd1 vccd1 vccd1 _18748_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_36_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17204__A1 _09436_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10827__A1 _10698_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09481_ _09481_/A _09592_/A vssd1 vssd1 vccd1 vccd1 _09482_/B sky130_fd_sc_hd__or2_2
XFILLER_224_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18679_ _18686_/CLK _18679_/D repeater252/X vssd1 vssd1 vccd1 vccd1 _18679_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_36_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18703__RESET_B hold351/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11723__A _11730_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12029__B1 _12028_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_205_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_220_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12201__B1 _12086_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17556__S _19498_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_127_HCLK_A clkbuf_4_4_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20006_ _20006_/CLK _20006_/D repeater240/X vssd1 vssd1 vccd1 vccd1 _20006_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_59_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16246__A2 _16597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09817_ _19969_/Q vssd1 vssd1 vccd1 vccd1 _09877_/A sky130_fd_sc_hd__inv_2
XFILLER_100_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17291__S _17512_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12268__B1 _12080_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09748_ _09748_/A _09748_/B vssd1 vssd1 vccd1 vccd1 _09772_/A sky130_fd_sc_hd__or2_1
XANTENNA__10818__A1 _20036_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09679_ _09646_/C _19412_/Q _19983_/Q _09676_/Y _09678_/X vssd1 vssd1 vccd1 vccd1
+ _09689_/B sky130_fd_sc_hd__o221a_1
XPHY_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11710_ _11738_/A vssd1 vssd1 vccd1 vccd1 _11731_/A sky130_fd_sc_hd__buf_2
XPHY_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12690_ _18972_/Q _12684_/X _12032_/A _12685_/X vssd1 vssd1 vccd1 vccd1 _18972_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_199_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11641_ _11641_/A _11641_/B _11645_/C vssd1 vssd1 vccd1 vccd1 _19549_/D sky130_fd_sc_hd__nor3_1
XPHY_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09103__A hold336/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14360_ _18423_/Q _14349_/X _14359_/X _14353_/X vssd1 vssd1 vccd1 vccd1 _18423_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_23_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11572_ _11572_/A _11615_/A vssd1 vssd1 vccd1 vccd1 _11573_/B sky130_fd_sc_hd__or2_2
XPHY_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13311_ _18854_/Q vssd1 vssd1 vccd1 vccd1 _13429_/B sky130_fd_sc_hd__inv_2
XFILLER_210_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10523_ _10735_/A vssd1 vssd1 vccd1 vccd1 _10527_/A sky130_fd_sc_hd__inv_2
Xinput19 HADDR[26] vssd1 vssd1 vccd1 vccd1 input19/X sky130_fd_sc_hd__buf_1
XPHY_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14291_ _18457_/Q _14288_/X _14273_/X _14290_/X vssd1 vssd1 vccd1 vccd1 _18457_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12464__A _12478_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_182_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13242_ _13242_/A vssd1 vssd1 vccd1 vccd1 _13243_/A sky130_fd_sc_hd__inv_2
XFILLER_6_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16030_ _18268_/Q vssd1 vssd1 vccd1 vccd1 _16030_/Y sky130_fd_sc_hd__inv_2
X_10454_ _19830_/Q _10450_/X _10418_/X _10452_/X vssd1 vssd1 vccd1 vccd1 _19830_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13279__B _19517_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_142_HCLK clkbuf_4_3_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _18465_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_184_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17466__S _17567_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13173_ _18912_/Q _13172_/Y _13162_/X _13173_/C1 vssd1 vssd1 vccd1 vccd1 _18912_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_124_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10385_ _19853_/Q _19852_/Q _08921_/X _08964_/X vssd1 vssd1 vccd1 vccd1 _10385_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_151_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12124_ _19299_/Q _12121_/X _11981_/X _12122_/X vssd1 vssd1 vccd1 vccd1 _19299_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19735__CLK _20051_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17981_ _20124_/CLK _17981_/D vssd1 vssd1 vccd1 vccd1 _17981_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19720_ _19720_/CLK _19720_/D repeater202/X vssd1 vssd1 vccd1 vccd1 _19720_/Q sky130_fd_sc_hd__dfrtp_1
X_12055_ _17611_/X _12055_/B vssd1 vssd1 vccd1 vccd1 _12056_/A sky130_fd_sc_hd__or2_2
X_16932_ _19476_/Q hold183/X _16946_/S vssd1 vssd1 vccd1 vccd1 _16932_/X sky130_fd_sc_hd__mux2_2
XANTENNA__10712__A hold322/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_238_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11006_ _19658_/Q _11006_/B vssd1 vssd1 vccd1 vccd1 _11006_/Y sky130_fd_sc_hd__nor2_1
X_19651_ _19859_/CLK _19651_/D repeater261/X vssd1 vssd1 vccd1 vccd1 _19651_/Q sky130_fd_sc_hd__dfrtp_1
X_16863_ _16862_/X _15648_/Y _17318_/S vssd1 vssd1 vccd1 vccd1 _16863_/X sky130_fd_sc_hd__mux2_1
XFILLER_238_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10431__B _16053_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_49_HCLK_A clkbuf_opt_2_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18602_ _19867_/CLK _18602_/D repeater263/X vssd1 vssd1 vccd1 vccd1 _18602_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_65_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15814_ _17953_/Q vssd1 vssd1 vccd1 vccd1 _15814_/Y sky130_fd_sc_hd__inv_2
X_19582_ _19582_/CLK _19582_/D hold348/A vssd1 vssd1 vccd1 vccd1 _19582_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__15996__A1 _17482_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16794_ _16717_/Y _19090_/Q _17544_/S vssd1 vssd1 vccd1 vccd1 _16794_/X sky130_fd_sc_hd__mux2_1
XANTENNA__15996__B2 _16513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18533_ _19771_/CLK _18533_/D repeater189/X vssd1 vssd1 vccd1 vccd1 _18533_/Q sky130_fd_sc_hd__dfrtp_1
X_15745_ _18483_/Q _18484_/Q _18485_/Q vssd1 vssd1 vccd1 vccd1 _18483_/D sky130_fd_sc_hd__o21ba_1
XFILLER_234_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12957_ _12968_/B vssd1 vssd1 vccd1 vccd1 _13060_/B sky130_fd_sc_hd__inv_2
XFILLER_45_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18464_ _18465_/CLK _18464_/D vssd1 vssd1 vccd1 vccd1 _18464_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13208__C1 _13176_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11908_ _19411_/Q _11905_/X _09075_/X _11906_/X vssd1 vssd1 vccd1 vccd1 _19411_/D
+ sky130_fd_sc_hd__a22o_1
X_15676_ _18612_/Q _15678_/B vssd1 vssd1 vccd1 vccd1 _15681_/B sky130_fd_sc_hd__or2_1
XPHY_4380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12888_ _12888_/A _12888_/B _12972_/A vssd1 vssd1 vccd1 vccd1 _12889_/A sky130_fd_sc_hd__or3_4
XPHY_4391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17415_ _15963_/X _12810_/Y _17534_/S vssd1 vssd1 vccd1 vccd1 _17415_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09013__A _12187_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14627_ _18266_/Q _14617_/A _14626_/X _14618_/A vssd1 vssd1 vccd1 vccd1 _18266_/D
+ sky130_fd_sc_hd__a22o_1
X_18395_ _18412_/CLK _18395_/D vssd1 vssd1 vccd1 vccd1 _18395_/Q sky130_fd_sc_hd__dfxtp_1
X_11839_ _12558_/B _15776_/A vssd1 vssd1 vccd1 vccd1 _11840_/S sky130_fd_sc_hd__or2_2
XANTENNA__09427__B2 _09426_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17346_ _16344_/X _18232_/Q _17564_/S vssd1 vssd1 vccd1 vccd1 _17346_/X sky130_fd_sc_hd__mux2_1
X_14558_ _14559_/A vssd1 vssd1 vccd1 vccd1 _14558_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__12431__B1 _12232_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13509_ _14629_/B _13506_/Y _13523_/A vssd1 vssd1 vccd1 vccd1 _13509_/X sky130_fd_sc_hd__o21a_1
XANTENNA__12374__A _12400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17277_ _16484_/X _10213_/Y _17566_/S vssd1 vssd1 vccd1 vccd1 _17277_/X sky130_fd_sc_hd__mux2_1
X_14489_ _19849_/Q _14489_/B _15318_/B vssd1 vssd1 vccd1 vccd1 _15094_/C sky130_fd_sc_hd__or3_4
XFILLER_146_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19016_ _19115_/CLK _19016_/D hold353/X vssd1 vssd1 vccd1 vccd1 _19016_/Q sky130_fd_sc_hd__dfrtp_4
X_16228_ _19760_/Q vssd1 vssd1 vccd1 vccd1 _16228_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17376__S _17567_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16159_ _18054_/Q vssd1 vssd1 vccd1 vccd1 _16159_/Y sky130_fd_sc_hd__inv_2
XANTENNA__10745__B1 _10448_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16476__A2 _15915_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08981_ _18870_/Q _09198_/A _17601_/X vssd1 vssd1 vccd1 vccd1 _08981_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__15684__B1 _15673_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19918_ _19937_/CLK _19918_/D repeater230/X vssd1 vssd1 vccd1 vccd1 _19918_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_87_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18955__RESET_B repeater257/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19849_ _19849_/CLK _19849_/D repeater258/X vssd1 vssd1 vccd1 vccd1 _19849_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__14239__B2 _17600_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_228_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09602_ _20015_/Q _09604_/A _09585_/X _09602_/C1 vssd1 vssd1 vccd1 vccd1 _20015_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_110_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09533_ _20025_/Q _09529_/Y _20021_/Q _16587_/A _09532_/X vssd1 vssd1 vccd1 vccd1
+ _09545_/A sky130_fd_sc_hd__o221a_1
XFILLER_209_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_23_HCLK clkbuf_4_9_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20066_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_25_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09464_ _09394_/Y _09417_/Y _09464_/C _09464_/D vssd1 vssd1 vccd1 vccd1 _09465_/B
+ sky130_fd_sc_hd__nand4bb_4
XFILLER_64_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09395_ _19913_/Q vssd1 vssd1 vccd1 vccd1 _10085_/A sky130_fd_sc_hd__inv_2
XPHY_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_196_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12422__B1 _12353_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19743__RESET_B repeater207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17286__S _17544_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10170_ _19886_/Q _10166_/X _09079_/X _10168_/X vssd1 vssd1 vccd1 vccd1 _19886_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_121_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16203__B _16344_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14004__A _14004_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18696__RESET_B hold351/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13860_ _19214_/Q vssd1 vssd1 vccd1 vccd1 _13860_/Y sky130_fd_sc_hd__inv_2
XFILLER_47_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09106__B1 _09105_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12811_ _18816_/Q vssd1 vssd1 vccd1 vccd1 _13539_/A sky130_fd_sc_hd__inv_2
XFILLER_74_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_216_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13791_ _18721_/Q vssd1 vssd1 vccd1 vccd1 _13910_/B sky130_fd_sc_hd__inv_2
XFILLER_170_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20115__CLK _20115_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15530_ _15530_/A _15530_/B vssd1 vssd1 vccd1 vccd1 _15530_/Y sky130_fd_sc_hd__nor2_1
X_12742_ _18823_/Q vssd1 vssd1 vccd1 vccd1 _13546_/A sky130_fd_sc_hd__inv_2
XFILLER_27_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13281__C _15190_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12673_ _18985_/Q _12670_/X hold308/X _12671_/X vssd1 vssd1 vccd1 vccd1 _18985_/D
+ sky130_fd_sc_hd__a22o_1
X_15461_ _18560_/Q vssd1 vssd1 vccd1 vccd1 _15463_/A sky130_fd_sc_hd__inv_2
XANTENNA__09409__B2 _19395_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17200_ _15963_/X _12822_/Y _17534_/S vssd1 vssd1 vccd1 vccd1 _17200_/X sky130_fd_sc_hd__mux2_1
XPHY_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14412_ _18393_/Q _14409_/X _14351_/X _14411_/X vssd1 vssd1 vccd1 vccd1 _18393_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_8_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11624_ _11624_/A _11624_/B vssd1 vssd1 vccd1 vccd1 _11629_/A sky130_fd_sc_hd__or2_1
XPHY_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18180_ _18216_/CLK _18180_/D vssd1 vssd1 vccd1 vccd1 _18180_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15392_ _18529_/Q _18528_/Q _13217_/B vssd1 vssd1 vccd1 vccd1 _15392_/X sky130_fd_sc_hd__a21bo_1
XPHY_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19484__RESET_B repeater260/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17131_ _17130_/X _19207_/Q _17545_/S vssd1 vssd1 vccd1 vccd1 _17131_/X sky130_fd_sc_hd__mux2_2
X_11555_ _11577_/A _11576_/A _11578_/A _11575_/A vssd1 vssd1 vccd1 vccd1 _11556_/D
+ sky130_fd_sc_hd__or4_4
X_14343_ _18429_/Q _14336_/X _14326_/X _14338_/X vssd1 vssd1 vccd1 vccd1 _18429_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19413__RESET_B repeater193/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10506_ _19533_/Q vssd1 vssd1 vccd1 vccd1 _10508_/A sky130_fd_sc_hd__inv_2
XFILLER_144_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17062_ _17061_/X _11358_/Y _17493_/S vssd1 vssd1 vccd1 vccd1 _17062_/X sky130_fd_sc_hd__mux2_1
X_14274_ _14274_/A vssd1 vssd1 vccd1 vccd1 _14275_/A sky130_fd_sc_hd__inv_2
XFILLER_128_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11486_ _11486_/A _11486_/B vssd1 vssd1 vccd1 vccd1 _11494_/A sky130_fd_sc_hd__or2_1
X_13225_ _18538_/Q _13225_/B vssd1 vssd1 vccd1 vccd1 _13226_/B sky130_fd_sc_hd__or2_1
X_16013_ _18036_/Q vssd1 vssd1 vccd1 vccd1 _16013_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17196__S _17548_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10437_ _19840_/Q _10433_/X _09061_/X _10435_/X vssd1 vssd1 vccd1 vccd1 _19840_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18670__SET_B repeater222/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10727__B1 _10421_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13156_ _19159_/Q vssd1 vssd1 vccd1 vccd1 _13156_/Y sky130_fd_sc_hd__inv_2
XFILLER_151_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10368_ _10368_/A vssd1 vssd1 vccd1 vccd1 _10368_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_124_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12107_ hold277/X vssd1 vssd1 vccd1 vccd1 _12107_/X sky130_fd_sc_hd__clkbuf_4
X_17964_ _19842_/CLK _17964_/D vssd1 vssd1 vccd1 vccd1 _17964_/Q sky130_fd_sc_hd__dfxtp_1
X_13087_ _13087_/A _13087_/B vssd1 vssd1 vccd1 vccd1 _13166_/A sky130_fd_sc_hd__or2_1
X_10299_ _18594_/Q _15597_/A vssd1 vssd1 vccd1 vccd1 _15601_/A sky130_fd_sc_hd__or2_1
XFILLER_214_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19703_ _20055_/CLK _19703_/D repeater202/X vssd1 vssd1 vccd1 vccd1 _19703_/Q sky130_fd_sc_hd__dfstp_1
X_16915_ _17473_/A0 _16631_/Y _17042_/S vssd1 vssd1 vccd1 vccd1 _16915_/X sky130_fd_sc_hd__mux2_1
X_12038_ hold250/X vssd1 vssd1 vccd1 vccd1 _12038_/X sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_46_HCLK clkbuf_opt_2_HCLK/A vssd1 vssd1 vccd1 vccd1 _19814_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_clkbuf_leaf_110_HCLK_A clkbuf_opt_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_238_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17895_ _15940_/Y _15941_/Y _15942_/Y _15943_/Y _17908_/S0 _18759_/Q vssd1 vssd1
+ vccd1 vccd1 _17895_/X sky130_fd_sc_hd__mux4_2
XANTENNA__15418__B1 _17584_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19634_ _19851_/CLK _19634_/D repeater258/X vssd1 vssd1 vccd1 vccd1 _19634_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_66_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16846_ _16845_/X _12929_/Y _17487_/S vssd1 vssd1 vccd1 vccd1 _16846_/X sky130_fd_sc_hd__mux2_1
XFILLER_66_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_225_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15969__B2 _15867_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19565_ _19576_/CLK _19565_/D repeater255/X vssd1 vssd1 vccd1 vccd1 _19565_/Q sky130_fd_sc_hd__dfrtp_1
X_16777_ _16776_/X _09494_/A _17414_/S vssd1 vssd1 vccd1 vccd1 _16777_/X sky130_fd_sc_hd__mux2_1
X_13989_ _18685_/Q vssd1 vssd1 vccd1 vccd1 _14015_/A sky130_fd_sc_hd__inv_2
XFILLER_241_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18516_ _19825_/CLK _19755_/Q repeater229/X vssd1 vssd1 vccd1 vccd1 _18516_/Q sky130_fd_sc_hd__dfrtp_1
X_15728_ _20038_/Q vssd1 vssd1 vccd1 vccd1 _15728_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19496_ _19859_/CLK hold253/X repeater262/X vssd1 vssd1 vccd1 vccd1 _19496_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12652__B1 _12599_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_234_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_206_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18447_ _19855_/CLK _18447_/D vssd1 vssd1 vccd1 vccd1 _18447_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_221_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15659_ _18608_/Q vssd1 vssd1 vccd1 vccd1 _15661_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_178_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09180_ _14709_/A vssd1 vssd1 vccd1 vccd1 _09180_/X sky130_fd_sc_hd__clkbuf_2
X_18378_ _19515_/CLK _18378_/D vssd1 vssd1 vccd1 vccd1 _18378_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__19900__CLK _19900_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17329_ _17328_/X _13534_/A _17536_/S vssd1 vssd1 vccd1 vccd1 _17329_/X sky130_fd_sc_hd__mux2_2
XFILLER_174_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16146__B2 _15999_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18035__CLK _19851_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08964_ _10321_/B vssd1 vssd1 vccd1 vccd1 _08964_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_124_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15862__B _15863_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_229_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16606__C1 _16605_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18185__CLK _18198_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_32_HCLK_A _18641_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19995__RESET_B repeater192/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_95_HCLK_A clkbuf_4_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_213_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09516_ _20006_/Q _09513_/Y _09467_/A _19296_/Q _09515_/X vssd1 vssd1 vccd1 vccd1
+ _09516_/X sky130_fd_sc_hd__a221o_1
XFILLER_25_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19924__RESET_B repeater230/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09447_ _19911_/Q vssd1 vssd1 vccd1 vccd1 _10083_/A sky130_fd_sc_hd__inv_2
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_224_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11911__A hold260/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09378_ _10044_/A _19388_/Q _10042_/A _19386_/Q vssd1 vssd1 vccd1 vccd1 _09378_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_40_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16913__S _17385_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11340_ _11464_/A _18965_/Q _19581_/Q _11337_/Y _11339_/X vssd1 vssd1 vccd1 vccd1
+ _11347_/B sky130_fd_sc_hd__o221a_1
XFILLER_181_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11271_ _19009_/Q vssd1 vssd1 vccd1 vccd1 _16582_/A sky130_fd_sc_hd__inv_2
X_13010_ _13008_/A _13008_/B _13008_/Y _12986_/A vssd1 vssd1 vccd1 vccd1 _18929_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_3_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18877__RESET_B repeater208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10222_ _19839_/Q _10966_/A _10218_/Y _19654_/Q _10221_/X vssd1 vssd1 vccd1 vccd1
+ _10247_/C sky130_fd_sc_hd__o221a_1
XFILLER_152_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_69_HCLK clkbuf_opt_3_HCLK/A vssd1 vssd1 vccd1 vccd1 _18886_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__18806__RESET_B repeater231/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17744__S _18508_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11358__A _18991_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10153_ _12436_/C _10186_/B vssd1 vssd1 vccd1 vccd1 _10155_/A sky130_fd_sc_hd__or2_4
XFILLER_160_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10084_ _10084_/A _10084_/B vssd1 vssd1 vccd1 vccd1 _10094_/A sky130_fd_sc_hd__or2_1
XANTENNA_input36_A HTRANS[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14961_ _18075_/Q _14953_/A _14935_/X _14954_/A vssd1 vssd1 vccd1 vccd1 _18075_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_248_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16700_ _19052_/Q vssd1 vssd1 vccd1 vccd1 _16700_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13912_ _13912_/A _13912_/B _13912_/C _13912_/D vssd1 vssd1 vccd1 vccd1 _13914_/C
+ sky130_fd_sc_hd__or4_4
X_17680_ _15513_/X _19455_/Q _17683_/S vssd1 vssd1 vccd1 vccd1 _18572_/D sky130_fd_sc_hd__mux2_1
XFILLER_101_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14892_ _18115_/Q _14884_/A _14816_/X _14885_/A vssd1 vssd1 vccd1 vccd1 _18115_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_235_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_207_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16073__B1 _17467_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16631_ _19460_/Q vssd1 vssd1 vccd1 vccd1 _16631_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16612__A2 _15889_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13843_ _13837_/X _13839_/X _13843_/C _13843_/D vssd1 vssd1 vccd1 vccd1 _13850_/B
+ sky130_fd_sc_hd__nand4bb_2
XFILLER_223_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19350_ _19352_/CLK _19350_/D hold373/X vssd1 vssd1 vccd1 vccd1 _19350_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12634__B1 _12408_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16562_ _17114_/X _16505_/A _17124_/X _16506_/A vssd1 vssd1 vccd1 vccd1 _16562_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10986_ _10986_/A vssd1 vssd1 vccd1 vccd1 _19664_/D sky130_fd_sc_hd__inv_2
XFILLER_62_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13774_ _18737_/Q _18738_/Q _13775_/S vssd1 vssd1 vccd1 vccd1 _18738_/D sky130_fd_sc_hd__mux2_1
X_18301_ _18431_/CLK _18301_/D vssd1 vssd1 vccd1 vccd1 _18301_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17799__S1 _19648_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15513_ _15510_/Y _15511_/Y _15512_/X vssd1 vssd1 vccd1 vccd1 _15513_/X sky130_fd_sc_hd__o21a_1
XFILLER_188_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12725_ _18954_/Q vssd1 vssd1 vccd1 vccd1 _14814_/A sky130_fd_sc_hd__clkbuf_2
X_19281_ _19282_/CLK _19281_/D repeater216/X vssd1 vssd1 vccd1 vccd1 _19281_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_231_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16493_ _16493_/A vssd1 vssd1 vccd1 vccd1 _16493_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_repeater175_A _17513_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18232_ _18412_/CLK _18232_/D vssd1 vssd1 vccd1 vccd1 _18232_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11821__A _11821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_231_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15444_ _19399_/Q vssd1 vssd1 vccd1 vccd1 _15571_/A sky130_fd_sc_hd__inv_2
XPHY_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12656_ _18994_/Q _12650_/X _12538_/X _12651_/X vssd1 vssd1 vccd1 vccd1 _18994_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11607_ _19565_/Q _11606_/Y _11592_/X _11579_/B vssd1 vssd1 vccd1 vccd1 _19565_/D
+ sky130_fd_sc_hd__o211a_1
X_18163_ _18165_/CLK _18163_/D vssd1 vssd1 vccd1 vccd1 _18163_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15375_ _19791_/Q _10651_/B _10652_/B vssd1 vssd1 vccd1 vccd1 _15375_/X sky130_fd_sc_hd__a21bo_1
X_12587_ _19039_/Q _12583_/X hold281/X _12584_/X vssd1 vssd1 vccd1 vccd1 _19039_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16823__S _17529_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17114_ _16484_/X _08928_/Y _17566_/S vssd1 vssd1 vccd1 vccd1 _17114_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_184_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14326_ hold331/X vssd1 vssd1 vccd1 vccd1 _14326_/X sky130_fd_sc_hd__clkbuf_2
X_18094_ _20090_/CLK _18094_/D vssd1 vssd1 vccd1 vccd1 _18094_/Q sky130_fd_sc_hd__dfxtp_1
X_11538_ _11538_/A vssd1 vssd1 vccd1 vccd1 _11538_/Y sky130_fd_sc_hd__inv_2
XFILLER_128_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17045_ _17044_/X _15672_/Y _17318_/S vssd1 vssd1 vccd1 vccd1 _17045_/X sky130_fd_sc_hd__mux2_1
X_11469_ _11469_/A _11525_/A vssd1 vssd1 vccd1 vccd1 _11470_/B sky130_fd_sc_hd__or2_2
X_14257_ _14490_/A _14963_/B _15034_/C vssd1 vssd1 vccd1 vccd1 _14259_/A sky130_fd_sc_hd__or3_4
XFILLER_109_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13208_ _18892_/Q _13207_/Y _13208_/B1 _13176_/X vssd1 vssd1 vccd1 vccd1 _18892_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_131_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14188_ _19120_/Q _18699_/Q _14187_/Y _14029_/A vssd1 vssd1 vccd1 vccd1 _14193_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_124_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17654__S _17655_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15963__A _17539_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13139_ _19184_/Q _13085_/A _13135_/Y _18887_/Q _13138_/X vssd1 vssd1 vccd1 vccd1
+ _13144_/C sky130_fd_sc_hd__o221a_1
XFILLER_225_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18996_ _19137_/CLK _18996_/D repeater249/X vssd1 vssd1 vccd1 vccd1 _18996_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_86_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14311__B1 _13678_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater203 repeater204/X vssd1 vssd1 vccd1 vccd1 repeater203/X sky130_fd_sc_hd__buf_6
X_17947_ _18765_/CLK _17947_/D vssd1 vssd1 vccd1 vccd1 _17947_/Q sky130_fd_sc_hd__dfxtp_1
Xrepeater214 repeater215/X vssd1 vssd1 vccd1 vccd1 repeater214/X sky130_fd_sc_hd__buf_8
Xrepeater225 repeater227/X vssd1 vssd1 vccd1 vccd1 repeater225/X sky130_fd_sc_hd__buf_8
XFILLER_227_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13483__A _13483_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater236 repeater238/X vssd1 vssd1 vccd1 vccd1 repeater236/X sky130_fd_sc_hd__buf_8
Xrepeater247 hold371/A vssd1 vssd1 vccd1 vccd1 hold372/A sky130_fd_sc_hd__buf_4
Xrepeater258 repeater259/X vssd1 vssd1 vccd1 vccd1 repeater258/X sky130_fd_sc_hd__buf_8
X_17878_ _16109_/Y _16110_/Y _16111_/Y _16112_/Y _17908_/S0 _18759_/Q vssd1 vssd1
+ vccd1 vccd1 _17878_/X sky130_fd_sc_hd__mux4_2
Xrepeater269 repeater273/X vssd1 vssd1 vccd1 vccd1 repeater269/X sky130_fd_sc_hd__buf_8
XFILLER_65_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16603__A2 _16394_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19617_ _19937_/CLK _19617_/D repeater230/X vssd1 vssd1 vccd1 vccd1 _19617_/Q sky130_fd_sc_hd__dfrtp_1
X_16829_ _16828_/X _18833_/Q _17386_/S vssd1 vssd1 vccd1 vccd1 _16829_/X sky130_fd_sc_hd__mux2_2
XFILLER_81_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19548_ _19582_/CLK _19548_/D hold346/A vssd1 vssd1 vccd1 vccd1 _19548_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12625__B1 _12392_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09301_ _18658_/Q _09329_/A vssd1 vssd1 vccd1 vccd1 _09302_/A sky130_fd_sc_hd__nand2_1
XFILLER_206_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19479_ _19506_/CLK hold182/X repeater256/X vssd1 vssd1 vccd1 vccd1 _19479_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_22_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11731__A _11731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09232_ _09229_/Y _15710_/A _19882_/Q _09231_/A vssd1 vssd1 vccd1 vccd1 _09232_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_221_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09163_ _09164_/A vssd1 vssd1 vccd1 vccd1 _09163_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_119_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09094_ _12232_/A vssd1 vssd1 vccd1 vccd1 _09094_/X sky130_fd_sc_hd__buf_4
XFILLER_119_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18970__RESET_B hold348/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11178__A _11192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17564__S _17564_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09996_ _19944_/Q _09995_/Y _09854_/B _09964_/X vssd1 vssd1 vccd1 vccd1 _19944_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_88_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08947_ _18781_/Q vssd1 vssd1 vccd1 vccd1 _08947_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19946__CLK _19976_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16908__S _17541_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10840_ _10715_/X _19717_/Q _10840_/S vssd1 vssd1 vccd1 vccd1 _19717_/D sky130_fd_sc_hd__mux2_1
XFILLER_71_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_232_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10771_ _10771_/A _10771_/B vssd1 vssd1 vccd1 vccd1 _10773_/A sky130_fd_sc_hd__or2_2
XFILLER_52_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12510_ _19079_/Q _12505_/X _12408_/X _12506_/X vssd1 vssd1 vccd1 vccd1 _19079_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_44_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_240_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13490_ _13483_/A _13483_/B _18837_/Q _13432_/X _13426_/X vssd1 vssd1 vccd1 vccd1
+ _18837_/D sky130_fd_sc_hd__o221a_1
XFILLER_185_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19005__RESET_B hold346/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_233_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12441_ _12457_/A vssd1 vssd1 vccd1 vccd1 _12441_/X sky130_fd_sc_hd__buf_1
XFILLER_8_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17739__S _18508_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10257__A _14300_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12372_ _12372_/A _12659_/B vssd1 vssd1 vccd1 vccd1 _12427_/A sky130_fd_sc_hd__or2_2
X_15160_ _15160_/A vssd1 vssd1 vccd1 vccd1 _15160_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_181_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15767__B _18514_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11323_ _11488_/A _18990_/Q _19608_/Q _11320_/Y _11322_/X vssd1 vssd1 vccd1 vccd1
+ _11331_/B sky130_fd_sc_hd__o221a_1
X_14111_ _14111_/A vssd1 vssd1 vccd1 vccd1 _14111_/Y sky130_fd_sc_hd__clkinv_1
X_15091_ _17996_/Q _15084_/A hold263/X _15085_/A vssd1 vssd1 vccd1 vccd1 _17996_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_176_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14042_ _19088_/Q vssd1 vssd1 vccd1 vccd1 _14042_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14541__B1 _14513_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11254_ _19590_/Q _19004_/Q _11470_/A _11253_/Y vssd1 vssd1 vccd1 vccd1 _11261_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10704__B _10704_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17474__S _17474_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10205_ _19831_/Q _19658_/Q _10203_/Y _10958_/A vssd1 vssd1 vccd1 vccd1 _10209_/C
+ sky130_fd_sc_hd__o22a_1
X_18850_ _18866_/CLK _18850_/D repeater232/X vssd1 vssd1 vccd1 vccd1 _18850_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_192_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11185_ _11192_/A vssd1 vssd1 vccd1 vccd1 _11185_/X sky130_fd_sc_hd__clkbuf_2
X_17801_ _18186_/Q _18178_/Q _18170_/Q _18154_/Q _17918_/S0 _18750_/Q vssd1 vssd1
+ vccd1 vccd1 _17801_/X sky130_fd_sc_hd__mux4_2
X_10136_ _10136_/A vssd1 vssd1 vccd1 vccd1 _10136_/X sky130_fd_sc_hd__clkbuf_2
X_18781_ _19865_/CLK _18781_/D repeater265/X vssd1 vssd1 vccd1 vccd1 _18781_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_48_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15993_ _16634_/A vssd1 vssd1 vccd1 vccd1 _16512_/A sky130_fd_sc_hd__buf_2
XFILLER_248_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17732_ _15377_/X _19713_/Q _18508_/D vssd1 vssd1 vccd1 vccd1 _17732_/X sky130_fd_sc_hd__mux2_1
X_10067_ _10042_/A _10042_/B _10032_/A _10065_/Y vssd1 vssd1 vccd1 vccd1 _19926_/D
+ sky130_fd_sc_hd__a211oi_2
X_14944_ _18087_/Q _14939_/X _14927_/X _14941_/X vssd1 vssd1 vccd1 vccd1 _18087_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_248_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19846__RESET_B repeater270/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17663_ _15582_/Y _19026_/Q _17664_/S vssd1 vssd1 vccd1 vccd1 _18589_/D sky130_fd_sc_hd__mux2_1
X_14875_ _18128_/Q _14871_/X _14703_/X _14873_/X vssd1 vssd1 vccd1 vccd1 _18128_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16818__S _17536_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_235_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19402_ _19984_/CLK _19402_/D repeater244/X vssd1 vssd1 vccd1 vccd1 _19402_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_211_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16614_ _16572_/X _16614_/B _16614_/C vssd1 vssd1 vccd1 vccd1 _16614_/Y sky130_fd_sc_hd__nand3b_4
XFILLER_90_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12607__B1 _12541_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13826_ _13912_/C _13924_/A vssd1 vssd1 vccd1 vccd1 _13827_/B sky130_fd_sc_hd__or2_2
X_17594_ _15348_/X _19709_/Q _17600_/S vssd1 vssd1 vccd1 vccd1 _17594_/X sky130_fd_sc_hd__mux2_1
XFILLER_35_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19333_ _20013_/CLK _19333_/D repeater243/X vssd1 vssd1 vccd1 vccd1 _19333_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_232_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16545_ _16616_/A vssd1 vssd1 vccd1 vccd1 _16583_/B sky130_fd_sc_hd__buf_6
X_13757_ _13757_/A vssd1 vssd1 vccd1 vccd1 _13757_/Y sky130_fd_sc_hd__inv_2
X_10969_ _12053_/B vssd1 vssd1 vccd1 vccd1 _17614_/S sky130_fd_sc_hd__buf_4
XFILLER_203_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12708_ _15222_/A _12708_/B _12708_/C vssd1 vssd1 vccd1 vccd1 _12710_/A sky130_fd_sc_hd__or3_4
X_19264_ _19952_/CLK _19264_/D repeater245/X vssd1 vssd1 vccd1 vccd1 _19264_/Q sky130_fd_sc_hd__dfrtp_1
X_16476_ _09308_/Y _15915_/X _09217_/Y _15884_/X vssd1 vssd1 vccd1 vccd1 _16476_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_203_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13688_ _18770_/Q _13685_/X _13676_/X _13686_/Y vssd1 vssd1 vccd1 vccd1 _18770_/D
+ sky130_fd_sc_hd__a22o_1
X_18215_ _19849_/CLK _18215_/D vssd1 vssd1 vccd1 vccd1 _18215_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09021__A hold291/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15427_ _19618_/Q _11163_/B _11164_/B vssd1 vssd1 vccd1 vccd1 _15427_/X sky130_fd_sc_hd__a21bo_1
XFILLER_176_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17649__S _17655_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12639_ _19007_/Q _12636_/X hold233/X _12637_/X vssd1 vssd1 vccd1 vccd1 _19007_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19195_ _19222_/CLK _19195_/D repeater188/X vssd1 vssd1 vccd1 vccd1 _19195_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18799__RESET_B repeater258/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18146_ _19851_/CLK _18146_/D vssd1 vssd1 vccd1 vccd1 _18146_/Q sky130_fd_sc_hd__dfxtp_1
X_15358_ _15358_/A _17590_/X vssd1 vssd1 vccd1 vccd1 _18500_/D sky130_fd_sc_hd__and2_1
XFILLER_184_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18728__RESET_B repeater253/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14309_ _18446_/Q _14303_/X _13674_/X _14305_/X vssd1 vssd1 vccd1 vccd1 _18446_/D
+ sky130_fd_sc_hd__a22o_1
Xhold205 hold205/A vssd1 vssd1 vccd1 vccd1 hold205/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18077_ _18137_/CLK _18077_/D vssd1 vssd1 vccd1 vccd1 _18077_/Q sky130_fd_sc_hd__dfxtp_1
X_15289_ _15289_/A _15289_/B vssd1 vssd1 vccd1 vccd1 _15290_/A sky130_fd_sc_hd__or2_1
XANTENNA__12382__A hold289/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold216 hold216/A vssd1 vssd1 vccd1 vccd1 hold216/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold227 hold227/A vssd1 vssd1 vccd1 vccd1 hold227/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16521__B2 _16235_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold238 HWDATA[6] vssd1 vssd1 vccd1 vccd1 input66/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold249 HWDATA[7] vssd1 vssd1 vccd1 vccd1 input67/A sky130_fd_sc_hd__dlygate4sd3_1
X_17028_ _17027_/X _19947_/Q _17518_/S vssd1 vssd1 vccd1 vccd1 _17028_/X sky130_fd_sc_hd__mux2_2
XFILLER_113_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17384__S _17414_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09850_ _09850_/A _09850_/B vssd1 vssd1 vccd1 vccd1 _09998_/A sky130_fd_sc_hd__or2_1
XFILLER_113_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18843__CLK _18866_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09781_ _09781_/A vssd1 vssd1 vccd1 vccd1 _09781_/Y sky130_fd_sc_hd__inv_2
X_18979_ _19597_/CLK _18979_/D hold273/X vssd1 vssd1 vccd1 vccd1 _18979_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_105_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17880__S0 _17913_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_222_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17559__S _17564_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20074__RESET_B repeater196/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09215_ _18650_/Q _09214_/B _09214_/Y vssd1 vssd1 vccd1 vccd1 _15715_/A sky130_fd_sc_hd__o21ai_1
XFILLER_195_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09146_ _09146_/A vssd1 vssd1 vccd1 vccd1 _09146_/Y sky130_fd_sc_hd__inv_2
XFILLER_108_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09077_ hold268/X vssd1 vssd1 vccd1 vccd1 _09077_/X sky130_fd_sc_hd__buf_6
XFILLER_107_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17294__S _17543_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09979_ _19954_/Q _09978_/Y _09968_/X _09863_/B vssd1 vssd1 vccd1 vccd1 _19954_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__16211__B _16212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20099_ _20122_/CLK _20099_/D repeater234/X vssd1 vssd1 vccd1 vccd1 _20099_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_162_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12990_ _12965_/B _12879_/B _12988_/Y _12986_/X vssd1 vssd1 vccd1 vccd1 _18937_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_183_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11941_ _11979_/A vssd1 vssd1 vccd1 vccd1 _11956_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_91_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16579__A1 _17263_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16579__B2 _15887_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_217_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_232_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14660_ _18248_/Q _14656_/X _14604_/X _14658_/X vssd1 vssd1 vccd1 vccd1 _18248_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_205_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17871__S0 _17913_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11872_ _12371_/A _15888_/A vssd1 vssd1 vccd1 vccd1 _11998_/A sky130_fd_sc_hd__or2_4
XFILLER_214_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13611_ _18805_/Q _13610_/Y _13591_/A _13530_/B vssd1 vssd1 vccd1 vccd1 _18805_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_189_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10823_ _17750_/X vssd1 vssd1 vccd1 vccd1 _10823_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14591_ _18288_/Q _14587_/X _14535_/X _14589_/X vssd1 vssd1 vccd1 vccd1 _18288_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_60_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10076__B1 _10079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16330_ _18032_/Q vssd1 vssd1 vccd1 vccd1 _16330_/Y sky130_fd_sc_hd__inv_2
X_13542_ _13542_/A _13586_/A vssd1 vssd1 vccd1 vccd1 _13543_/B sky130_fd_sc_hd__or2_2
XFILLER_111_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10754_ _10754_/A vssd1 vssd1 vccd1 vccd1 _10754_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17469__S _17565_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16261_ _18015_/Q vssd1 vssd1 vccd1 vccd1 _16261_/Y sky130_fd_sc_hd__inv_2
X_13473_ _13473_/A vssd1 vssd1 vccd1 vccd1 _13473_/Y sky130_fd_sc_hd__inv_2
X_10685_ _19500_/Q _14245_/C vssd1 vssd1 vccd1 vccd1 _15829_/B sky130_fd_sc_hd__or2_1
XFILLER_71_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18000_ _18465_/CLK _18000_/D vssd1 vssd1 vccd1 vccd1 _18000_/Q sky130_fd_sc_hd__dfxtp_1
X_15212_ _19722_/Q _15209_/X _15216_/C _15211_/Y vssd1 vssd1 vccd1 vccd1 _15213_/B
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__12368__A2 _12334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_185_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12424_ _19135_/Q _12420_/X _12223_/X _12421_/X vssd1 vssd1 vccd1 vccd1 _19135_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14762__B1 _14745_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16192_ _18086_/Q vssd1 vssd1 vccd1 vccd1 _16192_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18821__RESET_B repeater231/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15143_ _17962_/Q _15135_/A _09339_/X _15136_/A vssd1 vssd1 vccd1 vccd1 _17962_/D
+ sky130_fd_sc_hd__a22o_1
X_12355_ _19169_/Q _12352_/X _12353_/X _12354_/X vssd1 vssd1 vccd1 vccd1 _19169_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10715__A _14793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18866__CLK _18866_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11306_ _19597_/Q _11305_/Y _11472_/A _18974_/Q vssd1 vssd1 vccd1 vccd1 _11306_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__14514__B1 _14513_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15074_ _18009_/Q _15071_/X hold247/X _15073_/X vssd1 vssd1 vccd1 vccd1 _18009_/D
+ sky130_fd_sc_hd__a22o_1
X_12286_ _19208_/Q _12283_/X _12026_/X _12284_/X vssd1 vssd1 vccd1 vccd1 _19208_/D
+ sky130_fd_sc_hd__a22o_1
X_19951_ _19952_/CLK _19951_/D repeater244/X vssd1 vssd1 vccd1 vccd1 _19951_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_153_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14025_ _14025_/A _14111_/A vssd1 vssd1 vccd1 vccd1 _14026_/B sky130_fd_sc_hd__or2_2
X_11237_ _19583_/Q vssd1 vssd1 vccd1 vccd1 _11464_/A sky130_fd_sc_hd__inv_2
X_18902_ _19956_/CLK _18902_/D repeater245/X vssd1 vssd1 vccd1 vccd1 _18902_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_206_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19882_ _20059_/CLK _19882_/D repeater199/X vssd1 vssd1 vccd1 vccd1 _19882_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12930__A _19266_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11168_ _19623_/Q _11168_/B vssd1 vssd1 vccd1 vccd1 _11169_/B sky130_fd_sc_hd__or2_1
X_18833_ _19255_/CLK _18833_/D repeater237/X vssd1 vssd1 vccd1 vccd1 _18833_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_67_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10119_ _18567_/Q _15486_/A vssd1 vssd1 vccd1 vccd1 _15490_/A sky130_fd_sc_hd__or2_2
X_18764_ _18765_/CLK _18764_/D repeater196/X vssd1 vssd1 vccd1 vccd1 _18764_/Q sky130_fd_sc_hd__dfrtp_4
X_15976_ _16055_/A vssd1 vssd1 vccd1 vccd1 _15976_/X sky130_fd_sc_hd__clkbuf_2
X_11099_ _11061_/X _11098_/X _11061_/X _11098_/X vssd1 vssd1 vccd1 vccd1 _11103_/C
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_222_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17715_ _15425_/X _19526_/Q _18546_/D vssd1 vssd1 vccd1 vccd1 _17715_/X sky130_fd_sc_hd__mux2_1
XFILLER_76_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09016__A hold284/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14927_ _20079_/Q vssd1 vssd1 vccd1 vccd1 _14927_/X sky130_fd_sc_hd__clkbuf_2
X_18695_ _19119_/CLK _18695_/D hold351/X vssd1 vssd1 vccd1 vccd1 _18695_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_64_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18246__CLK _19847_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17646_ _15652_/X _19043_/Q _17655_/S vssd1 vssd1 vccd1 vccd1 _18606_/D sky130_fd_sc_hd__mux2_1
XFILLER_91_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17862__S0 _17913_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14858_ _14859_/A vssd1 vssd1 vccd1 vccd1 _14858_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_212_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13809_ _18712_/Q vssd1 vssd1 vccd1 vccd1 _13949_/A sky130_fd_sc_hd__inv_2
XANTENNA__13253__A0 _12313_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17577_ _15406_/X _19766_/Q _17584_/S vssd1 vssd1 vccd1 vccd1 _17577_/X sky130_fd_sc_hd__mux2_1
X_14789_ _18176_/Q _14785_/X _14749_/X _14787_/X vssd1 vssd1 vccd1 vccd1 _18176_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_211_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19316_ _19324_/CLK _19316_/D repeater213/X vssd1 vssd1 vccd1 vccd1 _19316_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__11281__A _19012_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16528_ _17199_/X _15904_/X _17190_/X _16509_/X vssd1 vssd1 vccd1 vccd1 _16528_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_220_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18909__RESET_B repeater188/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19247_ _19320_/CLK _19247_/D repeater214/X vssd1 vssd1 vccd1 vccd1 _19247_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__17379__S _17474_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16459_ _17314_/X _15900_/A _17083_/X _16234_/A vssd1 vssd1 vccd1 vccd1 _16459_/X
+ sky130_fd_sc_hd__o22a_2
XANTENNA__16742__B2 _16235_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09000_ _19498_/Q vssd1 vssd1 vccd1 vccd1 _15749_/A sky130_fd_sc_hd__buf_1
X_19178_ _19288_/CLK _19178_/D repeater212/X vssd1 vssd1 vccd1 vccd1 _19178_/Q sky130_fd_sc_hd__dfrtp_4
X_18129_ _20090_/CLK _18129_/D vssd1 vssd1 vccd1 vccd1 _18129_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17917__S1 _18750_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13001__A _13021_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09902_ _09873_/A _19357_/Q _19950_/Q _09901_/Y vssd1 vssd1 vccd1 vccd1 _09902_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_99_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20022_ _20091_/CLK _20022_/D repeater238/X vssd1 vssd1 vccd1 vccd1 _20022_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__13655__B _15169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09833_ _19953_/Q vssd1 vssd1 vccd1 vccd1 _09861_/A sky130_fd_sc_hd__inv_2
X_09764_ _19998_/Q _09758_/C _09763_/X _09761_/A vssd1 vssd1 vccd1 vccd1 _19998_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_55_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11175__B _18546_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_2_0_0_HCLK_A clkbuf_2_1_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09695_ _20001_/Q _19430_/Q _20001_/Q _19430_/Q vssd1 vssd1 vccd1 vccd1 _09695_/X
+ sky130_fd_sc_hd__a2bb2o_1
Xrebuffer20 _13070_/B vssd1 vssd1 vccd1 vccd1 _13196_/A sky130_fd_sc_hd__dlygate4sd1_1
XPHY_4017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer31 _13069_/C vssd1 vssd1 vccd1 vccd1 _13198_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_4028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrebuffer42 _11468_/C vssd1 vssd1 vccd1 vccd1 _11529_/A sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_242_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer53 _11467_/B vssd1 vssd1 vccd1 vccd1 _11533_/C1 sky130_fd_sc_hd__dlygate4sd1_1
XANTENNA__17853__S0 _17913_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrebuffer64 _13064_/B vssd1 vssd1 vccd1 vccd1 _13211_/C1 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrebuffer75 _13073_/B vssd1 vssd1 vccd1 vccd1 _13192_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_242_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrebuffer86 _14028_/B vssd1 vssd1 vccd1 vccd1 _14109_/C1 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrebuffer97 _14026_/B vssd1 vssd1 vccd1 vccd1 _14113_/B1 sky130_fd_sc_hd__dlygate4sd1_1
XANTENNA__18739__CLK _20051_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13244__B1 _12596_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11191__A _11191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17289__S _17413_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16733__B2 _16002_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer110 _14020_/B vssd1 vssd1 vccd1 vccd1 _14122_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_109_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10470_ _18548_/Q _10470_/B vssd1 vssd1 vccd1 vccd1 _19823_/D sky130_fd_sc_hd__or2_1
Xrebuffer121 _09857_/C vssd1 vssd1 vccd1 vccd1 _09988_/A sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_6_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17908__S1 _18759_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09129_ _09133_/C _09136_/B vssd1 vssd1 vccd1 vccd1 _09129_/Y sky130_fd_sc_hd__nor2_1
XFILLER_108_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16921__S _17318_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16497__B1 _17227_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12140_ _19291_/Q _12134_/X _12076_/X _12137_/X vssd1 vssd1 vccd1 vccd1 _19291_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_2_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12071_ _12122_/A vssd1 vssd1 vccd1 vccd1 _12096_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_89_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11022_ _11029_/A vssd1 vssd1 vccd1 vccd1 _11022_/X sky130_fd_sc_hd__buf_1
XFILLER_89_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19438__RESET_B repeater210/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15830_ _15830_/A vssd1 vssd1 vccd1 vccd1 _15831_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__11366__A _19129_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15761_ _15765_/C _18526_/D _18527_/Q vssd1 vssd1 vccd1 vccd1 _18522_/D sky130_fd_sc_hd__and3_1
XANTENNA__17749__A0 _15753_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12973_ _18946_/Q _12972_/Y _12888_/B _12972_/A _12958_/X vssd1 vssd1 vccd1 vccd1
+ _18946_/D sky130_fd_sc_hd__o221a_1
X_17500_ _17499_/X _15956_/Y _17565_/S vssd1 vssd1 vccd1 vccd1 _17500_/X sky130_fd_sc_hd__mux2_1
X_14712_ _18220_/Q _14700_/A _14711_/X _14701_/A vssd1 vssd1 vccd1 vccd1 _18220_/D
+ sky130_fd_sc_hd__a22o_1
X_18480_ _20049_/CLK _18480_/D repeater202/X vssd1 vssd1 vccd1 vccd1 _18480_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17844__S0 _19633_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11924_ _12238_/A vssd1 vssd1 vccd1 vccd1 _11924_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_206_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15692_ _18616_/Q vssd1 vssd1 vccd1 vccd1 _15692_/Y sky130_fd_sc_hd__inv_2
XPHY_4540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17431_ _17430_/X _08952_/Y _17566_/S vssd1 vssd1 vccd1 vccd1 _17431_/X sky130_fd_sc_hd__mux2_1
XPHY_4562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14643_ _14644_/A vssd1 vssd1 vccd1 vccd1 _14643_/X sky130_fd_sc_hd__clkbuf_2
XPHY_4573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11855_ _11855_/A vssd1 vssd1 vccd1 vccd1 _15201_/B sky130_fd_sc_hd__clkbuf_2
XPHY_4584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output105_A _16251_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17362_ _17361_/X _13065_/A _17488_/S vssd1 vssd1 vccd1 vccd1 _17362_/X sky130_fd_sc_hd__mux2_1
X_10806_ _10806_/A vssd1 vssd1 vccd1 vccd1 _17621_/S sky130_fd_sc_hd__clkbuf_4
XPHY_3872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14574_ _14574_/A vssd1 vssd1 vccd1 vccd1 _14574_/X sky130_fd_sc_hd__clkbuf_2
XPHY_3883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11786_ _11822_/A vssd1 vssd1 vccd1 vccd1 _11801_/A sky130_fd_sc_hd__buf_2
XFILLER_220_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19101_ _19585_/CLK _19101_/D hold365/X vssd1 vssd1 vccd1 vccd1 _19101_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__11797__B1 hold305/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_186_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16313_ _16312_/Y _16303_/X _15751_/Y _15850_/B vssd1 vssd1 vccd1 vccd1 _16313_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__17199__S _17548_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13525_ _18761_/Q _13524_/X _18761_/Q _13524_/X vssd1 vssd1 vccd1 vccd1 _13525_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_10737_ _10519_/D _10733_/Y _11653_/B _11650_/B _10736_/X vssd1 vssd1 vccd1 vccd1
+ _15271_/D sky130_fd_sc_hd__a2111o_1
XFILLER_159_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17293_ _16484_/X _08924_/Y _17566_/S vssd1 vssd1 vccd1 vccd1 _17293_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19032_ _19577_/CLK _19032_/D repeater269/X vssd1 vssd1 vccd1 vccd1 _19032_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__14735__B1 _14600_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16244_ _16530_/A vssd1 vssd1 vccd1 vccd1 _16597_/A sky130_fd_sc_hd__clkinv_4
X_13456_ _13456_/A vssd1 vssd1 vccd1 vccd1 _13456_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10668_ _17733_/X _10661_/X _19792_/Q _10663_/X vssd1 vssd1 vccd1 vccd1 _19792_/D
+ sky130_fd_sc_hd__a22o_1
X_12407_ _19145_/Q _12400_/X _12406_/X _12402_/X vssd1 vssd1 vccd1 vccd1 _19145_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_154_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16175_ _18230_/Q vssd1 vssd1 vccd1 vccd1 _16175_/Y sky130_fd_sc_hd__inv_2
X_10599_ _18482_/Q vssd1 vssd1 vccd1 vccd1 _15224_/A sky130_fd_sc_hd__clkbuf_2
X_13387_ _18865_/Q vssd1 vssd1 vccd1 vccd1 _13387_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16831__S _17488_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_217_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput107 _16397_/Y vssd1 vssd1 vccd1 vccd1 HRDATA[6] sky130_fd_sc_hd__clkbuf_2
Xoutput118 _16758_/LO vssd1 vssd1 vccd1 vccd1 IRQ[15] sky130_fd_sc_hd__clkbuf_2
X_15126_ _17975_/Q _15122_/X _14925_/X _15124_/X vssd1 vssd1 vccd1 vccd1 _17975_/D
+ sky130_fd_sc_hd__a22o_1
Xoutput129 _19732_/Q vssd1 vssd1 vccd1 vccd1 MSO_S3 sky130_fd_sc_hd__clkbuf_2
XFILLER_142_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12338_ _19177_/Q _12334_/X _12100_/X _12335_/X vssd1 vssd1 vccd1 vccd1 _19177_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_99_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19934_ _19937_/CLK _19934_/D repeater189/X vssd1 vssd1 vccd1 vccd1 _19934_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_142_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15057_ _18018_/Q _15048_/A _15020_/X _15049_/A vssd1 vssd1 vccd1 vccd1 _18018_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12660__A _12698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12269_ _12276_/A vssd1 vssd1 vccd1 vccd1 _12269_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_96_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14008_ _14008_/A _14142_/A vssd1 vssd1 vccd1 vccd1 _14009_/B sky130_fd_sc_hd__or2_1
X_19865_ _19865_/CLK _19865_/D repeater262/X vssd1 vssd1 vccd1 vccd1 _19865_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__19179__RESET_B repeater212/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18816_ _18856_/CLK _18816_/D repeater217/X vssd1 vssd1 vccd1 vccd1 _18816_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_233_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19796_ _19810_/CLK _19796_/D repeater226/X vssd1 vssd1 vccd1 vccd1 _19796_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_56_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14266__A2 _14259_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18747_ _20059_/CLK _18747_/D repeater198/X vssd1 vssd1 vccd1 vccd1 _18747_/Q sky130_fd_sc_hd__dfrtp_4
X_15959_ _15961_/A vssd1 vssd1 vccd1 vccd1 _16204_/A sky130_fd_sc_hd__buf_1
XFILLER_48_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09480_ _09480_/A _09480_/B vssd1 vssd1 vccd1 vccd1 _09592_/A sky130_fd_sc_hd__or2_1
XANTENNA__17835__S0 _17908_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18678_ _18686_/CLK _18678_/D repeater252/X vssd1 vssd1 vccd1 vccd1 _18678_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_224_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17629_ _19890_/Q _19743_/Q _17630_/S vssd1 vssd1 vccd1 vccd1 _17629_/X sky130_fd_sc_hd__mux2_1
XFILLER_51_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_196_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11788__B1 _09016_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_192_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19949__RESET_B hold371/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11960__B1 _09049_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_207_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19531__RESET_B repeater221/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17572__S _17584_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20005_ _20091_/CLK _20005_/D repeater236/X vssd1 vssd1 vccd1 vccd1 _20005_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_59_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09816_ _19971_/Q _09607_/X _09815_/Y vssd1 vssd1 vccd1 vccd1 _19971_/D sky130_fd_sc_hd__o21a_1
XFILLER_143_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_4_5_0_HCLK clkbuf_4_5_0_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_opt_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_100_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09747_ _09747_/A _09775_/A vssd1 vssd1 vccd1 vccd1 _09748_/B sky130_fd_sc_hd__or2_2
XFILLER_246_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18561__CLK _19992_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17826__S0 _17918_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09678_ _20003_/Q _09677_/Y _09670_/Y _19432_/Q vssd1 vssd1 vccd1 vccd1 _09678_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA_hold348_A hold348/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16916__S _17474_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11640_ _11548_/B _11642_/A _11548_/A vssd1 vssd1 vccd1 vccd1 _11641_/B sky130_fd_sc_hd__o21a_1
XPHY_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11571_ _11571_/A _11571_/B vssd1 vssd1 vccd1 vccd1 _11615_/A sky130_fd_sc_hd__or2_1
XFILLER_52_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13310_ _18855_/Q vssd1 vssd1 vccd1 vccd1 _13429_/A sky130_fd_sc_hd__inv_6
XPHY_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10522_ _11655_/A _10522_/B _19529_/Q _10734_/C vssd1 vssd1 vccd1 vccd1 _10735_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_168_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14290_ _14290_/A vssd1 vssd1 vccd1 vccd1 _14290_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13241_ _13242_/A vssd1 vssd1 vccd1 vccd1 _13241_/X sky130_fd_sc_hd__clkbuf_2
X_10453_ _19831_/Q _10450_/X _10451_/X _10452_/X vssd1 vssd1 vccd1 vccd1 _19831_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_182_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10384_ _10345_/X _10321_/C _10368_/X _10383_/X vssd1 vssd1 vccd1 vccd1 _19854_/D
+ sky130_fd_sc_hd__o22ai_1
X_13172_ _13172_/A vssd1 vssd1 vccd1 vccd1 _13172_/Y sky130_fd_sc_hd__inv_2
XFILLER_184_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19619__RESET_B repeater230/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11951__B1 _09033_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12123_ _19300_/Q _12121_/X _11978_/X _12122_/X vssd1 vssd1 vccd1 vccd1 _19300_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_184_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17980_ _20124_/CLK _17980_/D vssd1 vssd1 vccd1 vccd1 _17980_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12054_ _17614_/S _12052_/X _11853_/A _12053_/Y vssd1 vssd1 vccd1 vccd1 _12055_/B
+ sky130_fd_sc_hd__o22a_1
X_16931_ _19475_/Q hold196/X _16950_/S vssd1 vssd1 vccd1 vccd1 _16931_/X sky130_fd_sc_hd__mux2_4
XFILLER_96_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17482__S _17482_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11005_ _11005_/A vssd1 vssd1 vccd1 vccd1 _11006_/B sky130_fd_sc_hd__inv_2
XFILLER_77_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_238_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19650_ _19859_/CLK _19650_/D repeater262/X vssd1 vssd1 vccd1 vccd1 _19650_/Q sky130_fd_sc_hd__dfrtp_1
X_16862_ _17473_/A0 _16602_/Y _17547_/S vssd1 vssd1 vccd1 vccd1 _16862_/X sky130_fd_sc_hd__mux2_1
XFILLER_238_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18601_ _19867_/CLK _18601_/D repeater263/X vssd1 vssd1 vccd1 vccd1 _18601_/Q sky130_fd_sc_hd__dfrtp_1
X_15813_ _17977_/Q vssd1 vssd1 vccd1 vccd1 _15813_/Y sky130_fd_sc_hd__inv_2
X_19581_ _19591_/CLK _19581_/D hold363/X vssd1 vssd1 vccd1 vccd1 _19581_/Q sky130_fd_sc_hd__dfrtp_1
X_16793_ _16792_/X _13894_/Y _17545_/S vssd1 vssd1 vccd1 vccd1 _16793_/X sky130_fd_sc_hd__mux2_1
XFILLER_225_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_203_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15996__A2 _16512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18532_ _19937_/CLK _18532_/D repeater189/X vssd1 vssd1 vccd1 vccd1 _18532_/Q sky130_fd_sc_hd__dfrtp_1
X_15744_ _15747_/C _15744_/B _18489_/Q vssd1 vssd1 vccd1 vccd1 _18485_/D sky130_fd_sc_hd__nor3_1
XANTENNA__20106__RESET_B repeater230/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17817__S0 _17918_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12956_ _12956_/A _12956_/B _12956_/C _12956_/D vssd1 vssd1 vccd1 vccd1 _12968_/B
+ sky130_fd_sc_hd__and4_2
XFILLER_33_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_234_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18463_ _18465_/CLK _18463_/D vssd1 vssd1 vccd1 vccd1 _18463_/Q sky130_fd_sc_hd__dfxtp_1
X_11907_ _19412_/Q _11905_/X _09071_/X _11906_/X vssd1 vssd1 vccd1 vccd1 _19412_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_33_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15675_ _18612_/Q vssd1 vssd1 vccd1 vccd1 _15675_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16826__S _17523_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12887_ _12887_/A _12975_/A _12887_/C vssd1 vssd1 vccd1 vccd1 _12972_/A sky130_fd_sc_hd__or3_4
XFILLER_221_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17414_ _17413_/X _09468_/A _17414_/S vssd1 vssd1 vccd1 vccd1 _17414_/X sky130_fd_sc_hd__mux2_1
XPHY_4392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14626_ _20074_/Q vssd1 vssd1 vccd1 vccd1 _14626_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__09013__B _12659_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18394_ _18412_/CLK _18394_/D vssd1 vssd1 vccd1 vccd1 _18394_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11838_ _12183_/B vssd1 vssd1 vccd1 vccd1 _15776_/A sky130_fd_sc_hd__clkbuf_4
XPHY_3680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17345_ _16345_/X _19832_/Q _17566_/S vssd1 vssd1 vccd1 vccd1 _17345_/X sky130_fd_sc_hd__mux2_1
XFILLER_186_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14557_ _14598_/A _19643_/Q _14557_/C vssd1 vssd1 vccd1 vccd1 _14559_/A sky130_fd_sc_hd__or3_4
XANTENNA__12431__A1 _19130_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11769_ hold190/X _11764_/X _19477_/Q _11765_/X vssd1 vssd1 vccd1 vccd1 hold192/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_202_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13508_ _14695_/A _14696_/B vssd1 vssd1 vccd1 vccd1 _13523_/A sky130_fd_sc_hd__or2_2
Xclkbuf_opt_4_HCLK clkbuf_opt_4_HCLK/A vssd1 vssd1 vccd1 vccd1 _18545_/CLK sky130_fd_sc_hd__clkbuf_16
X_17276_ _16484_/X _10219_/Y _17566_/S vssd1 vssd1 vccd1 vccd1 _17276_/X sky130_fd_sc_hd__mux2_1
X_14488_ _18346_/Q _14479_/A _14268_/X _14480_/A vssd1 vssd1 vccd1 vccd1 _18346_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_133_HCLK_A clkbuf_4_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19015_ _19115_/CLK _19015_/D hold353/X vssd1 vssd1 vccd1 vccd1 _19015_/Q sky130_fd_sc_hd__dfrtp_4
X_16227_ _18876_/Q vssd1 vssd1 vccd1 vccd1 _16227_/Y sky130_fd_sc_hd__inv_2
X_13439_ _13439_/A vssd1 vssd1 vccd1 vccd1 _13439_/Y sky130_fd_sc_hd__inv_2
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12195__B1 _12076_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16158_ _18038_/Q vssd1 vssd1 vccd1 vccd1 _16158_/Y sky130_fd_sc_hd__inv_2
XFILLER_154_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15109_ _15109_/A _15109_/B _15121_/C vssd1 vssd1 vccd1 vccd1 _15111_/A sky130_fd_sc_hd__or3_4
XFILLER_114_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12390__A _12402_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16089_ _18349_/Q vssd1 vssd1 vccd1 vccd1 _16089_/Y sky130_fd_sc_hd__inv_2
X_08980_ _08982_/B vssd1 vssd1 vccd1 vccd1 _08980_/Y sky130_fd_sc_hd__inv_2
XFILLER_170_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19917_ _19937_/CLK _19917_/D repeater190/X vssd1 vssd1 vccd1 vccd1 _19917_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17392__S _17548_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19848_ _19849_/CLK _19848_/D repeater257/X vssd1 vssd1 vccd1 vccd1 _19848_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_84_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09601_ _09601_/A vssd1 vssd1 vccd1 vccd1 _09604_/A sky130_fd_sc_hd__inv_2
XFILLER_228_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19779_ _19780_/CLK _19779_/D repeater218/X vssd1 vssd1 vccd1 vccd1 _19779_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_113_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09532_ _09479_/A _19309_/Q _20019_/Q _09531_/Y vssd1 vssd1 vccd1 vccd1 _09532_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_71_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17808__S0 _17918_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18924__RESET_B repeater212/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09463_ _09463_/A _09463_/B _09463_/C _09463_/D vssd1 vssd1 vccd1 vccd1 _09464_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_224_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09394_ _09379_/X _09385_/X _09394_/C _09394_/D vssd1 vssd1 vccd1 vccd1 _09394_/Y
+ sky130_fd_sc_hd__nand4bb_2
Xclkbuf_4_13_0_HCLK clkbuf_3_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_13_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_12_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_196_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_220_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17361__A1 _12945_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14175__A1 _19123_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17567__S _17567_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14175__B2 _18673_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14780__A _14780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19783__RESET_B repeater203/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_55_HCLK_A clkbuf_opt_3_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11909__A hold268/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_235_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12810_ _19230_/Q vssd1 vssd1 vccd1 vccd1 _12810_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13790_ _18722_/Q vssd1 vssd1 vccd1 vccd1 _13910_/A sky130_fd_sc_hd__inv_2
XANTENNA__12110__B1 _12026_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_216_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18307__CLK _19847_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12741_ _19250_/Q vssd1 vssd1 vccd1 vccd1 _12741_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_1_0_0_HCLK clkbuf_0_HCLK/X vssd1 vssd1 vccd1 vccd1 clkbuf_1_0_1_HCLK/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__16927__A1 hold193/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_231_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15460_ _15463_/B _15458_/X _15459_/X vssd1 vssd1 vccd1 vccd1 _15460_/X sky130_fd_sc_hd__o21a_1
XFILLER_231_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12672_ _18986_/Q _12670_/X hold303/X _12671_/X vssd1 vssd1 vccd1 vccd1 _18986_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14402__A2 _14395_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14411_ _14411_/A vssd1 vssd1 vccd1 vccd1 _14411_/X sky130_fd_sc_hd__clkbuf_2
XPHY_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11623_ _11623_/A _11632_/A vssd1 vssd1 vccd1 vccd1 _11624_/B sky130_fd_sc_hd__or2_1
XPHY_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15391_ _15391_/A _17584_/X vssd1 vssd1 vccd1 vccd1 _18528_/D sky130_fd_sc_hd__nor2_1
XPHY_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09814__C1 _09759_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17130_ _16543_/Y _19075_/Q _17490_/S vssd1 vssd1 vccd1 vccd1 _17130_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10424__B1 _10423_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13277__A1_N _18750_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14342_ _18430_/Q _14336_/X hold324/X _14338_/X vssd1 vssd1 vccd1 vccd1 _18430_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11554_ _11580_/A _11579_/A _11572_/A _11571_/A vssd1 vssd1 vccd1 vccd1 _11556_/C
+ sky130_fd_sc_hd__or4_4
XPHY_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09290__B1 _09082_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10505_ _10528_/C _19537_/Q _10505_/C vssd1 vssd1 vccd1 vccd1 _10736_/A sky130_fd_sc_hd__nor3_4
X_17061_ _15768_/Y _11258_/Y _17546_/S vssd1 vssd1 vccd1 vccd1 _17061_/X sky130_fd_sc_hd__mux2_1
XANTENNA__17477__S _17543_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15363__B1 _17600_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14273_ _14273_/A vssd1 vssd1 vccd1 vccd1 _14273_/X sky130_fd_sc_hd__buf_2
X_11485_ _11485_/A _11497_/A vssd1 vssd1 vccd1 vccd1 _11486_/B sky130_fd_sc_hd__or2_2
XFILLER_109_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12177__B1 _11922_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16012_ _18068_/Q vssd1 vssd1 vccd1 vccd1 _16012_/Y sky130_fd_sc_hd__inv_2
X_13224_ _18537_/Q _13224_/B vssd1 vssd1 vccd1 vccd1 _13225_/B sky130_fd_sc_hd__or2_1
XFILLER_109_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17104__A1 _19069_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10436_ _19841_/Q _10433_/X _09058_/X _10435_/X vssd1 vssd1 vccd1 vccd1 _19841_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_3_3_0_HCLK_A clkbuf_3_3_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19453__RESET_B repeater272/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13155_ _13152_/Y _18893_/Q _13153_/Y _18903_/Q _13154_/X vssd1 vssd1 vccd1 vccd1
+ _13159_/C sky130_fd_sc_hd__o221a_1
X_10367_ _19858_/Q _10367_/B vssd1 vssd1 vccd1 vccd1 _10367_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_repeater218_A repeater219/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12106_ _12121_/A vssd1 vssd1 vccd1 vccd1 _12106_/X sky130_fd_sc_hd__clkbuf_2
X_10298_ _18593_/Q _15593_/A vssd1 vssd1 vccd1 vccd1 _15597_/A sky130_fd_sc_hd__or2_1
X_13086_ _13086_/A _13169_/A vssd1 vssd1 vccd1 vccd1 _13087_/B sky130_fd_sc_hd__or2_2
X_17963_ _20036_/CLK _17963_/D vssd1 vssd1 vccd1 vccd1 _17963_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13677__B1 _13676_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19702_ _20055_/CLK _19702_/D repeater202/X vssd1 vssd1 vccd1 vccd1 _19702_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_214_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16914_ _16913_/X _18826_/Q _17386_/S vssd1 vssd1 vccd1 vccd1 _16914_/X sky130_fd_sc_hd__mux2_2
XFILLER_66_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12037_ _19342_/Q _12034_/X _12035_/X _12036_/X vssd1 vssd1 vccd1 vccd1 _19342_/D
+ sky130_fd_sc_hd__a22o_1
X_17894_ _17890_/X _17891_/X _17892_/X _17893_/X _19633_/Q _19634_/Q vssd1 vssd1 vccd1
+ vccd1 _17894_/X sky130_fd_sc_hd__mux4_2
XFILLER_66_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19633_ _19851_/CLK _19633_/D repeater258/X vssd1 vssd1 vccd1 vccd1 _19633_/Q sky130_fd_sc_hd__dfrtp_2
X_16845_ _17486_/A0 _13119_/Y _17543_/S vssd1 vssd1 vccd1 vccd1 _16845_/X sky130_fd_sc_hd__mux2_1
XFILLER_225_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16776_ _16775_/X _09391_/Y _17413_/S vssd1 vssd1 vccd1 vccd1 _16776_/X sky130_fd_sc_hd__mux2_1
X_19564_ _19576_/CLK _19564_/D repeater268/X vssd1 vssd1 vccd1 vccd1 _19564_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_230_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13988_ _18686_/Q vssd1 vssd1 vccd1 vccd1 _14016_/A sky130_fd_sc_hd__inv_4
XANTENNA__12101__B1 _12100_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18515_ _19822_/CLK _18515_/D repeater227/X vssd1 vssd1 vccd1 vccd1 _18515_/Q sky130_fd_sc_hd__dfrtp_1
X_15727_ _15727_/A _15727_/B vssd1 vssd1 vccd1 vccd1 _18660_/D sky130_fd_sc_hd__nor2_1
X_12939_ _12938_/Y _12891_/A _19292_/Q _18949_/Q vssd1 vssd1 vccd1 vccd1 _12939_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16918__A1 _09431_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19495_ _19515_/CLK hold262/X repeater260/X vssd1 vssd1 vccd1 vccd1 _19495_/Q sky130_fd_sc_hd__dfrtp_1
X_15658_ _15656_/Y _15657_/Y _15643_/X vssd1 vssd1 vccd1 vccd1 _15658_/X sky130_fd_sc_hd__o21a_1
X_18446_ _19855_/CLK _18446_/D vssd1 vssd1 vccd1 vccd1 _18446_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_221_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14609_ _18277_/Q _14599_/X _14580_/X _14602_/X vssd1 vssd1 vccd1 vccd1 _18277_/D
+ sky130_fd_sc_hd__a22o_1
X_18377_ _18441_/CLK _18377_/D vssd1 vssd1 vccd1 vccd1 _18377_/Q sky130_fd_sc_hd__dfxtp_1
X_15589_ _18590_/Q _15584_/A _18591_/Q vssd1 vssd1 vccd1 vccd1 _15589_/X sky130_fd_sc_hd__o21a_1
XFILLER_30_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19382__CLK _19920_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17328_ _17327_/X _13394_/Y _17535_/S vssd1 vssd1 vccd1 vccd1 _17328_/X sky130_fd_sc_hd__mux2_1
XFILLER_202_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17387__S _17487_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17259_ _16582_/Y _18977_/Q _17493_/S vssd1 vssd1 vccd1 vccd1 _17259_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12168__B1 _11909_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19194__RESET_B repeater188/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16854__A0 _17473_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08963_ _19852_/Q vssd1 vssd1 vccd1 vccd1 _10321_/B sky130_fd_sc_hd__inv_2
XANTENNA__13668__B1 hold259/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_229_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12340__B1 _12104_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_132_HCLK clkbuf_4_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19970_/CLK sky130_fd_sc_hd__clkbuf_16
X_09515_ _20017_/Q _19307_/Q _09477_/A _09514_/Y vssd1 vssd1 vccd1 vccd1 _09515_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_37_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17031__A0 _17473_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09446_ _19367_/Q vssd1 vssd1 vccd1 vccd1 _09446_/Y sky130_fd_sc_hd__inv_2
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09377_ _19926_/Q vssd1 vssd1 vccd1 vccd1 _10042_/A sky130_fd_sc_hd__inv_2
XFILLER_178_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09272__B1 _09082_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17297__S _17517_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12159__B1 _12107_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09024__B1 hold288/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11270_ _19599_/Q vssd1 vssd1 vccd1 vccd1 _11479_/A sky130_fd_sc_hd__inv_2
XFILLER_118_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10221_ _10219_/Y _19665_/Q _19838_/Q _10965_/A vssd1 vssd1 vccd1 vccd1 _10221_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_3_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16845__A0 _17486_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10152_ _10147_/X _19896_/Q _10152_/S vssd1 vssd1 vccd1 vccd1 _19896_/D sky130_fd_sc_hd__mux2_1
XFILLER_239_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13659__B1 hold233/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10083_ _10083_/A _10097_/A vssd1 vssd1 vccd1 vccd1 _10084_/B sky130_fd_sc_hd__or2_1
X_14960_ _18076_/Q _14953_/A _14933_/X _14954_/A vssd1 vssd1 vccd1 vccd1 _18076_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_48_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12331__B1 _12088_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18846__RESET_B repeater233/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13911_ _13911_/A _13911_/B _13911_/C _13911_/D vssd1 vssd1 vccd1 vccd1 _13912_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_102_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14891_ _18116_/Q _14884_/A _14814_/X _14885_/A vssd1 vssd1 vccd1 vccd1 _18116_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16073__A1 _17460_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17270__A0 _17473_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16073__B2 _15999_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16630_ _19283_/Q vssd1 vssd1 vccd1 vccd1 _16630_/Y sky130_fd_sc_hd__inv_2
XFILLER_207_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13842_ _19218_/Q _13914_/A _19207_/Q _13911_/B vssd1 vssd1 vccd1 vccd1 _13843_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_74_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16561_ _19040_/Q vssd1 vssd1 vccd1 vccd1 _16561_/Y sky130_fd_sc_hd__inv_2
X_13773_ _18738_/Q _18739_/Q _13775_/S vssd1 vssd1 vccd1 vccd1 _18739_/D sky130_fd_sc_hd__mux2_1
X_10985_ _10980_/B _10978_/X _10984_/Y _10408_/X _10964_/A vssd1 vssd1 vccd1 vccd1
+ _10986_/A sky130_fd_sc_hd__o32a_1
XFILLER_188_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17022__A0 _17486_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18300_ _18431_/CLK _18300_/D vssd1 vssd1 vccd1 vccd1 _18300_/Q sky130_fd_sc_hd__dfxtp_1
X_15512_ _15512_/A vssd1 vssd1 vccd1 vccd1 _15512_/X sky130_fd_sc_hd__clkbuf_2
X_12724_ _14812_/A _12709_/X _12723_/X _12711_/X vssd1 vssd1 vccd1 vccd1 _18955_/D
+ sky130_fd_sc_hd__a22o_1
X_19280_ _19283_/CLK _19280_/D repeater216/X vssd1 vssd1 vccd1 vccd1 _19280_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_15_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16492_ _16492_/A _16492_/B vssd1 vssd1 vccd1 vccd1 _16492_/X sky130_fd_sc_hd__or2_1
XANTENNA__17573__A1 _19770_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_231_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18231_ _18412_/CLK _18231_/D vssd1 vssd1 vccd1 vccd1 _18231_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15443_ _15443_/A _15443_/B vssd1 vssd1 vccd1 vccd1 _18551_/D sky130_fd_sc_hd__nor2_1
XFILLER_188_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12655_ _18995_/Q _12650_/X _12536_/X _12651_/X vssd1 vssd1 vccd1 vccd1 _18995_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10718__A _10718_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_repeater168_A _17548_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11606_ _11606_/A vssd1 vssd1 vccd1 vccd1 _11606_/Y sky130_fd_sc_hd__inv_2
XPHY_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18162_ _18954_/CLK _18162_/D vssd1 vssd1 vccd1 vccd1 _18162_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15374_ _19790_/Q _10650_/B _10651_/B vssd1 vssd1 vccd1 vccd1 _15374_/X sky130_fd_sc_hd__a21bo_1
XPHY_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12586_ _19040_/Q _12583_/X _12344_/X _12584_/X vssd1 vssd1 vccd1 vccd1 _19040_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19634__RESET_B repeater258/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17113_ _17112_/X _15628_/Y _17318_/S vssd1 vssd1 vccd1 vccd1 _17113_/X sky130_fd_sc_hd__mux2_2
XPHY_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14325_ _18438_/Q _14318_/X hold324/X _14320_/X vssd1 vssd1 vccd1 vccd1 _18438_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11537_ _11463_/A _11537_/A2 _11523_/X _11535_/Y vssd1 vssd1 vccd1 vccd1 _19582_/D
+ sky130_fd_sc_hd__a211oi_4
X_18093_ _18765_/CLK _18093_/D vssd1 vssd1 vccd1 vccd1 _18093_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16533__C1 _16532_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17000__S _17546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17044_ _17473_/A0 _16659_/Y _17547_/S vssd1 vssd1 vccd1 vccd1 _17044_/X sky130_fd_sc_hd__mux2_1
XANTENNA_output97_A _16698_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14256_ _14256_/A _14489_/B _15318_/B vssd1 vssd1 vccd1 vccd1 _15034_/C sky130_fd_sc_hd__or3_4
XFILLER_128_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11468_ _11468_/A _11468_/B _11468_/C vssd1 vssd1 vccd1 vccd1 _11525_/A sky130_fd_sc_hd__or3_1
Xclkbuf_leaf_13_HCLK clkbuf_4_2_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20123_/CLK sky130_fd_sc_hd__clkbuf_16
X_13207_ _13207_/A vssd1 vssd1 vccd1 vccd1 _13207_/Y sky130_fd_sc_hd__clkinv_1
X_10419_ _10419_/A vssd1 vssd1 vccd1 vccd1 _10419_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14187_ _19120_/Q vssd1 vssd1 vccd1 vccd1 _14187_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11399_ _19554_/Q _11396_/Y _11624_/A _19134_/Q _11398_/X vssd1 vssd1 vccd1 vccd1
+ _11412_/B sky130_fd_sc_hd__o221a_1
XFILLER_225_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13138_ _13136_/Y _18912_/Q _13137_/Y _18898_/Q vssd1 vssd1 vccd1 vccd1 _13138_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__15963__B _17537_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18995_ _19137_/CLK _18995_/D repeater249/X vssd1 vssd1 vccd1 vccd1 _18995_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_140_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13069_ _13069_/A _13069_/B _13069_/C vssd1 vssd1 vccd1 vccd1 _13070_/B sky130_fd_sc_hd__or3_1
X_17946_ _18260_/CLK _17946_/D vssd1 vssd1 vccd1 vccd1 _17946_/Q sky130_fd_sc_hd__dfxtp_1
Xrepeater204 repeater205/X vssd1 vssd1 vccd1 vccd1 repeater204/X sky130_fd_sc_hd__clkbuf_8
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11125__A1 _19634_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_227_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater215 repeater216/X vssd1 vssd1 vccd1 vccd1 repeater215/X sky130_fd_sc_hd__buf_4
XANTENNA__12322__B1 _12069_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater226 repeater227/X vssd1 vssd1 vccd1 vccd1 repeater226/X sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_155_HCLK clkbuf_4_1_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _18431_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__18587__RESET_B repeater271/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater237 repeater239/X vssd1 vssd1 vccd1 vccd1 repeater237/X sky130_fd_sc_hd__buf_6
XFILLER_94_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater248 hold370/A vssd1 vssd1 vccd1 vccd1 hold371/A sky130_fd_sc_hd__buf_6
XFILLER_120_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17877_ _16105_/Y _16106_/Y _16107_/Y _16108_/Y _17908_/S0 _18759_/Q vssd1 vssd1
+ vccd1 vccd1 _17877_/X sky130_fd_sc_hd__mux4_1
Xrepeater259 repeater260/X vssd1 vssd1 vccd1 vccd1 repeater259/X sky130_fd_sc_hd__buf_6
XANTENNA__17261__A0 _17486_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17670__S _17683_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19616_ _19937_/CLK _19616_/D repeater190/X vssd1 vssd1 vccd1 vccd1 _19616_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_241_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16828_ _16719_/Y _20120_/Q _17385_/S vssd1 vssd1 vccd1 vccd1 _16828_/X sky130_fd_sc_hd__mux2_1
XANTENNA__19748__CLK _20070_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19547_ _19576_/CLK _19547_/D repeater282/X vssd1 vssd1 vccd1 vccd1 _19547_/Q sky130_fd_sc_hd__dfrtp_1
X_16759_ vssd1 vssd1 vccd1 vccd1 _16759_/HI _16759_/LO sky130_fd_sc_hd__conb_1
X_09300_ _18654_/Q _18655_/Q _18656_/Q _18657_/Q vssd1 vssd1 vccd1 vccd1 _09329_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_62_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19478_ _19506_/CLK hold188/X repeater256/X vssd1 vssd1 vccd1 vccd1 _19478_/Q sky130_fd_sc_hd__dfrtp_1
X_09231_ _09231_/A vssd1 vssd1 vccd1 vccd1 _15710_/A sky130_fd_sc_hd__inv_2
X_18429_ _18795_/CLK _18429_/D vssd1 vssd1 vccd1 vccd1 _18429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_221_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19898__CLK _19900_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09162_ _09162_/A _15319_/A vssd1 vssd1 vccd1 vccd1 _09164_/A sky130_fd_sc_hd__or2_4
XFILLER_119_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16524__C1 _16523_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09093_ _14791_/A vssd1 vssd1 vccd1 vccd1 _12232_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_163_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15873__B _15878_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18152__CLK _18169_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09995_ _09995_/A vssd1 vssd1 vccd1 vccd1 _09995_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13674__A hold325/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08946_ _18773_/Q vssd1 vssd1 vccd1 vccd1 _08946_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17580__S _17584_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_hold163_A HADDR[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11922__A _13678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10770_ _19750_/Q _10766_/B _10758_/B _10761_/A vssd1 vssd1 vccd1 vccd1 _19750_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_40_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16209__B _16212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09429_ _19906_/Q vssd1 vssd1 vccd1 vccd1 _10013_/A sky130_fd_sc_hd__inv_2
XFILLER_240_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16924__S _17414_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12440_ _12478_/A vssd1 vssd1 vccd1 vccd1 _12457_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__17307__A1 _13845_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_36_HCLK _18641_/CLK vssd1 vssd1 vccd1 vccd1 _20081_/CLK sky130_fd_sc_hd__clkbuf_16
X_12371_ _12371_/A _15902_/A vssd1 vssd1 vccd1 vccd1 _12659_/B sky130_fd_sc_hd__or2_2
XFILLER_193_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14110_ _14026_/A _14110_/A2 _14108_/Y _14135_/B vssd1 vssd1 vccd1 vccd1 _18696_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_176_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11322_ _11484_/A _18986_/Q _19589_/Q _11321_/Y vssd1 vssd1 vccd1 vccd1 _11322_/X
+ sky130_fd_sc_hd__o22a_1
X_15090_ _17997_/Q _15083_/X _14793_/X _15085_/X vssd1 vssd1 vccd1 vccd1 _17997_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_181_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14041_ _14038_/Y _18690_/Q _19084_/Q _14025_/A _14040_/X vssd1 vssd1 vccd1 vccd1
+ _14049_/B sky130_fd_sc_hd__a221o_1
X_11253_ _19004_/Q vssd1 vssd1 vccd1 vccd1 _11253_/Y sky130_fd_sc_hd__inv_2
X_10204_ _19658_/Q vssd1 vssd1 vccd1 vccd1 _10958_/A sky130_fd_sc_hd__inv_2
XFILLER_79_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11184_ _11191_/A vssd1 vssd1 vccd1 vccd1 _11184_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_192_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17491__A0 _17490_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17800_ _18330_/Q _18210_/Q _18202_/Q _18194_/Q _17918_/S0 _18750_/Q vssd1 vssd1
+ vccd1 vccd1 _17800_/X sky130_fd_sc_hd__mux4_2
XFILLER_121_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_192_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10135_ _10136_/A vssd1 vssd1 vccd1 vccd1 _10138_/A sky130_fd_sc_hd__inv_2
X_18780_ _19855_/CLK _18780_/D repeater265/X vssd1 vssd1 vccd1 vccd1 _18780_/Q sky130_fd_sc_hd__dfrtp_1
X_15992_ _15990_/Y _15884_/X _15991_/Y _15915_/X vssd1 vssd1 vccd1 vccd1 _15992_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_209_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12304__B1 _12232_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18680__RESET_B hold359/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17731_ _15378_/X _19714_/Q _18508_/D vssd1 vssd1 vccd1 vccd1 _17731_/X sky130_fd_sc_hd__mux2_1
X_10066_ _19927_/Q _10065_/Y _10057_/X _10044_/B vssd1 vssd1 vccd1 vccd1 _19927_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_76_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14943_ _18088_/Q _14939_/X _14925_/X _14941_/X vssd1 vssd1 vccd1 vccd1 _18088_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_output135_A _15732_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_208_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17243__A0 _17242_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17490__S _17490_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14874_ _18129_/Q _14871_/X _14699_/X _14873_/X vssd1 vssd1 vccd1 vccd1 _18129_/D
+ sky130_fd_sc_hd__a22o_1
X_17662_ _15586_/Y _19027_/Q _17664_/S vssd1 vssd1 vccd1 vccd1 _18590_/D sky130_fd_sc_hd__mux2_1
XFILLER_36_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19401_ _19976_/CLK _19401_/D hold371/X vssd1 vssd1 vccd1 vccd1 _19401_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_35_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16613_ _16869_/X _16577_/X _17004_/X _16578_/X _16612_/X vssd1 vssd1 vccd1 vccd1
+ _16614_/C sky130_fd_sc_hd__o221a_1
X_13825_ _13912_/D _13825_/B vssd1 vssd1 vccd1 vccd1 _13924_/A sky130_fd_sc_hd__or2_1
XFILLER_235_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17593_ _15351_/X _19710_/Q _17600_/S vssd1 vssd1 vccd1 vccd1 _17593_/X sky130_fd_sc_hd__mux2_1
XFILLER_211_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09005__C _11842_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11832__A _15823_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19332_ _19956_/CLK _19332_/D repeater245/X vssd1 vssd1 vccd1 vccd1 _19332_/Q sky130_fd_sc_hd__dfrtp_1
X_16544_ _16544_/A _16544_/B vssd1 vssd1 vccd1 vccd1 _16544_/Y sky130_fd_sc_hd__nor2_1
X_13756_ _13756_/A _13756_/B vssd1 vssd1 vccd1 vccd1 _13757_/A sky130_fd_sc_hd__nand2_1
XFILLER_44_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10968_ _10968_/A vssd1 vssd1 vccd1 vccd1 _10968_/Y sky130_fd_sc_hd__inv_2
XFILLER_149_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12707_ _18959_/Q vssd1 vssd1 vccd1 vccd1 _14802_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_203_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16475_ _08962_/Y _16505_/A _10236_/Y _16506_/A vssd1 vssd1 vccd1 vccd1 _16475_/X
+ sky130_fd_sc_hd__o22a_1
X_19263_ _19283_/CLK _19263_/D repeater212/X vssd1 vssd1 vccd1 vccd1 _19263_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__16834__S _17386_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13687_ _18771_/Q _13685_/X _13674_/X _13686_/Y vssd1 vssd1 vccd1 vccd1 _18771_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10448__A _10448_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10899_ _19689_/Q _10893_/X _10861_/X _10895_/X vssd1 vssd1 vccd1 vccd1 _19689_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_203_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15426_ _19617_/Q _11162_/B _11163_/B vssd1 vssd1 vccd1 vccd1 _15426_/X sky130_fd_sc_hd__a21bo_1
X_18214_ _19630_/CLK _18214_/D vssd1 vssd1 vccd1 vccd1 _18214_/Q sky130_fd_sc_hd__dfxtp_1
X_12638_ _19008_/Q _12636_/X _12413_/X _12637_/X vssd1 vssd1 vccd1 vccd1 _19008_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19194_ _19214_/CLK _19194_/D repeater188/X vssd1 vssd1 vccd1 vccd1 _19194_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15958__B _16344_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15357_ _18500_/Q _14230_/B _14231_/B vssd1 vssd1 vccd1 vccd1 _15357_/X sky130_fd_sc_hd__a21bo_1
X_18145_ _18145_/CLK _18145_/D vssd1 vssd1 vccd1 vccd1 _18145_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12663__A _12699_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12569_ _12576_/A vssd1 vssd1 vccd1 vccd1 _12569_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_184_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16135__A _19773_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14308_ _18447_/Q _14303_/X _14279_/X _14305_/X vssd1 vssd1 vccd1 vccd1 _18447_/D
+ sky130_fd_sc_hd__a22o_1
X_18076_ _18198_/CLK _18076_/D vssd1 vssd1 vccd1 vccd1 _18076_/Q sky130_fd_sc_hd__dfxtp_1
X_15288_ _19780_/Q _18517_/D _15268_/C _15254_/Y _10754_/A vssd1 vssd1 vccd1 vccd1
+ _15289_/B sky130_fd_sc_hd__o32a_1
XFILLER_172_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold206 input26/X vssd1 vssd1 vccd1 vccd1 hold206/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__18175__CLK _18198_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold217 hold217/A vssd1 vssd1 vccd1 vccd1 hold217/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold228 hold228/A vssd1 vssd1 vccd1 vccd1 hold228/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17665__S _17683_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17027_ _16472_/Y _19409_/Q _17523_/S vssd1 vssd1 vccd1 vccd1 _17027_/X sky130_fd_sc_hd__mux2_1
X_14239_ _18668_/Q _14236_/X _18507_/Q _17600_/S vssd1 vssd1 vccd1 vccd1 _18668_/D
+ sky130_fd_sc_hd__a22o_1
Xhold239 hold239/A vssd1 vssd1 vccd1 vccd1 hold239/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09780_ _09744_/A _09744_/B _09734_/A _09778_/Y vssd1 vssd1 vccd1 vccd1 _19988_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_140_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18978_ _19600_/CLK _18978_/D hold273/X vssd1 vssd1 vccd1 vccd1 _18978_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__14296__B1 _13678_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_239_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17929_ _18623_/CLK hold368/X vssd1 vssd1 vccd1 vccd1 _17929_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_239_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17234__A0 _17486_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_227_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_242_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17880__S1 _19632_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11742__A _11742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17537__A1 _13021_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_6_0_HCLK_A clkbuf_4_7_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_59_HCLK clkbuf_4_12_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19971_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__19556__RESET_B hold346/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_201_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09214_ _18650_/Q _09214_/B vssd1 vssd1 vccd1 vccd1 _09214_/Y sky130_fd_sc_hd__nand2_1
XFILLER_195_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14220__B1 _18671_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09145_ _09138_/A _17605_/S _17603_/X vssd1 vssd1 vccd1 vccd1 _09146_/A sky130_fd_sc_hd__a21oi_2
XFILLER_175_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12782__B1 _19233_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09076_ _20101_/Q _09069_/X _09075_/X _09072_/X vssd1 vssd1 vccd1 vccd1 _20101_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_30_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17575__S _17584_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12534__B1 _12533_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17473__A0 _17473_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15079__A2 _15072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold280_A HWDATA[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09978_ _09978_/A vssd1 vssd1 vccd1 vccd1 _09978_/Y sky130_fd_sc_hd__inv_2
X_08929_ _19866_/Q vssd1 vssd1 vccd1 vccd1 _10332_/A sky130_fd_sc_hd__inv_2
XFILLER_58_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20098_ _20107_/CLK _20098_/D repeater234/X vssd1 vssd1 vccd1 vccd1 _20098_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__16919__S _17482_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10848__B1 _10451_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11940_ _11977_/A vssd1 vssd1 vccd1 vccd1 _11979_/A sky130_fd_sc_hd__inv_2
XANTENNA__16579__A2 _15889_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_217_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11871_ _12130_/A _11935_/B _12256_/C vssd1 vssd1 vccd1 vccd1 _15888_/A sky130_fd_sc_hd__or3_1
XANTENNA__17871__S1 _19632_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_232_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13610_ _13610_/A vssd1 vssd1 vccd1 vccd1 _13610_/Y sky130_fd_sc_hd__inv_2
X_10822_ _10831_/B vssd1 vssd1 vccd1 vccd1 _17750_/S sky130_fd_sc_hd__inv_2
XFILLER_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14590_ _18289_/Q _14587_/X _14531_/X _14589_/X vssd1 vssd1 vccd1 vccd1 _18289_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_32_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_232_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19297__RESET_B repeater241/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13541_ _13541_/A _13541_/B vssd1 vssd1 vccd1 vccd1 _13586_/A sky130_fd_sc_hd__or2_1
X_10753_ _18519_/Q _15436_/A vssd1 vssd1 vccd1 vccd1 _10754_/A sky130_fd_sc_hd__nand2_1
XFILLER_186_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10268__A _19647_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19226__RESET_B repeater257/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_200_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16260_ _18167_/Q vssd1 vssd1 vccd1 vccd1 _16260_/Y sky130_fd_sc_hd__inv_2
X_13472_ _13470_/A _13470_/B _13470_/Y _13437_/X vssd1 vssd1 vccd1 vccd1 _18847_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_201_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_200_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18198__CLK _18198_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10684_ _11842_/D vssd1 vssd1 vccd1 vccd1 _15858_/C sky130_fd_sc_hd__buf_1
X_15211_ _15211_/A _15215_/B vssd1 vssd1 vccd1 vccd1 _15211_/Y sky130_fd_sc_hd__nor2_1
X_12423_ _19136_/Q _12420_/X _12356_/X _12421_/X vssd1 vssd1 vccd1 vccd1 _19136_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19443__CLK _19992_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16191_ _17957_/Q vssd1 vssd1 vccd1 vccd1 _16191_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15142_ _17963_/Q _15135_/A _10423_/A _15136_/A vssd1 vssd1 vccd1 vccd1 _17963_/D
+ sky130_fd_sc_hd__a22o_1
X_12354_ _12362_/A vssd1 vssd1 vccd1 vccd1 _12354_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_138_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17485__S _17536_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11305_ _18979_/Q vssd1 vssd1 vccd1 vccd1 _11305_/Y sky130_fd_sc_hd__inv_2
XFILLER_114_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15073_ _15073_/A vssd1 vssd1 vccd1 vccd1 _15073_/X sky130_fd_sc_hd__clkbuf_2
X_19950_ _19964_/CLK _19950_/D hold371/X vssd1 vssd1 vccd1 vccd1 _19950_/Q sky130_fd_sc_hd__dfrtp_1
X_12285_ _19209_/Q _12283_/X _12107_/X _12284_/X vssd1 vssd1 vccd1 vccd1 _19209_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_107_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18861__RESET_B repeater231/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14024_ _14024_/A _14024_/B vssd1 vssd1 vccd1 vccd1 _14111_/A sky130_fd_sc_hd__or2_1
X_18901_ _19352_/CLK _18901_/D repeater188/X vssd1 vssd1 vccd1 vccd1 _18901_/Q sky130_fd_sc_hd__dfrtp_1
X_11236_ _18993_/Q vssd1 vssd1 vccd1 vccd1 _11236_/Y sky130_fd_sc_hd__inv_2
X_19881_ _20050_/CLK _19881_/D repeater200/X vssd1 vssd1 vccd1 vccd1 _19881_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_150_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18832_ _19255_/CLK _18832_/D repeater237/X vssd1 vssd1 vccd1 vccd1 _18832_/Q sky130_fd_sc_hd__dfrtp_1
X_11167_ _19622_/Q _11167_/B vssd1 vssd1 vccd1 vccd1 _11168_/B sky130_fd_sc_hd__or2_1
XANTENNA__14278__B1 _14277_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10118_ _18566_/Q _15481_/A vssd1 vssd1 vccd1 vccd1 _15486_/A sky130_fd_sc_hd__or2_1
XFILLER_121_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18763_ _20123_/CLK _18763_/D repeater195/X vssd1 vssd1 vccd1 vccd1 _18763_/Q sky130_fd_sc_hd__dfrtp_4
X_15975_ _19674_/Q vssd1 vssd1 vccd1 vccd1 _15975_/Y sky130_fd_sc_hd__inv_2
X_11098_ _14963_/B _14476_/A _10400_/B vssd1 vssd1 vccd1 vccd1 _11098_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__16829__S _17386_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17216__A0 _17486_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17714_ _15426_/X _19527_/Q _18546_/D vssd1 vssd1 vccd1 vccd1 _17714_/X sky130_fd_sc_hd__mux2_1
X_10049_ _10049_/A vssd1 vssd1 vccd1 vccd1 _10049_/Y sky130_fd_sc_hd__inv_2
X_14926_ _18096_/Q _14920_/X _14925_/X _14923_/X vssd1 vssd1 vccd1 vccd1 _18096_/D
+ sky130_fd_sc_hd__a22o_1
X_18694_ _19119_/CLK _18694_/D hold351/X vssd1 vssd1 vccd1 vccd1 _18694_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_209_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17645_ _15658_/X _19044_/Q _17655_/S vssd1 vssd1 vccd1 vccd1 _18607_/D sky130_fd_sc_hd__mux2_1
XANTENNA__17862__S1 _19632_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14857_ _14857_/A _15109_/B _15145_/C vssd1 vssd1 vccd1 vccd1 _14859_/A sky130_fd_sc_hd__or3_4
X_13808_ _18713_/Q vssd1 vssd1 vccd1 vccd1 _13950_/A sky130_fd_sc_hd__inv_2
X_17576_ _15408_/X _19767_/Q _17584_/S vssd1 vssd1 vccd1 vccd1 _17576_/X sky130_fd_sc_hd__mux2_1
X_14788_ _18177_/Q _14785_/X _14745_/X _14787_/X vssd1 vssd1 vccd1 vccd1 _18177_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_90_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17519__A1 _09807_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19315_ _19315_/CLK _19315_/D repeater214/X vssd1 vssd1 vccd1 vccd1 _19315_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_50_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_220_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16527_ _17106_/X _16505_/X _17276_/X _16506_/X vssd1 vssd1 vccd1 vccd1 _16527_/X
+ sky130_fd_sc_hd__o22a_1
X_13739_ _18752_/Q _13741_/A _13255_/Y _13738_/A vssd1 vssd1 vccd1 vccd1 _18752_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_176_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19246_ _19320_/CLK _19246_/D repeater214/X vssd1 vssd1 vccd1 vccd1 _19246_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_176_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16458_ _17310_/X _15884_/A _17309_/X _15915_/A vssd1 vssd1 vccd1 vccd1 _16458_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__14202__B1 _19122_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16742__A2 _15904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15409_ _15413_/A _17576_/X vssd1 vssd1 vccd1 vccd1 _18536_/D sky130_fd_sc_hd__and2_1
X_19177_ _19288_/CLK _19177_/D repeater212/X vssd1 vssd1 vccd1 vccd1 _19177_/Q sky130_fd_sc_hd__dfrtp_1
X_16389_ _17340_/X _15884_/A _17339_/X _15915_/A vssd1 vssd1 vccd1 vccd1 _16389_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_185_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18810__CLK _20115_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18128_ _20090_/CLK _18128_/D vssd1 vssd1 vccd1 vccd1 _18128_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17395__S _17564_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18059_ _18460_/CLK _18059_/D vssd1 vssd1 vccd1 vccd1 _18059_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12516__B1 hold281/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09901_ _19342_/Q vssd1 vssd1 vccd1 vccd1 _09901_/Y sky130_fd_sc_hd__inv_2
XFILLER_160_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20021_ _20032_/CLK _20021_/D repeater238/X vssd1 vssd1 vccd1 vccd1 _20021_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17455__A0 _15768_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09832_ _19954_/Q vssd1 vssd1 vccd1 vccd1 _09862_/A sky130_fd_sc_hd__inv_2
XFILLER_113_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_246_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09763_ _09848_/B vssd1 vssd1 vccd1 vccd1 _09763_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_132_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09694_ _19410_/Q vssd1 vssd1 vccd1 vccd1 _09694_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrebuffer10 _13075_/B vssd1 vssd1 vccd1 vccd1 _13189_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_4007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer21 _14012_/C vssd1 vssd1 vccd1 vccd1 _14136_/A sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_94_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19737__RESET_B repeater207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer32 _11566_/B vssd1 vssd1 vccd1 vccd1 _11543_/A sky130_fd_sc_hd__dlygate4sd1_1
XPHY_4029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer43 _11468_/C vssd1 vssd1 vccd1 vccd1 _11530_/A2 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer54 _11467_/B vssd1 vssd1 vccd1 vccd1 _11531_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XANTENNA__17853__S1 _19632_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_242_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_214_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrebuffer65 _13064_/B vssd1 vssd1 vccd1 vccd1 _13209_/A2 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer76 _13419_/A vssd1 vssd1 vccd1 vccd1 _13423_/A sky130_fd_sc_hd__dlygate4sd1_1
XPHY_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_242_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_214_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13244__A1 _15419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrebuffer87 _14028_/B vssd1 vssd1 vccd1 vccd1 _14107_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrebuffer98 _14026_/B vssd1 vssd1 vccd1 vccd1 _14110_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16733__A2 _16513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrebuffer100 _11482_/B vssd1 vssd1 vccd1 vccd1 _11502_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_195_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrebuffer111 _09858_/B vssd1 vssd1 vccd1 vccd1 _09984_/A sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_195_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrebuffer122 _09857_/C vssd1 vssd1 vccd1 vccd1 _09989_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_109_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09128_ _15321_/B _09162_/A _17602_/X _09127_/X vssd1 vssd1 vccd1 vccd1 _09136_/B
+ sky130_fd_sc_hd__or4b_4
XFILLER_135_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18619__RESET_B repeater269/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16497__B2 _15908_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09059_ _20106_/Q _09053_/X _09058_/X _09055_/X vssd1 vssd1 vccd1 vccd1 _20106_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12507__B1 _12401_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12070_ _12121_/A vssd1 vssd1 vccd1 vccd1 _12122_/A sky130_fd_sc_hd__inv_2
XFILLER_132_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17446__A0 _15963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16249__A1 _11742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11021_ _19653_/Q _10955_/Y _10954_/A _10211_/X vssd1 vssd1 vccd1 vccd1 _19653_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_89_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_238_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_246_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15760_ _18527_/D vssd1 vssd1 vccd1 vccd1 _15765_/C sky130_fd_sc_hd__inv_2
X_12972_ _12972_/A vssd1 vssd1 vccd1 vccd1 _12972_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17749__A1 _18879_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14711_ _14711_/A vssd1 vssd1 vccd1 vccd1 _14711_/X sky130_fd_sc_hd__clkbuf_2
X_11923_ _19403_/Q _11914_/X _11922_/X _11915_/X vssd1 vssd1 vccd1 vccd1 _19403_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_233_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15691_ _15690_/Y _15687_/A _18615_/Q _15687_/Y _15643_/A vssd1 vssd1 vccd1 vccd1
+ _15691_/X sky130_fd_sc_hd__o221a_1
XANTENNA__17844__S1 _19634_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12478__A _12478_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17430_ _17429_/X _16113_/Y _17565_/S vssd1 vssd1 vccd1 vccd1 _17430_/X sky130_fd_sc_hd__mux2_1
X_14642_ _14642_/A _14668_/B _14951_/C vssd1 vssd1 vccd1 vccd1 _14644_/A sky130_fd_sc_hd__or3_4
XPHY_4563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11854_ _11869_/A _13641_/B vssd1 vssd1 vccd1 vccd1 _11855_/A sky130_fd_sc_hd__or2_1
XFILLER_61_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14432__B1 _14419_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10805_ _10805_/A _18653_/Q vssd1 vssd1 vccd1 vccd1 _10806_/A sky130_fd_sc_hd__or2_1
XFILLER_202_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14573_ _14573_/A vssd1 vssd1 vccd1 vccd1 _14574_/A sky130_fd_sc_hd__inv_2
X_17361_ _17360_/X _12945_/Y _17487_/S vssd1 vssd1 vccd1 vccd1 _17361_/X sky130_fd_sc_hd__mux2_1
XPHY_3873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11785_ _11821_/A vssd1 vssd1 vccd1 vccd1 _11822_/A sky130_fd_sc_hd__inv_2
XPHY_3884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19060__RESET_B repeater257/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19100_ _19109_/CLK _19100_/D hold361/X vssd1 vssd1 vccd1 vccd1 _19100_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_3895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16312_ _19526_/Q vssd1 vssd1 vccd1 vccd1 _16312_/Y sky130_fd_sc_hd__inv_2
X_13524_ _14642_/A _14668_/B _13506_/A _14857_/A _13523_/Y vssd1 vssd1 vccd1 vccd1
+ _13524_/X sky130_fd_sc_hd__o32a_1
X_10736_ _10736_/A _10736_/B vssd1 vssd1 vccd1 vccd1 _10736_/X sky130_fd_sc_hd__or2_1
XFILLER_14_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17292_ _17291_/X _15491_/A _17513_/S vssd1 vssd1 vccd1 vccd1 _17292_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16724__A2 _15887_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19031_ _19855_/CLK _19031_/D repeater265/X vssd1 vssd1 vccd1 vccd1 _19031_/Q sky130_fd_sc_hd__dfrtp_1
X_16243_ _17394_/X _15883_/A _17393_/X _15914_/A vssd1 vssd1 vccd1 vccd1 _16243_/X
+ sky130_fd_sc_hd__o22a_2
X_13455_ _13429_/D _13340_/B _13453_/Y _13445_/X vssd1 vssd1 vccd1 vccd1 _18853_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_174_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10667_ _17732_/X _10661_/X _19793_/Q _10663_/X vssd1 vssd1 vccd1 vccd1 _19793_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_repeater150_A _17487_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12406_ hold318/X vssd1 vssd1 vccd1 vccd1 _12406_/X sky130_fd_sc_hd__clkbuf_2
X_16174_ _19846_/Q vssd1 vssd1 vccd1 vccd1 _16174_/Y sky130_fd_sc_hd__inv_2
XFILLER_127_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13386_ _13376_/X _13386_/B _13386_/C _13386_/D vssd1 vssd1 vccd1 vccd1 _13418_/B
+ sky130_fd_sc_hd__and4b_1
X_10598_ _10598_/A vssd1 vssd1 vccd1 vccd1 _10598_/Y sky130_fd_sc_hd__inv_2
X_15125_ _17976_/Q _15122_/X _14921_/X _15124_/X vssd1 vssd1 vccd1 vccd1 _17976_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_217_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput108 _16465_/Y vssd1 vssd1 vccd1 vccd1 HRDATA[7] sky130_fd_sc_hd__clkbuf_2
X_12337_ _19178_/Q _12334_/X _12098_/X _12335_/X vssd1 vssd1 vccd1 vccd1 _19178_/D
+ sky130_fd_sc_hd__a22o_1
Xoutput119 _16750_/Y vssd1 vssd1 vccd1 vccd1 IRQ[1] sky130_fd_sc_hd__clkbuf_2
XANTENNA__17780__S0 _17923_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19933_ _19933_/CLK _19933_/D repeater236/X vssd1 vssd1 vccd1 vccd1 _19933_/Q sky130_fd_sc_hd__dfrtp_4
X_15056_ _18019_/Q _15048_/A _15006_/X _15049_/A vssd1 vssd1 vccd1 vccd1 _18019_/D
+ sky130_fd_sc_hd__a22o_1
X_12268_ _19220_/Q _12260_/X _12080_/X _12263_/X vssd1 vssd1 vccd1 vccd1 _19220_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_130_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14007_ _14007_/A _14007_/B vssd1 vssd1 vccd1 vccd1 _14142_/A sky130_fd_sc_hd__or2_1
XFILLER_96_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11219_ _19585_/Q vssd1 vssd1 vccd1 vccd1 _11466_/A sky130_fd_sc_hd__inv_2
X_19864_ _19865_/CLK _19864_/D repeater267/X vssd1 vssd1 vccd1 vccd1 _19864_/Q sky130_fd_sc_hd__dfrtp_1
X_12199_ _12206_/A vssd1 vssd1 vccd1 vccd1 _12199_/X sky130_fd_sc_hd__buf_1
XFILLER_233_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput90 _16006_/Y vssd1 vssd1 vccd1 vccd1 HRDATA[1] sky130_fd_sc_hd__clkbuf_2
XFILLER_110_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18815_ _20115_/CLK _18815_/D repeater239/X vssd1 vssd1 vccd1 vccd1 _18815_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__09027__A hold286/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19795_ _19795_/CLK _19795_/D repeater219/X vssd1 vssd1 vccd1 vccd1 _19795_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_56_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16660__A1 _16974_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18746_ _20036_/CLK _18746_/D repeater199/X vssd1 vssd1 vccd1 vccd1 _18746_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_83_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15958_ _17938_/Q _16344_/B vssd1 vssd1 vccd1 vccd1 _15958_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_156_HCLK_A clkbuf_4_1_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19830__RESET_B repeater270/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_224_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14909_ _14909_/A vssd1 vssd1 vccd1 vccd1 _14910_/A sky130_fd_sc_hd__inv_2
XANTENNA__17835__S1 _18759_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18677_ _18686_/CLK _18677_/D repeater252/X vssd1 vssd1 vccd1 vccd1 _18677_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__12388__A _12400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15889_ _16637_/A vssd1 vssd1 vccd1 vccd1 _15889_/X sky130_fd_sc_hd__buf_2
XANTENNA__11292__A _18994_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17628_ _19891_/Q _19744_/Q _17630_/S vssd1 vssd1 vccd1 vccd1 _17628_/X sky130_fd_sc_hd__mux2_1
XFILLER_224_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13777__A2 _13202_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17559_ _15820_/Y _15819_/Y _17564_/S vssd1 vssd1 vccd1 vccd1 _17559_/X sky130_fd_sc_hd__mux2_1
XFILLER_220_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19229_ _19314_/CLK _19229_/D repeater214/X vssd1 vssd1 vccd1 vccd1 _19229_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_118_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18712__RESET_B repeater253/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17771__S0 _17923_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15151__B2 _15148_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19989__RESET_B repeater192/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_207_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11712__A1 _15858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19918__RESET_B repeater230/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20004_ _20091_/CLK _20004_/D repeater236/X vssd1 vssd1 vccd1 vccd1 _20004_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__11712__B2 _16950_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09815_ _19326_/Q vssd1 vssd1 vccd1 vccd1 _09815_/Y sky130_fd_sc_hd__inv_2
XFILLER_247_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_228_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13682__A _14405_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09746_ _09746_/A _09746_/B vssd1 vssd1 vccd1 vccd1 _09775_/A sky130_fd_sc_hd__or2_1
XFILLER_27_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_227_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09677_ _19432_/Q vssd1 vssd1 vccd1 vccd1 _09677_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17826__S1 _18750_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_15_HCLK_A clkbuf_4_2_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_hold243_A RsRx_S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_78_HCLK_A clkbuf_4_13_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_3_HCLK_A clkbuf_4_0_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10249__C _12053_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11570_ _11570_/A _11570_/B vssd1 vssd1 vccd1 vccd1 _11571_/B sky130_fd_sc_hd__or2_2
XPHY_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16217__B _17473_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10521_ _19532_/Q _19531_/Q _10521_/C vssd1 vssd1 vccd1 vccd1 _10734_/C sky130_fd_sc_hd__or3_1
XFILLER_183_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16932__S _16946_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13240_ _15973_/A _13252_/D vssd1 vssd1 vccd1 vccd1 _13242_/A sky130_fd_sc_hd__or2_2
XFILLER_182_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10452_ _10452_/A vssd1 vssd1 vccd1 vccd1 _10452_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_136_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_182_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13171_ _13085_/A _13171_/A2 _13202_/A _13169_/Y vssd1 vssd1 vccd1 vccd1 _18913_/D
+ sky130_fd_sc_hd__a211oi_4
X_10383_ _19853_/Q _19852_/Q _19854_/Q _10382_/X vssd1 vssd1 vccd1 vccd1 _10383_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_109_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_184_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12122_ _12122_/A vssd1 vssd1 vccd1 vccd1 _12122_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_151_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12053_ _15233_/A _12053_/B vssd1 vssd1 vccd1 vccd1 _12053_/Y sky130_fd_sc_hd__nor2_1
X_16930_ _19474_/Q hold206/X _16950_/S vssd1 vssd1 vccd1 vccd1 _16930_/X sky130_fd_sc_hd__mux2_4
XFILLER_117_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11004_ _11004_/A vssd1 vssd1 vccd1 vccd1 _19659_/D sky130_fd_sc_hd__inv_2
XANTENNA__19659__RESET_B repeater270/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16861_ _16860_/X _15517_/Y _17513_/S vssd1 vssd1 vccd1 vccd1 _16861_/X sky130_fd_sc_hd__mux2_1
XFILLER_238_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18600_ _19867_/CLK _18600_/D repeater263/X vssd1 vssd1 vccd1 vccd1 _18600_/Q sky130_fd_sc_hd__dfrtp_4
X_15812_ _18258_/Q vssd1 vssd1 vccd1 vccd1 _15812_/Y sky130_fd_sc_hd__inv_2
X_19580_ _19591_/CLK _19580_/D hold346/X vssd1 vssd1 vccd1 vccd1 _19580_/Q sky130_fd_sc_hd__dfrtp_1
X_16792_ _16791_/X _16736_/Y _17490_/S vssd1 vssd1 vccd1 vccd1 _16792_/X sky130_fd_sc_hd__mux2_2
XFILLER_133_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18531_ _19937_/CLK _18531_/D repeater189/X vssd1 vssd1 vccd1 vccd1 _18531_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_46_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_246_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15743_ _15747_/C _18488_/D _18489_/Q vssd1 vssd1 vccd1 vccd1 _18484_/D sky130_fd_sc_hd__and3_1
XFILLER_218_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12955_ _12944_/X _12955_/B _12955_/C _12955_/D vssd1 vssd1 vccd1 vccd1 _12956_/D
+ sky130_fd_sc_hd__and4b_1
XFILLER_46_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17817__S1 _18750_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19241__RESET_B repeater239/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11906_ _11915_/A vssd1 vssd1 vccd1 vccd1 _11906_/X sky130_fd_sc_hd__buf_1
X_18462_ _19842_/CLK _18462_/D vssd1 vssd1 vccd1 vccd1 _18462_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_234_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15674_ _18611_/Q _15669_/Y _15672_/Y _15669_/A _15673_/X vssd1 vssd1 vccd1 vccd1
+ _15674_/X sky130_fd_sc_hd__o221a_1
X_12886_ _18945_/Q vssd1 vssd1 vccd1 vccd1 _12887_/C sky130_fd_sc_hd__inv_2
XPHY_4360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17413_ _17412_/X _16119_/Y _17413_/S vssd1 vssd1 vccd1 vccd1 _17413_/X sky130_fd_sc_hd__mux2_1
XPHY_4393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14625_ _18267_/Q _14617_/A _09185_/X _14618_/A vssd1 vssd1 vccd1 vccd1 _18267_/D
+ sky130_fd_sc_hd__a22o_1
X_11837_ _15867_/A _15839_/A vssd1 vssd1 vccd1 vccd1 _12183_/B sky130_fd_sc_hd__or2_2
XFILLER_33_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18393_ _18441_/CLK _18393_/D vssd1 vssd1 vccd1 vccd1 _18393_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_199_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17003__S _17547_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14556_ _18306_/Q _14547_/A _14474_/X _14548_/A vssd1 vssd1 vccd1 vccd1 _18306_/D
+ sky130_fd_sc_hd__a22o_1
X_17344_ _16346_/Y _17854_/X _17568_/S vssd1 vssd1 vccd1 vccd1 _17344_/X sky130_fd_sc_hd__mux2_1
XFILLER_202_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11768_ hold186/X _11764_/X _19478_/Q _11765_/X vssd1 vssd1 vccd1 vccd1 hold188/A
+ sky130_fd_sc_hd__o22a_1
XPHY_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10719_ _15971_/A _13252_/D vssd1 vssd1 vccd1 vccd1 _10721_/A sky130_fd_sc_hd__or2_2
XPHY_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13507_ _18764_/Q vssd1 vssd1 vccd1 vccd1 _14695_/A sky130_fd_sc_hd__inv_2
XANTENNA__16842__S _17546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17275_ _17274_/X _11435_/Y _17548_/S vssd1 vssd1 vccd1 vccd1 _17275_/X sky130_fd_sc_hd__mux2_1
X_14487_ _18347_/Q _14479_/A _12731_/X _14480_/A vssd1 vssd1 vccd1 vccd1 _18347_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14708__B2 _14701_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11699_ _19522_/Q _11691_/A _10868_/X _11692_/A vssd1 vssd1 vccd1 vccd1 _19522_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_228_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19014_ _19115_/CLK _19014_/D hold353/X vssd1 vssd1 vccd1 vccd1 _19014_/Q sky130_fd_sc_hd__dfrtp_4
X_13438_ _13350_/A _13350_/B _13437_/X _13352_/C vssd1 vssd1 vccd1 vccd1 _18863_/D
+ sky130_fd_sc_hd__a211oi_4
X_16226_ _19769_/Q vssd1 vssd1 vccd1 vccd1 _16226_/Y sky130_fd_sc_hd__inv_2
Xrebuffer1 rebuffer1/A vssd1 vssd1 vccd1 vccd1 _12985_/A sky130_fd_sc_hd__dlygate4sd1_1
XANTENNA__13392__B1 _20113_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08938__A2 _08937_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16157_ _18070_/Q vssd1 vssd1 vccd1 vccd1 _16157_/Y sky130_fd_sc_hd__inv_2
X_13369_ _20107_/Q vssd1 vssd1 vccd1 vccd1 _13369_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15108_ _18526_/D _11173_/C _18527_/D _17985_/Q _15107_/X vssd1 vssd1 vccd1 vccd1
+ _17985_/D sky130_fd_sc_hd__a32o_1
X_16088_ _18149_/Q vssd1 vssd1 vccd1 vccd1 _16088_/Y sky130_fd_sc_hd__inv_2
XFILLER_170_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17673__S _17683_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19916_ _19937_/CLK _19916_/D repeater189/X vssd1 vssd1 vccd1 vccd1 _19916_/Q sky130_fd_sc_hd__dfrtp_1
X_15039_ _18032_/Q _15035_/X _14996_/X _15037_/X vssd1 vssd1 vccd1 vccd1 _18032_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_102_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19847_ _19847_/CLK _19847_/D repeater264/X vssd1 vssd1 vccd1 vccd1 _19847_/Q sky130_fd_sc_hd__dfrtp_1
X_09600_ _09476_/A _09600_/A2 _09598_/Y _09587_/X vssd1 vssd1 vccd1 vccd1 _20016_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_84_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19778_ _19780_/CLK _19778_/D repeater218/X vssd1 vssd1 vccd1 vccd1 _19778_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_243_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09531_ _19309_/Q vssd1 vssd1 vccd1 vccd1 _09531_/Y sky130_fd_sc_hd__inv_2
X_18729_ _19224_/CLK _18729_/D repeater253/X vssd1 vssd1 vccd1 vccd1 _18729_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17808__S1 _18750_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_243_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_236_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09462_ _10035_/A _19379_/Q _19919_/Q _09458_/Y _09461_/X vssd1 vssd1 vccd1 vccd1
+ _09463_/D sky130_fd_sc_hd__o221a_1
XFILLER_25_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16397__B1 _15859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_212_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09393_ _10101_/C _19367_/Q _10011_/A _19369_/Q _09392_/X vssd1 vssd1 vccd1 vccd1
+ _09394_/D sky130_fd_sc_hd__o221a_1
XFILLER_178_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11750__A _11771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18964__RESET_B hold370/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16149__B1 _17417_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19504__CLK _19510_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16053__A _16053_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17583__S _17584_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19752__RESET_B repeater196/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11697__B1 _10863_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_235_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_228_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09729_ _09729_/A vssd1 vssd1 vccd1 vccd1 _09848_/B sky130_fd_sc_hd__inv_2
XANTENNA__16927__S _16950_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_243_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12740_ _18822_/Q vssd1 vssd1 vccd1 vccd1 _13545_/A sky130_fd_sc_hd__inv_2
XFILLER_216_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12671_ _12678_/A vssd1 vssd1 vccd1 vccd1 _12671_/X sky130_fd_sc_hd__buf_1
XPHY_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14410_ _14410_/A vssd1 vssd1 vccd1 vccd1 _14411_/A sky130_fd_sc_hd__inv_2
XPHY_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11622_ _11622_/A _11622_/B vssd1 vssd1 vccd1 vccd1 _11632_/A sky130_fd_sc_hd__or2_1
XPHY_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15390_ _19523_/Q vssd1 vssd1 vccd1 vccd1 _15390_/Y sky130_fd_sc_hd__inv_2
XPHY_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20011__CLK _20013_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14341_ _18431_/Q _14336_/X _14279_/X _14338_/X vssd1 vssd1 vccd1 vccd1 _18431_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11553_ _19560_/Q vssd1 vssd1 vccd1 vccd1 _11573_/A sky130_fd_sc_hd__inv_2
XPHY_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10504_ _19545_/Q _19540_/Q _19539_/Q _11654_/A vssd1 vssd1 vccd1 vccd1 _10505_/C
+ sky130_fd_sc_hd__or4_4
X_17060_ _17059_/X _18828_/Q _17386_/S vssd1 vssd1 vccd1 vccd1 _17060_/X sky130_fd_sc_hd__mux2_2
XPHY_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14272_ _14274_/A vssd1 vssd1 vccd1 vccd1 _14272_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_183_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11484_ _11484_/A _11484_/B vssd1 vssd1 vccd1 vccd1 _11497_/A sky130_fd_sc_hd__or2_1
XFILLER_137_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16011_ _17988_/Q vssd1 vssd1 vccd1 vccd1 _16011_/Y sky130_fd_sc_hd__inv_2
X_13223_ _18536_/Q _13223_/B vssd1 vssd1 vccd1 vccd1 _13224_/B sky130_fd_sc_hd__or2_1
XFILLER_171_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10435_ _10452_/A vssd1 vssd1 vccd1 vccd1 _10435_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__10188__A0 _10147_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13154_ _19166_/Q _13068_/A _19183_/Q _13084_/A vssd1 vssd1 vccd1 vccd1 _13154_/X
+ sky130_fd_sc_hd__o22a_1
X_10366_ _10366_/A vssd1 vssd1 vccd1 vccd1 _10367_/B sky130_fd_sc_hd__inv_2
XFILLER_3_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12105_ _19311_/Q _12094_/X _12104_/X _12096_/X vssd1 vssd1 vccd1 vccd1 _19311_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17493__S _17493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13085_ _13085_/A _13085_/B vssd1 vssd1 vccd1 vccd1 _13169_/A sky130_fd_sc_hd__or2_1
X_17962_ _20036_/CLK _17962_/D vssd1 vssd1 vccd1 vccd1 _17962_/Q sky130_fd_sc_hd__dfxtp_1
X_10297_ _18592_/Q _15588_/A vssd1 vssd1 vccd1 vccd1 _15593_/A sky130_fd_sc_hd__or2_1
XFILLER_239_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19493__RESET_B repeater260/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19701_ _20055_/CLK _19701_/D repeater202/X vssd1 vssd1 vccd1 vccd1 _19701_/Q sky130_fd_sc_hd__dfstp_1
X_16913_ _16646_/Y _20113_/Q _17385_/S vssd1 vssd1 vccd1 vccd1 _16913_/X sky130_fd_sc_hd__mux2_1
X_12036_ _12044_/A vssd1 vssd1 vccd1 vccd1 _12036_/X sky130_fd_sc_hd__clkbuf_2
X_17893_ _16019_/Y _16020_/Y _16021_/Y _16022_/Y _17913_/S0 _19632_/Q vssd1 vssd1
+ vccd1 vccd1 _17893_/X sky130_fd_sc_hd__mux4_2
XANTENNA__19422__RESET_B repeater271/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16076__C1 _16074_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19632_ _19637_/CLK _19632_/D repeater258/X vssd1 vssd1 vccd1 vccd1 _19632_/Q sky130_fd_sc_hd__dfrtp_2
X_16844_ _16843_/X _11446_/Y _17548_/S vssd1 vssd1 vccd1 vccd1 _16844_/X sky130_fd_sc_hd__mux2_1
XANTENNA__14211__A _19123_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19563_ _19577_/CLK _19563_/D repeater268/X vssd1 vssd1 vccd1 vccd1 _19563_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_92_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16775_ _15963_/X _09517_/Y _17534_/S vssd1 vssd1 vccd1 vccd1 _16775_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12101__A1 _19313_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13987_ _18687_/Q vssd1 vssd1 vccd1 vccd1 _14017_/A sky130_fd_sc_hd__inv_2
XANTENNA__16837__S _17488_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18514_ _20048_/CLK _18514_/D repeater208/X vssd1 vssd1 vccd1 vccd1 _18514_/Q sky130_fd_sc_hd__dfrtp_1
X_15726_ _15726_/A _15727_/B vssd1 vssd1 vccd1 vccd1 _18659_/D sky130_fd_sc_hd__nor2_1
XFILLER_92_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19494_ _19515_/CLK hold141/X repeater260/X vssd1 vssd1 vccd1 vccd1 _19494_/Q sky130_fd_sc_hd__dfrtp_1
X_12938_ _19292_/Q vssd1 vssd1 vccd1 vccd1 _12938_/Y sky130_fd_sc_hd__inv_2
XFILLER_233_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18445_ _19865_/CLK _18445_/D vssd1 vssd1 vccd1 vccd1 _18445_/Q sky130_fd_sc_hd__dfxtp_1
X_15657_ _15657_/A _15657_/B vssd1 vssd1 vccd1 vccd1 _15657_/Y sky130_fd_sc_hd__nor2_1
XPHY_4190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_61_HCLK_A clkbuf_opt_3_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12869_ _18929_/Q vssd1 vssd1 vccd1 vccd1 _13008_/A sky130_fd_sc_hd__inv_2
XANTENNA__15051__B1 _14996_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_221_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14608_ _18278_/Q _14599_/X _14578_/X _14602_/X vssd1 vssd1 vccd1 vccd1 _18278_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13384__A1_N _20115_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18376_ _19637_/CLK _18376_/D vssd1 vssd1 vccd1 vccd1 _18376_/Q sky130_fd_sc_hd__dfxtp_1
X_15588_ _15588_/A vssd1 vssd1 vccd1 vccd1 _15594_/B sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_92_HCLK clkbuf_4_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19976_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_193_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17327_ _15963_/X _12821_/Y _17534_/S vssd1 vssd1 vccd1 vccd1 _17327_/X sky130_fd_sc_hd__mux2_1
XANTENNA__17668__S _17683_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14539_ _18318_/Q _14530_/X _14509_/X _14533_/X vssd1 vssd1 vccd1 vccd1 _18318_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_239_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17258_ _17257_/X _19210_/Q _17545_/S vssd1 vssd1 vccd1 vccd1 _17258_/X sky130_fd_sc_hd__mux2_1
XANTENNA__18551__CLK _19780_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16209_ _16209_/A _16212_/B vssd1 vssd1 vccd1 vccd1 _16209_/Y sky130_fd_sc_hd__nor2_1
X_17189_ _17188_/X _14069_/Y _17544_/S vssd1 vssd1 vccd1 vccd1 _17189_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10179__B1 _09105_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08962_ _18780_/Q vssd1 vssd1 vccd1 vccd1 _08962_/Y sky130_fd_sc_hd__inv_2
XFILLER_229_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_217_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20068__RESET_B repeater207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_225_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09514_ _19307_/Q vssd1 vssd1 vccd1 vccd1 _09514_/Y sky130_fd_sc_hd__inv_2
XFILLER_140_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_213_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_197_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09445_ _10034_/A _19378_/Q _19918_/Q _09442_/Y _09444_/X vssd1 vssd1 vccd1 vccd1
+ _09463_/A sky130_fd_sc_hd__o221a_1
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15042__B1 _15002_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09376_ _19928_/Q vssd1 vssd1 vccd1 vccd1 _10044_/A sky130_fd_sc_hd__inv_2
XFILLER_197_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17578__S _17584_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14791__A _14791_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10709__A2 _10704_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10220_ _19665_/Q vssd1 vssd1 vccd1 vccd1 _10965_/A sky130_fd_sc_hd__inv_2
XFILLER_79_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10151_ _10186_/A _10186_/B _15961_/A vssd1 vssd1 vccd1 vccd1 _10152_/S sky130_fd_sc_hd__or3_1
XFILLER_134_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10082_ _10082_/A _10099_/A vssd1 vssd1 vccd1 vccd1 _10097_/A sky130_fd_sc_hd__or2_2
XFILLER_121_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_247_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13910_ _13910_/A _13910_/B _13910_/C _13910_/D vssd1 vssd1 vccd1 vccd1 _13911_/D
+ sky130_fd_sc_hd__or4_4
XFILLER_87_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_247_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14890_ _18117_/Q _14883_/X _14812_/X _14885_/X vssd1 vssd1 vccd1 vccd1 _18117_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_102_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_207_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13841_ _13840_/Y _13832_/A _19223_/Q _18734_/Q vssd1 vssd1 vccd1 vccd1 _13843_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_207_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16560_ _19454_/Q vssd1 vssd1 vccd1 vccd1 _16560_/Y sky130_fd_sc_hd__inv_2
X_13772_ _18739_/Q _18740_/Q _13772_/S vssd1 vssd1 vccd1 vccd1 _18740_/D sky130_fd_sc_hd__mux2_1
XFILLER_28_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10984_ _19664_/Q _10984_/B vssd1 vssd1 vccd1 vccd1 _10984_/Y sky130_fd_sc_hd__nor2_1
XFILLER_74_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18815__RESET_B repeater239/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15511_ _15511_/A _15511_/B vssd1 vssd1 vccd1 vccd1 _15511_/Y sky130_fd_sc_hd__nor2_1
XFILLER_243_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12723_ _14810_/A vssd1 vssd1 vccd1 vccd1 _12723_/X sky130_fd_sc_hd__clkbuf_2
X_16491_ _16489_/Y _15884_/A _16490_/Y _15915_/A vssd1 vssd1 vccd1 vccd1 _16492_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__15033__B1 _15020_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18230_ _18412_/CLK _18230_/D vssd1 vssd1 vccd1 vccd1 _18230_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15442_ _15259_/Y _15257_/Y _15439_/A vssd1 vssd1 vccd1 vccd1 _18548_/D sky130_fd_sc_hd__o21a_1
XFILLER_188_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12654_ _18996_/Q _12650_/X _12533_/X _12651_/X vssd1 vssd1 vccd1 vccd1 _18996_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_231_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11605_ _11579_/A _11579_/B _11569_/A _11603_/Y vssd1 vssd1 vccd1 vccd1 _19566_/D
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__17488__S _17488_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09799__C1 _09813_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18161_ _18216_/CLK _18161_/D vssd1 vssd1 vccd1 vccd1 _18161_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15373_ _19789_/Q _10649_/B _10650_/B vssd1 vssd1 vccd1 vccd1 _15373_/X sky130_fd_sc_hd__a21bo_1
X_12585_ _19041_/Q _12583_/X _12413_/X _12584_/X vssd1 vssd1 vccd1 vccd1 _19041_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17112_ _17473_/A0 _16535_/Y _17547_/S vssd1 vssd1 vccd1 vccd1 _17112_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14324_ hold325/X vssd1 vssd1 vccd1 vccd1 hold324/A sky130_fd_sc_hd__clkbuf_2
XPHY_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11536_ _19583_/Q _11535_/Y _11521_/X _11465_/B vssd1 vssd1 vccd1 vccd1 _19583_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_129_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18092_ _18765_/CLK _18092_/D vssd1 vssd1 vccd1 vccd1 _18092_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_183_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14255_ _14255_/A vssd1 vssd1 vccd1 vccd1 _15318_/B sky130_fd_sc_hd__buf_1
X_17043_ _17042_/X _15541_/Y _17474_/S vssd1 vssd1 vccd1 vccd1 _17043_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_repeater230_A repeater233/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11467_ _11467_/A _11467_/B vssd1 vssd1 vccd1 vccd1 _11468_/C sky130_fd_sc_hd__or2_2
XFILLER_99_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13206_ _13066_/A _13206_/A2 _13204_/Y _13202_/X vssd1 vssd1 vccd1 vccd1 _18893_/D
+ sky130_fd_sc_hd__a211oi_2
X_10418_ _12232_/A vssd1 vssd1 vccd1 vccd1 _10418_/X sky130_fd_sc_hd__buf_4
X_14186_ _19124_/Q _18703_/Q _14185_/Y _14034_/Y vssd1 vssd1 vccd1 vccd1 _14193_/A
+ sky130_fd_sc_hd__o22a_1
X_11398_ _19570_/Q _19150_/Q _19570_/Q _19150_/Q vssd1 vssd1 vccd1 vccd1 _11398_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_152_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13137_ _19169_/Q vssd1 vssd1 vccd1 vccd1 _13137_/Y sky130_fd_sc_hd__inv_2
XFILLER_225_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10349_ _19863_/Q _10349_/B vssd1 vssd1 vccd1 vccd1 _10349_/Y sky130_fd_sc_hd__nor2_1
X_18994_ _19208_/CLK _18994_/D repeater249/X vssd1 vssd1 vccd1 vccd1 _18994_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__15963__C _17548_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_239_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13068_ _13068_/A _13068_/B vssd1 vssd1 vccd1 vccd1 _13069_/C sky130_fd_sc_hd__or2_2
X_17945_ _18260_/CLK _17945_/D vssd1 vssd1 vccd1 vccd1 _17945_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrepeater205 repeater207/X vssd1 vssd1 vccd1 vccd1 repeater205/X sky130_fd_sc_hd__clkbuf_8
XFILLER_239_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12019_ _19351_/Q _12016_/X hold300/X _12017_/X vssd1 vssd1 vccd1 vccd1 _19351_/D
+ sky130_fd_sc_hd__a22o_1
Xrepeater216 repeater242/X vssd1 vssd1 vccd1 vccd1 repeater216/X sky130_fd_sc_hd__clkbuf_8
Xrepeater227 repeater228/X vssd1 vssd1 vccd1 vccd1 repeater227/X sky130_fd_sc_hd__buf_6
Xrepeater238 repeater239/X vssd1 vssd1 vccd1 vccd1 repeater238/X sky130_fd_sc_hd__buf_6
X_17876_ _16101_/Y _16102_/Y _16103_/Y _16104_/Y _17908_/S0 _18759_/Q vssd1 vssd1
+ vccd1 vccd1 _17876_/X sky130_fd_sc_hd__mux4_2
XFILLER_241_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xrepeater249 hold370/X vssd1 vssd1 vccd1 vccd1 repeater249/X sky130_fd_sc_hd__clkbuf_8
XFILLER_227_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19615_ _19937_/CLK _19615_/D repeater190/X vssd1 vssd1 vccd1 vccd1 _19615_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__09035__A hold306/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16827_ _16826_/X _09874_/A _17524_/S vssd1 vssd1 vccd1 vccd1 _16827_/X sky130_fd_sc_hd__mux2_2
XFILLER_38_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19546_ _19595_/CLK _19546_/D hold346/A vssd1 vssd1 vccd1 vccd1 _19546_/Q sky130_fd_sc_hd__dfrtp_1
X_16758_ vssd1 vssd1 vccd1 vccd1 _16758_/HI _16758_/LO sky130_fd_sc_hd__conb_1
XFILLER_0_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_234_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18556__RESET_B repeater193/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15709_ _15709_/A _15713_/B vssd1 vssd1 vccd1 vccd1 _18644_/D sky130_fd_sc_hd__nor2_1
X_19477_ _19506_/CLK hold192/X repeater256/X vssd1 vssd1 vccd1 vccd1 _19477_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12396__A hold296/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16689_ _17054_/X _16637_/X _17037_/X _16638_/X vssd1 vssd1 vccd1 vccd1 _16689_/X
+ sky130_fd_sc_hd__o22a_1
X_09230_ _18644_/Q _09226_/X _18644_/Q _09226_/X vssd1 vssd1 vccd1 vccd1 _09231_/A
+ sky130_fd_sc_hd__o2bb2a_1
X_18428_ _18795_/CLK _18428_/D vssd1 vssd1 vccd1 vccd1 _18428_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16772__A0 _15963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09161_ _20081_/Q vssd1 vssd1 vccd1 vccd1 _14699_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__17398__S _17567_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18359_ _19849_/CLK _18359_/D vssd1 vssd1 vccd1 vccd1 _18359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_187_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_175_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09092_ hold326/X vssd1 vssd1 vccd1 vccd1 _14791_/A sky130_fd_sc_hd__buf_4
XFILLER_119_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_175_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19344__RESET_B repeater244/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09994_ _09854_/A _09854_/B _09992_/Y _09990_/X vssd1 vssd1 vccd1 vccd1 _19945_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_131_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08945_ _18772_/Q vssd1 vssd1 vccd1 vccd1 _08945_/Y sky130_fd_sc_hd__inv_2
XFILLER_229_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16460__C1 _16459_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12077__B1 _12076_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_232_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11824__B1 _10885_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15015__B1 _14998_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09428_ _10015_/C _19377_/Q _19917_/Q _09424_/Y _09427_/X vssd1 vssd1 vccd1 vccd1
+ _09440_/B sky130_fd_sc_hd__o221a_1
XANTENNA__16763__A0 _15963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_hold323_A HWDATA[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09359_ _20018_/Q vssd1 vssd1 vccd1 vccd1 _09478_/A sky130_fd_sc_hd__inv_2
XFILLER_12_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16506__A _16506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17101__S _17530_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12370_ _12370_/A _12370_/B _12370_/C vssd1 vssd1 vccd1 vccd1 _15902_/A sky130_fd_sc_hd__or3_4
XFILLER_165_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19992__CLK _19992_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_219_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11321_ _18971_/Q vssd1 vssd1 vccd1 vccd1 _11321_/Y sky130_fd_sc_hd__inv_2
XFILLER_166_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16940__S _16946_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14040_ _14039_/Y _18691_/Q _19075_/Q _14016_/A vssd1 vssd1 vccd1 vccd1 _14040_/X
+ sky130_fd_sc_hd__a22o_1
X_11252_ _19590_/Q vssd1 vssd1 vccd1 vccd1 _11470_/A sky130_fd_sc_hd__inv_2
X_10203_ _19831_/Q vssd1 vssd1 vccd1 vccd1 _10203_/Y sky130_fd_sc_hd__inv_2
XFILLER_134_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11183_ _17709_/X _11176_/X _19622_/Q _11178_/X vssd1 vssd1 vccd1 vccd1 _19622_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11088__C _12053_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14829__B1 _14780_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10134_ _10133_/A _10132_/B _13283_/C _10133_/X _09197_/B vssd1 vssd1 vccd1 vccd1
+ _10136_/A sky130_fd_sc_hd__a2111o_4
X_15991_ _17496_/X vssd1 vssd1 vccd1 vccd1 _15991_/Y sky130_fd_sc_hd__inv_2
XFILLER_192_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17730_ _15379_/X _19715_/Q _18508_/D vssd1 vssd1 vccd1 vccd1 _17730_/X sky130_fd_sc_hd__mux2_1
X_10065_ _10065_/A vssd1 vssd1 vccd1 vccd1 _10065_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14942_ _18089_/Q _14939_/X _14921_/X _14941_/X vssd1 vssd1 vccd1 vccd1 _18089_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_209_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17661_ _15591_/X _19028_/Q _17664_/S vssd1 vssd1 vccd1 vccd1 _18591_/D sky130_fd_sc_hd__mux2_1
XFILLER_75_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14873_ _14873_/A vssd1 vssd1 vccd1 vccd1 _14873_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_output128_A _19749_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19400_ _19905_/CLK _19400_/D repeater191/X vssd1 vssd1 vccd1 vccd1 _19400_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_62_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16612_ _16866_/X _15889_/X _17006_/X _15887_/X vssd1 vssd1 vccd1 vccd1 _16612_/X
+ sky130_fd_sc_hd__o22a_2
X_13824_ _13909_/A _13929_/A vssd1 vssd1 vccd1 vccd1 _13825_/B sky130_fd_sc_hd__or2_2
X_17592_ _15353_/X _19711_/Q _17600_/S vssd1 vssd1 vccd1 vccd1 _17592_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19331_ _19956_/CLK _19331_/D hold371/X vssd1 vssd1 vccd1 vccd1 _19331_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_189_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16543_ _16543_/A _16544_/B vssd1 vssd1 vccd1 vccd1 _16543_/Y sky130_fd_sc_hd__nor2_1
XFILLER_204_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_repeater180_A _17530_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10967_ _10967_/A _10973_/A vssd1 vssd1 vccd1 vccd1 _10968_/A sky130_fd_sc_hd__or2_1
X_13755_ _13745_/Y _17763_/S _18747_/Q _13287_/X vssd1 vssd1 vccd1 vccd1 _13756_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_189_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12706_ _18960_/Q _12677_/A _12543_/X _12678_/A vssd1 vssd1 vccd1 vccd1 _18960_/D
+ sky130_fd_sc_hd__a22o_1
X_19262_ _19283_/CLK _19262_/D repeater212/X vssd1 vssd1 vccd1 vccd1 _19262_/Q sky130_fd_sc_hd__dfrtp_1
X_16474_ _19033_/Q _17473_/S vssd1 vssd1 vccd1 vccd1 _16474_/Y sky130_fd_sc_hd__nand2_1
X_10898_ _19690_/Q _10893_/X _10885_/X _10895_/X vssd1 vssd1 vccd1 vccd1 _19690_/D
+ sky130_fd_sc_hd__a22o_1
X_13686_ _13686_/A vssd1 vssd1 vccd1 vccd1 _13686_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13568__B1 _13597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18213_ _18216_/CLK _18213_/D vssd1 vssd1 vccd1 vccd1 _18213_/Q sky130_fd_sc_hd__dfxtp_1
X_15425_ _19616_/Q _11161_/B _11162_/B vssd1 vssd1 vccd1 vccd1 _15425_/X sky130_fd_sc_hd__a21bo_1
XPHY_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12637_ _12651_/A vssd1 vssd1 vccd1 vccd1 _12637_/X sky130_fd_sc_hd__clkbuf_2
X_19193_ _19221_/CLK _19193_/D hold367/X vssd1 vssd1 vccd1 vccd1 _19193_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17011__S _17548_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18144_ _18169_/CLK _18144_/D vssd1 vssd1 vccd1 vccd1 _18144_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15356_ _15358_/A _17591_/X vssd1 vssd1 vccd1 vccd1 _18499_/D sky130_fd_sc_hd__and2_1
XFILLER_145_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12568_ _19052_/Q _12560_/X _12386_/X _12563_/X vssd1 vssd1 vccd1 vccd1 _19052_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11519_ _11472_/A _11519_/A2 _11506_/X _11517_/Y vssd1 vssd1 vccd1 vccd1 _19592_/D
+ sky130_fd_sc_hd__a211oi_2
X_14307_ _18448_/Q _14303_/X _14277_/X _14305_/X vssd1 vssd1 vccd1 vccd1 _18448_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_117_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18075_ _18260_/CLK _18075_/D vssd1 vssd1 vccd1 vccd1 _18075_/Q sky130_fd_sc_hd__dfxtp_1
X_15287_ _15439_/A _15443_/B _15287_/C vssd1 vssd1 vccd1 vccd1 _18629_/D sky130_fd_sc_hd__nand3_1
X_12499_ _12506_/A vssd1 vssd1 vccd1 vccd1 _12499_/X sky130_fd_sc_hd__buf_1
XANTENNA__16850__S _17545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold207 HADDR[3] vssd1 vssd1 vccd1 vccd1 input26/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold218 hold218/A vssd1 vssd1 vccd1 vccd1 hold218/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09539__A2 _19319_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold229 hold229/A vssd1 vssd1 vccd1 vccd1 hold229/X sky130_fd_sc_hd__dlygate4sd3_1
X_17026_ _17025_/X _20012_/Q _17414_/S vssd1 vssd1 vccd1 vccd1 _17026_/X sky130_fd_sc_hd__mux2_2
X_14238_ _18669_/Q _14236_/X _18668_/Q _17600_/S vssd1 vssd1 vccd1 vccd1 _18669_/D
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_122_HCLK clkbuf_4_4_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19597_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_113_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10003__C1 _09964_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14169_ _14167_/Y _18693_/Q _14168_/Y _18675_/Q vssd1 vssd1 vccd1 vccd1 _14169_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_124_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18977_ _19600_/CLK _18977_/D hold273/X vssd1 vssd1 vccd1 vccd1 _18977_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__11295__A _19021_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17681__S _17683_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17928_ _19437_/CLK _19437_/Q vssd1 vssd1 vccd1 vccd1 _17928_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_239_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_226_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17859_ _17855_/X _17856_/X _17857_/X _17858_/X _18760_/Q _18761_/Q vssd1 vssd1 vccd1
+ vccd1 _17859_/X sky130_fd_sc_hd__mux4_2
XFILLER_242_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16993__A0 _15768_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_242_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19529_ _19544_/CLK _19529_/D repeater221/X vssd1 vssd1 vccd1 vccd1 _19529_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_235_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11806__B1 _09051_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09213_ _09213_/A vssd1 vssd1 vccd1 vccd1 _09214_/B sky130_fd_sc_hd__inv_2
XFILLER_22_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_210_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09144_ _09154_/A _09149_/A _09144_/C _20085_/Q vssd1 vssd1 vccd1 vccd1 _15322_/C
+ sky130_fd_sc_hd__or4_4
XFILLER_182_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12231__B1 _11981_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17170__A0 _15963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09075_ hold250/X vssd1 vssd1 vccd1 vccd1 _09075_/X sky130_fd_sc_hd__buf_4
XFILLER_146_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20083__RESET_B repeater204/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09977_ _09863_/A _09863_/B _09975_/Y _09970_/X vssd1 vssd1 vccd1 vccd1 _19955_/D
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__10821__B _10841_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17591__S _17600_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08928_ _18787_/Q vssd1 vssd1 vccd1 vccd1 _08928_/Y sky130_fd_sc_hd__inv_2
X_20097_ _20107_/CLK _20097_/D repeater233/X vssd1 vssd1 vccd1 vccd1 _20097_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_85_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15405__A _15413_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11933__A _11933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11870_ _19433_/Q _11869_/Y _11867_/X vssd1 vssd1 vccd1 vccd1 _19433_/D sky130_fd_sc_hd__o21a_1
XANTENNA__17987__CLK _19851_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10821_ _15854_/A _10841_/A vssd1 vssd1 vccd1 vccd1 _10831_/B sky130_fd_sc_hd__or2_4
XFILLER_232_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16935__S _16946_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10752_ _18631_/Q vssd1 vssd1 vccd1 vccd1 _15436_/A sky130_fd_sc_hd__clkbuf_2
X_13540_ _13540_/A _13590_/A vssd1 vssd1 vccd1 vccd1 _13541_/B sky130_fd_sc_hd__or2_2
XFILLER_41_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12470__B1 hold270/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13471_ _18848_/Q _13470_/Y _13443_/A _13336_/B vssd1 vssd1 vccd1 vccd1 _18848_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_201_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10683_ _17744_/X _10676_/A _19781_/Q _10677_/A vssd1 vssd1 vccd1 vccd1 _19781_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_139_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_197_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16236__A _16633_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_200_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15210_ _19682_/Q _19681_/Q _19683_/Q vssd1 vssd1 vccd1 vccd1 _15216_/C sky130_fd_sc_hd__or3_4
X_12422_ _19137_/Q _12420_/X _12353_/X _12421_/X vssd1 vssd1 vccd1 vccd1 _19137_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12222__B1 _12038_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16190_ _10625_/Y _15277_/Y _16189_/X vssd1 vssd1 vccd1 vccd1 _18552_/D sky130_fd_sc_hd__o21ai_1
XFILLER_127_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_145_HCLK clkbuf_4_1_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19668_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__19266__RESET_B repeater212/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12353_ hold240/X vssd1 vssd1 vccd1 vccd1 _12353_/X sky130_fd_sc_hd__clkbuf_4
X_15141_ _17964_/Q _15134_/X _10715_/X _15136_/X vssd1 vssd1 vccd1 vccd1 _17964_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_181_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11304_ _18978_/Q vssd1 vssd1 vccd1 vccd1 _11304_/Y sky130_fd_sc_hd__inv_2
X_15072_ _15072_/A vssd1 vssd1 vccd1 vccd1 _15073_/A sky130_fd_sc_hd__inv_2
XANTENNA__19738__CLK _20051_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12284_ _12300_/A vssd1 vssd1 vccd1 vccd1 _12284_/X sky130_fd_sc_hd__clkbuf_2
X_14023_ _14023_/A _14115_/A vssd1 vssd1 vccd1 vccd1 _14024_/B sky130_fd_sc_hd__or2_2
X_18900_ _19352_/CLK _18900_/D hold373/X vssd1 vssd1 vccd1 vccd1 _18900_/Q sky130_fd_sc_hd__dfrtp_1
X_11235_ _19593_/Q _11230_/Y _11487_/A _19021_/Q _11234_/X vssd1 vssd1 vccd1 vccd1
+ _11248_/B sky130_fd_sc_hd__o221a_1
XFILLER_106_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19880_ _20059_/CLK _19880_/D repeater200/X vssd1 vssd1 vccd1 vccd1 _19880_/Q sky130_fd_sc_hd__dfrtp_1
X_18831_ _19255_/CLK _18831_/D repeater237/X vssd1 vssd1 vccd1 vccd1 _18831_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_96_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11166_ _19621_/Q _11166_/B vssd1 vssd1 vccd1 vccd1 _11167_/B sky130_fd_sc_hd__or2_1
XFILLER_49_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18762__CLK _20123_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10117_ _18565_/Q _18564_/Q _15474_/A vssd1 vssd1 vccd1 vccd1 _15481_/A sky130_fd_sc_hd__or3_1
XANTENNA__12289__B1 _12032_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18762_ _20123_/CLK _18762_/D repeater195/X vssd1 vssd1 vccd1 vccd1 _18762_/Q sky130_fd_sc_hd__dfrtp_1
X_15974_ _18479_/Q vssd1 vssd1 vccd1 vccd1 _15974_/Y sky130_fd_sc_hd__inv_2
X_11097_ _15094_/B vssd1 vssd1 vccd1 vccd1 _14963_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_48_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17713_ _15427_/X _19528_/Q _18546_/D vssd1 vssd1 vccd1 vccd1 _17713_/X sky130_fd_sc_hd__mux2_1
XANTENNA__18830__RESET_B repeater239/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10048_ _10048_/A _10055_/A vssd1 vssd1 vccd1 vccd1 _10049_/A sky130_fd_sc_hd__or2_2
X_14925_ _20080_/Q vssd1 vssd1 vccd1 vccd1 _14925_/X sky130_fd_sc_hd__clkbuf_2
X_18693_ _18701_/CLK _18693_/D hold359/X vssd1 vssd1 vccd1 vccd1 _18693_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_236_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17006__S _17513_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17644_ _15663_/Y _19045_/Q _17655_/S vssd1 vssd1 vccd1 vccd1 _18608_/D sky130_fd_sc_hd__mux2_1
X_14856_ _18764_/Q vssd1 vssd1 vccd1 vccd1 _15109_/B sky130_fd_sc_hd__buf_1
XFILLER_224_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13807_ _13948_/A _13947_/A _13946_/A _13964_/B vssd1 vssd1 vccd1 vccd1 _13813_/C
+ sky130_fd_sc_hd__or4_4
X_17575_ _15410_/X _19768_/Q _17584_/S vssd1 vssd1 vccd1 vccd1 _17575_/X sky130_fd_sc_hd__mux2_1
XFILLER_51_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14787_ _14787_/A vssd1 vssd1 vccd1 vccd1 _14787_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__16845__S _17543_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11999_ _12043_/A vssd1 vssd1 vccd1 vccd1 _12016_/A sky130_fd_sc_hd__buf_2
X_19314_ _19314_/CLK _19314_/D repeater214/X vssd1 vssd1 vccd1 vccd1 _19314_/Q sky130_fd_sc_hd__dfrtp_4
X_16526_ _19037_/Q vssd1 vssd1 vccd1 vccd1 _16526_/Y sky130_fd_sc_hd__inv_2
XFILLER_232_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12461__B1 _12406_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13738_ _13738_/A vssd1 vssd1 vccd1 vccd1 _13741_/A sky130_fd_sc_hd__inv_2
XANTENNA__16727__B1 _16829_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_220_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19245_ _19320_/CLK _19245_/D repeater214/X vssd1 vssd1 vccd1 vccd1 _19245_/Q sky130_fd_sc_hd__dfrtp_4
X_16457_ _15268_/A _15840_/X _16451_/X _16456_/X vssd1 vssd1 vccd1 vccd1 _16457_/X
+ sky130_fd_sc_hd__o211a_1
X_13669_ _18779_/Q _13664_/X _12596_/X _13665_/X vssd1 vssd1 vccd1 vccd1 _18779_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_31_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15408_ _18536_/Q _13223_/B _13224_/B vssd1 vssd1 vccd1 vccd1 _15408_/X sky130_fd_sc_hd__a21bo_1
X_19176_ _19288_/CLK _19176_/D repeater212/X vssd1 vssd1 vccd1 vccd1 _19176_/Q sky130_fd_sc_hd__dfrtp_1
X_16388_ _16380_/Y _15828_/X _16383_/X _16387_/X vssd1 vssd1 vccd1 vccd1 _16388_/X
+ sky130_fd_sc_hd__o211a_2
XANTENNA__12764__A1 _19229_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18127_ _20090_/CLK _18127_/D vssd1 vssd1 vccd1 vccd1 _18127_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_116_HCLK_A clkbuf_opt_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17676__S _17683_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15339_ _15347_/A _17599_/X vssd1 vssd1 vccd1 vccd1 _18491_/D sky130_fd_sc_hd__and2_1
XFILLER_8_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10775__B1 _19749_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18058_ _18460_/CLK _18058_/D vssd1 vssd1 vccd1 vccd1 _18058_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17009_ _15768_/Y _11286_/Y _17546_/S vssd1 vssd1 vccd1 vccd1 _17009_/X sky130_fd_sc_hd__mux2_1
X_09900_ _19361_/Q vssd1 vssd1 vccd1 vccd1 _09900_/Y sky130_fd_sc_hd__inv_2
XFILLER_99_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20020_ _20091_/CLK _20020_/D repeater240/X vssd1 vssd1 vccd1 vccd1 _20020_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18918__RESET_B repeater188/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09831_ _19955_/Q vssd1 vssd1 vccd1 vccd1 _09863_/A sky130_fd_sc_hd__inv_2
XANTENNA__16663__C1 _16662_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09762_ _19999_/Q _09761_/Y _09629_/B _09761_/A _09759_/X vssd1 vssd1 vccd1 vccd1
+ _19999_/D sky130_fd_sc_hd__o221a_1
XANTENNA__12819__A2 _13529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_227_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_239_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_26_HCLK clkbuf_4_9_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20070_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_55_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09693_ _09746_/A _19419_/Q _19990_/Q _09690_/Y _09692_/X vssd1 vssd1 vccd1 vccd1
+ _09693_/X sky130_fd_sc_hd__a221o_1
XFILLER_66_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrebuffer11 _13085_/B vssd1 vssd1 vccd1 vccd1 _13173_/C1 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_215_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18500__RESET_B repeater219/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrebuffer22 _14012_/C vssd1 vssd1 vccd1 vccd1 _14137_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_4019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer33 _11543_/A vssd1 vssd1 vccd1 vccd1 _11565_/A sky130_fd_sc_hd__buf_2
Xrebuffer44 _11468_/C vssd1 vssd1 vccd1 vccd1 _11527_/A2 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer55 _13081_/B vssd1 vssd1 vccd1 vccd1 _13181_/C1 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrebuffer66 _09488_/B vssd1 vssd1 vccd1 vccd1 _09582_/B1 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_25_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_214_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xrebuffer77 _09875_/B vssd1 vssd1 vccd1 vccd1 _09958_/C1 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer88 _09476_/B vssd1 vssd1 vccd1 vccd1 _09602_/C1 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrebuffer99 _11482_/B vssd1 vssd1 vccd1 vccd1 _11505_/C1 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_242_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12452__B1 _12389_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18635__CLK _19780_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrebuffer101 _09465_/B vssd1 vssd1 vccd1 vccd1 _09620_/A sky130_fd_sc_hd__dlygate4sd1_1
XANTENNA__12204__B1 _12092_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrebuffer112 _13087_/B vssd1 vssd1 vccd1 vccd1 _13170_/C1 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer123 _09857_/C vssd1 vssd1 vccd1 vccd1 _09986_/A2 sky130_fd_sc_hd__dlygate4sd1_1
X_09127_ _09127_/A _09133_/C _15319_/A _09139_/B vssd1 vssd1 vccd1 vccd1 _09127_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_109_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15895__A _15895_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09058_ hold233/X vssd1 vssd1 vccd1 vccd1 _09058_/X sky130_fd_sc_hd__buf_4
XANTENNA__16497__A2 _16148_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12507__A1 _19082_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11928__A _11933_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11020_ _10408_/X _10224_/X _10973_/B _11019_/X vssd1 vssd1 vccd1 vccd1 _19654_/D
+ sky130_fd_sc_hd__o22ai_1
XANTENNA__16249__A2 _16243_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18659__RESET_B repeater210/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_238_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18015__CLK _18169_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12971_ _18947_/Q _12970_/X _12962_/X _12889_/A vssd1 vssd1 vccd1 vccd1 _18947_/D
+ sky130_fd_sc_hd__o211a_1
X_14710_ _18221_/Q _14698_/X _14709_/X _14701_/X vssd1 vssd1 vccd1 vccd1 _18221_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_246_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11922_ _13678_/A vssd1 vssd1 vccd1 vccd1 _11922_/X sky130_fd_sc_hd__buf_2
X_15690_ _18615_/Q vssd1 vssd1 vccd1 vccd1 _15690_/Y sky130_fd_sc_hd__inv_2
XPHY_4520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14641_ _18763_/Q _14641_/B _15195_/B vssd1 vssd1 vccd1 vccd1 _14951_/C sky130_fd_sc_hd__or3_4
XPHY_4553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11853_ _11853_/A vssd1 vssd1 vccd1 vccd1 _13641_/B sky130_fd_sc_hd__inv_2
XPHY_4564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19410__CLK _19984_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10804_ _19733_/Q _10800_/B _10793_/B _10807_/A vssd1 vssd1 vccd1 vccd1 _19733_/D
+ sky130_fd_sc_hd__o211a_1
X_17360_ _17486_/A0 _13131_/Y _17543_/S vssd1 vssd1 vccd1 vccd1 _17360_/X sky130_fd_sc_hd__mux2_1
XPHY_4597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14572_ _14573_/A vssd1 vssd1 vccd1 vccd1 _14572_/X sky130_fd_sc_hd__clkbuf_2
X_11784_ _11800_/A vssd1 vssd1 vccd1 vccd1 _11784_/X sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_3863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16311_ _19761_/Q vssd1 vssd1 vccd1 vccd1 _16311_/Y sky130_fd_sc_hd__inv_2
XPHY_3896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13523_ _13523_/A vssd1 vssd1 vccd1 vccd1 _13523_/Y sky130_fd_sc_hd__inv_2
X_10735_ _10735_/A _10735_/B vssd1 vssd1 vccd1 vccd1 _11650_/B sky130_fd_sc_hd__nand2_1
XFILLER_198_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17291_ _17473_/A0 _16517_/Y _17512_/S vssd1 vssd1 vccd1 vccd1 _17291_/X sky130_fd_sc_hd__mux2_1
XFILLER_40_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19030_ _19667_/CLK _19030_/D repeater264/X vssd1 vssd1 vccd1 vccd1 _19030_/Q sky130_fd_sc_hd__dfrtp_1
X_16242_ _17380_/X _16638_/A _17404_/X _15901_/A _16241_/Y vssd1 vssd1 vccd1 vccd1
+ _16242_/X sky130_fd_sc_hd__o221a_1
X_13454_ _18854_/Q _13453_/Y _13342_/B _13443_/X vssd1 vssd1 vccd1 vccd1 _18854_/D
+ sky130_fd_sc_hd__o211a_1
X_10666_ _17731_/X _10661_/X _19794_/Q _10663_/X vssd1 vssd1 vccd1 vccd1 _19794_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_186_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12405_ _19146_/Q _12400_/X _12404_/X _12402_/X vssd1 vssd1 vccd1 vccd1 _19146_/D
+ sky130_fd_sc_hd__a22o_1
X_13385_ _13383_/Y _18844_/Q _20098_/Q _13467_/A _13384_/X vssd1 vssd1 vccd1 vccd1
+ _13386_/D sky130_fd_sc_hd__o221a_1
X_16173_ _19652_/Q _16095_/Y _16170_/X _16171_/X _16172_/Y vssd1 vssd1 vccd1 vccd1
+ _16173_/X sky130_fd_sc_hd__o221a_1
X_10597_ _10614_/B _10942_/A _15298_/A vssd1 vssd1 vccd1 vccd1 _10598_/A sky130_fd_sc_hd__or3_4
XFILLER_182_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15124_ _15124_/A vssd1 vssd1 vccd1 vccd1 _15124_/X sky130_fd_sc_hd__clkbuf_2
Xoutput109 _16482_/Y vssd1 vssd1 vccd1 vccd1 HRDATA[8] sky130_fd_sc_hd__clkbuf_2
X_12336_ _19179_/Q _12334_/X _12095_/X _12335_/X vssd1 vssd1 vccd1 vccd1 _19179_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_126_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_217_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17780__S1 _19646_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19932_ _19933_/CLK _19932_/D repeater189/X vssd1 vssd1 vccd1 vccd1 _19932_/Q sky130_fd_sc_hd__dfrtp_2
X_15055_ _18020_/Q _15048_/A _15004_/X _15049_/A vssd1 vssd1 vccd1 vccd1 _18020_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_5_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12267_ _19221_/Q _12260_/X _12078_/X _12263_/X vssd1 vssd1 vccd1 vccd1 _19221_/D
+ sky130_fd_sc_hd__a22o_1
X_11218_ _18992_/Q vssd1 vssd1 vccd1 vccd1 _11218_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17437__A1 _11059_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14006_ _14006_/A _14145_/A vssd1 vssd1 vccd1 vccd1 _14007_/B sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_49_HCLK clkbuf_opt_2_HCLK/A vssd1 vssd1 vccd1 vccd1 _19822_/CLK sky130_fd_sc_hd__clkbuf_16
X_19863_ _19865_/CLK _19863_/D repeater267/X vssd1 vssd1 vccd1 vccd1 _19863_/Q sky130_fd_sc_hd__dfrtp_1
X_12198_ _12205_/A vssd1 vssd1 vccd1 vccd1 _12198_/X sky130_fd_sc_hd__buf_1
Xoutput80 _16516_/Y vssd1 vssd1 vccd1 vccd1 HRDATA[10] sky130_fd_sc_hd__clkbuf_2
Xoutput91 _16629_/X vssd1 vssd1 vccd1 vccd1 HRDATA[20] sky130_fd_sc_hd__clkbuf_2
XFILLER_233_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18814_ _19314_/CLK _18814_/D repeater239/X vssd1 vssd1 vccd1 vccd1 _18814_/Q sky130_fd_sc_hd__dfrtp_1
X_11149_ _10263_/X _11148_/X _10263_/X _11148_/X vssd1 vssd1 vccd1 vccd1 _11150_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_19794_ _19794_/CLK _19794_/D repeater219/X vssd1 vssd1 vccd1 vccd1 _19794_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_209_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18745_ _20059_/CLK _18745_/D repeater199/X vssd1 vssd1 vccd1 vccd1 _18745_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18508__CLK _19780_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15957_ _17962_/Q vssd1 vssd1 vccd1 vccd1 _15957_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14908_ _14909_/A vssd1 vssd1 vccd1 vccd1 _14908_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_236_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12682__B1 hold310/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18676_ _18686_/CLK _18676_/D repeater252/X vssd1 vssd1 vccd1 vccd1 _18676_/Q sky130_fd_sc_hd__dfrtp_1
X_15888_ _15888_/A vssd1 vssd1 vccd1 vccd1 _16637_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_236_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17627_ _19892_/Q _19745_/Q _17630_/S vssd1 vssd1 vccd1 vccd1 _17627_/X sky130_fd_sc_hd__mux2_1
X_14839_ _18149_/Q _14832_/X _14812_/X _14834_/X vssd1 vssd1 vccd1 vccd1 _18149_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_224_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19870__RESET_B repeater210/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12434__B1 _12238_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17558_ _17557_/X _19896_/Q _17558_/S vssd1 vssd1 vccd1 vccd1 _17558_/X sky130_fd_sc_hd__mux2_1
XFILLER_211_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19903__CLK _20123_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16509_ _16509_/A vssd1 vssd1 vccd1 vccd1 _16509_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_176_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17489_ _15768_/Y _14171_/Y _17546_/S vssd1 vssd1 vccd1 vccd1 _17489_/X sky130_fd_sc_hd__mux2_1
XFILLER_176_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19228_ _19320_/CLK _19228_/D repeater237/X vssd1 vssd1 vccd1 vccd1 _19228_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_164_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17125__A0 _17473_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19159_ _19214_/CLK _19159_/D repeater188/X vssd1 vssd1 vccd1 vccd1 _19159_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__10748__B1 _10421_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17771__S1 _19646_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18038__CLK _18169_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15151__A2 _15146_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18752__RESET_B repeater195/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16636__C1 _16635_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20003_ _20003_/CLK _20003_/D repeater185/X vssd1 vssd1 vccd1 vccd1 _20003_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_143_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09814_ _09807_/A _09807_/B _19972_/Q _09736_/A _09759_/X vssd1 vssd1 vccd1 vccd1
+ _19972_/D sky130_fd_sc_hd__o221a_1
XFILLER_59_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09745_ _09745_/A _09778_/A vssd1 vssd1 vccd1 vccd1 _09746_/B sky130_fd_sc_hd__or2_2
XFILLER_228_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_243_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_228_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12673__B1 hold308/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09676_ _19412_/Q vssd1 vssd1 vccd1 vccd1 _09676_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11228__B2 _19023_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12425__B1 _12225_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09888__A _19360_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19540__RESET_B repeater221/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_196_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10520_ _19530_/Q vssd1 vssd1 vccd1 vccd1 _10522_/B sky130_fd_sc_hd__inv_2
XFILLER_10_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10451_ _10451_/A vssd1 vssd1 vccd1 vccd1 _10451_/X sky130_fd_sc_hd__buf_4
XANTENNA__10739__A0 _19764_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13170_ _18914_/Q _13169_/Y _13162_/X _13170_/C1 vssd1 vssd1 vccd1 vccd1 _18914_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_201_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10382_ _08921_/X _08964_/X _10321_/C vssd1 vssd1 vccd1 vccd1 _10382_/X sky130_fd_sc_hd__o21a_1
XFILLER_151_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_162_HCLK_A clkbuf_4_0_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12121_ _12121_/A vssd1 vssd1 vccd1 vccd1 _12121_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_190_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_184_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17419__A1 _12937_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12052_ _11848_/Y _11863_/A _11856_/A _13641_/A vssd1 vssd1 vccd1 vccd1 _12052_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_78_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11003_ _10999_/B _11002_/Y _10973_/B _10989_/X _10959_/A vssd1 vssd1 vccd1 vccd1
+ _11004_/A sky130_fd_sc_hd__o32a_1
XFILLER_78_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16860_ _17473_/A0 _16601_/Y _17512_/S vssd1 vssd1 vccd1 vccd1 _16860_/X sky130_fd_sc_hd__mux2_1
XFILLER_77_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09109__B1 _09108_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15811_ _18074_/Q vssd1 vssd1 vccd1 vccd1 _15811_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16791_ _15768_/Y _14185_/Y _17546_/S vssd1 vssd1 vccd1 vccd1 _16791_/X sky130_fd_sc_hd__mux2_1
XFILLER_92_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18530_ _19771_/CLK _18530_/D repeater189/X vssd1 vssd1 vccd1 vccd1 _18530_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_92_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15742_ _18489_/D vssd1 vssd1 vccd1 vccd1 _15747_/C sky130_fd_sc_hd__inv_2
X_12954_ _12951_/Y _18932_/Q _19275_/Q _12964_/D _12953_/X vssd1 vssd1 vccd1 vccd1
+ _12955_/D sky130_fd_sc_hd__o221a_1
XFILLER_246_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18800__CLK _19900_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19628__RESET_B repeater257/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18461_ _19842_/CLK _18461_/D vssd1 vssd1 vccd1 vccd1 _18461_/Q sky130_fd_sc_hd__dfxtp_1
X_11905_ _11914_/A vssd1 vssd1 vccd1 vccd1 _11905_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_output110_A _16499_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15673_ _19437_/Q vssd1 vssd1 vccd1 vccd1 _15673_/X sky130_fd_sc_hd__clkbuf_2
XPHY_4350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12885_ _12885_/A _12885_/B vssd1 vssd1 vccd1 vccd1 _12975_/A sky130_fd_sc_hd__or2_2
XPHY_4361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17412_ _15963_/X _09534_/Y _17534_/S vssd1 vssd1 vccd1 vccd1 _17412_/X sky130_fd_sc_hd__mux2_1
XPHY_4372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14624_ _18268_/Q _14617_/A _09183_/X _14618_/A vssd1 vssd1 vccd1 vccd1 _18268_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18392_ _18441_/CLK _18392_/D vssd1 vssd1 vccd1 vccd1 _18392_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12416__B1 _12344_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11836_ _11996_/A vssd1 vssd1 vccd1 vccd1 _15867_/A sky130_fd_sc_hd__buf_6
XPHY_4394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17343_ _16363_/X _17967_/Q _17564_/S vssd1 vssd1 vccd1 vccd1 _17343_/X sky130_fd_sc_hd__mux2_1
XPHY_3682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_repeater260_A repeater261/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14555_ _18307_/Q _14547_/A hold334/X _14548_/A vssd1 vssd1 vccd1 vccd1 _18307_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11767_ hold180/X _11764_/X _19479_/Q _11765_/X vssd1 vssd1 vccd1 vccd1 hold182/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_13_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13506_ _13506_/A vssd1 vssd1 vccd1 vccd1 _13506_/Y sky130_fd_sc_hd__inv_2
XFILLER_186_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17274_ _17273_/X _11321_/Y _17490_/S vssd1 vssd1 vccd1 vccd1 _17274_/X sky130_fd_sc_hd__mux2_1
X_10718_ _10718_/A vssd1 vssd1 vccd1 vccd1 _13252_/D sky130_fd_sc_hd__buf_2
XANTENNA__15905__B2 _15904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14486_ _18348_/Q _14479_/A _12729_/X _14480_/A vssd1 vssd1 vccd1 vccd1 _18348_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_186_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11698_ _19523_/Q _11691_/A _10866_/X _11692_/A vssd1 vssd1 vccd1 vccd1 _19523_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_146_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19013_ _19597_/CLK _19013_/D repeater281/X vssd1 vssd1 vccd1 vccd1 _19013_/Q sky130_fd_sc_hd__dfrtp_2
X_16225_ _15226_/Y _15840_/X _16218_/Y _15836_/A _16224_/X vssd1 vssd1 vccd1 vccd1
+ _16225_/X sky130_fd_sc_hd__o221a_2
XFILLER_228_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13437_ _13445_/A vssd1 vssd1 vccd1 vccd1 _13437_/X sky130_fd_sc_hd__clkbuf_4
X_10649_ _19789_/Q _10649_/B vssd1 vssd1 vccd1 vccd1 _10650_/B sky130_fd_sc_hd__or2_1
XFILLER_155_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrebuffer2 _12985_/A vssd1 vssd1 vccd1 vccd1 _12960_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__13392__A1 _20111_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19306__CLK _20115_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16156_ _17990_/Q vssd1 vssd1 vccd1 vccd1 _16156_/Y sky130_fd_sc_hd__inv_2
X_13368_ _13365_/Y _18837_/Q _20091_/Q _13327_/A _13367_/X vssd1 vssd1 vccd1 vccd1
+ _13372_/C sky130_fd_sc_hd__o221a_1
XFILLER_115_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15107_ _15762_/B _18526_/Q vssd1 vssd1 vccd1 vccd1 _15107_/X sky130_fd_sc_hd__or2_1
X_12319_ _12361_/A vssd1 vssd1 vccd1 vccd1 _12362_/A sky130_fd_sc_hd__inv_2
X_16087_ _18013_/Q vssd1 vssd1 vccd1 vccd1 _16087_/Y sky130_fd_sc_hd__inv_2
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13299_ _13299_/A _13299_/B _13299_/C _13299_/D vssd1 vssd1 vccd1 vccd1 _13299_/X
+ sky130_fd_sc_hd__or4_4
XFILLER_244_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_21_HCLK_A clkbuf_4_3_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19915_ _20006_/CLK _19915_/D repeater191/X vssd1 vssd1 vccd1 vccd1 _19915_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__14341__B1 _14279_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15038_ _18033_/Q _15035_/X _14992_/X _15037_/X vssd1 vssd1 vccd1 vccd1 _18033_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_130_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_84_HCLK_A clkbuf_4_13_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19846_ _19846_/CLK _19846_/D repeater270/X vssd1 vssd1 vccd1 vccd1 _19846_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__10902__B1 _10868_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19777_ _19780_/CLK _19777_/D repeater227/X vssd1 vssd1 vccd1 vccd1 _19777_/Q sky130_fd_sc_hd__dfrtp_1
X_16989_ _16988_/X _11409_/Y _17548_/S vssd1 vssd1 vccd1 vccd1 _16989_/X sky130_fd_sc_hd__mux2_1
XFILLER_110_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09530_ _19311_/Q vssd1 vssd1 vccd1 vccd1 _16587_/A sky130_fd_sc_hd__inv_2
XFILLER_95_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12655__B1 _12536_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18728_ _19224_/CLK _18728_/D repeater253/X vssd1 vssd1 vccd1 vccd1 _18728_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_83_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_224_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19369__RESET_B repeater241/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09461_ _10045_/A _19389_/Q _19929_/Q _09460_/Y vssd1 vssd1 vccd1 vccd1 _09461_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_236_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18659_ _20048_/CLK _18659_/D repeater210/X vssd1 vssd1 vccd1 vccd1 _18659_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_36_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16397__A1 _15846_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16397__B2 _16388_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09392_ _10023_/A _09391_/Y _19936_/Q _19396_/Q vssd1 vssd1 vccd1 vccd1 _09392_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12407__B1 _12406_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_224_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09501__A _19313_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16149__B2 _16003_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14332__B1 _14314_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_247_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_235_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19792__RESET_B repeater219/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09728_ _09728_/A _09728_/B _09728_/C _09728_/D vssd1 vssd1 vccd1 vccd1 _09729_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__12646__B1 hold250/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12102__A hold310/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_228_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09659_ _09746_/A _09745_/A _09747_/A _09744_/A vssd1 vssd1 vccd1 vccd1 _09660_/D
+ sky130_fd_sc_hd__or4_4
XFILLER_42_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11941__A _11979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17104__S _17544_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_243_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15413__A _15413_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12670_ _12677_/A vssd1 vssd1 vccd1 vccd1 _12670_/X sky130_fd_sc_hd__buf_1
XPHY_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_230_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_203_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11621_ _11621_/A _11635_/A vssd1 vssd1 vccd1 vccd1 _11622_/B sky130_fd_sc_hd__or2_1
XPHY_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16943__S _16946_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14340_ _18432_/Q _14336_/X _14277_/X _14338_/X vssd1 vssd1 vccd1 vccd1 _18432_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11552_ _11620_/A _11619_/C _11552_/C _11552_/D vssd1 vssd1 vccd1 vccd1 _11570_/B
+ sky130_fd_sc_hd__or4_4
XPHY_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10503_ _19538_/Q vssd1 vssd1 vccd1 vccd1 _10528_/C sky130_fd_sc_hd__inv_2
XPHY_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11483_ _11483_/A _11500_/A vssd1 vssd1 vccd1 vccd1 _11484_/B sky130_fd_sc_hd__or2_2
X_14271_ _14366_/A _14758_/B _14784_/C vssd1 vssd1 vccd1 vccd1 _14274_/A sky130_fd_sc_hd__or3_4
XPHY_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16010_ _18116_/Q vssd1 vssd1 vccd1 vccd1 _16010_/Y sky130_fd_sc_hd__inv_2
X_13222_ _18535_/Q _13222_/B vssd1 vssd1 vccd1 vccd1 _13223_/B sky130_fd_sc_hd__or2_1
XFILLER_183_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18674__RESET_B repeater252/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10434_ _10450_/A vssd1 vssd1 vccd1 vccd1 _10452_/A sky130_fd_sc_hd__inv_2
XFILLER_164_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10365_ _10361_/B _10335_/B _10364_/X _10319_/A _19859_/Q vssd1 vssd1 vccd1 vccd1
+ _19859_/D sky130_fd_sc_hd__a32o_1
X_13153_ _19174_/Q vssd1 vssd1 vccd1 vccd1 _13153_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14323__B1 _14279_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12104_ hold294/X vssd1 vssd1 vccd1 vccd1 _12104_/X sky130_fd_sc_hd__buf_2
X_17961_ _18869_/CLK _17961_/D vssd1 vssd1 vccd1 vccd1 _17961_/Q sky130_fd_sc_hd__dfxtp_1
X_13084_ _13084_/A _13172_/A vssd1 vssd1 vccd1 vccd1 _13085_/B sky130_fd_sc_hd__or2_2
X_10296_ _18590_/Q _15584_/A _18591_/Q vssd1 vssd1 vccd1 vccd1 _15588_/A sky130_fd_sc_hd__or3_1
XFILLER_239_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19700_ _19720_/CLK _19700_/D repeater201/X vssd1 vssd1 vccd1 vccd1 _19700_/Q sky130_fd_sc_hd__dfrtp_2
X_12035_ hold239/X vssd1 vssd1 vccd1 vccd1 _12035_/X sky130_fd_sc_hd__clkbuf_4
X_16912_ _16911_/X _09868_/A _17524_/S vssd1 vssd1 vccd1 vccd1 _16912_/X sky130_fd_sc_hd__mux2_2
XFILLER_78_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17892_ _16015_/Y _16016_/Y _16017_/Y _16018_/Y _17913_/S0 _19632_/Q vssd1 vssd1
+ vccd1 vccd1 _17892_/X sky130_fd_sc_hd__mux4_1
X_16843_ _16842_/X _11325_/Y _17493_/S vssd1 vssd1 vccd1 vccd1 _16843_/X sky130_fd_sc_hd__mux2_1
X_19631_ _19637_/CLK _19631_/D repeater258/X vssd1 vssd1 vccd1 vccd1 _19631_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_19_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19562_ _19577_/CLK _19562_/D repeater268/X vssd1 vssd1 vccd1 vccd1 _19562_/Q sky130_fd_sc_hd__dfrtp_1
X_16774_ _16773_/X _13557_/A _17386_/S vssd1 vssd1 vccd1 vccd1 _16774_/X sky130_fd_sc_hd__mux2_1
X_13986_ _18688_/Q vssd1 vssd1 vccd1 vccd1 _14018_/A sky130_fd_sc_hd__inv_2
XFILLER_81_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18513_ _19780_/CLK _18513_/D repeater227/X vssd1 vssd1 vccd1 vccd1 _18513_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_218_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15725_ _15725_/A _15725_/B vssd1 vssd1 vccd1 vccd1 _18658_/D sky130_fd_sc_hd__nor2_1
X_19493_ _19515_/CLK hold138/X repeater260/X vssd1 vssd1 vccd1 vccd1 _19493_/Q sky130_fd_sc_hd__dfrtp_1
X_12937_ _19265_/Q vssd1 vssd1 vccd1 vccd1 _12937_/Y sky130_fd_sc_hd__inv_2
XFILLER_233_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17014__S _17524_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18444_ _19865_/CLK _18444_/D vssd1 vssd1 vccd1 vccd1 _18444_/Q sky130_fd_sc_hd__dfxtp_1
X_15656_ _15661_/B vssd1 vssd1 vccd1 vccd1 _15656_/Y sky130_fd_sc_hd__inv_2
XPHY_4180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12868_ _18930_/Q vssd1 vssd1 vccd1 vccd1 _12870_/C sky130_fd_sc_hd__inv_2
XFILLER_233_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14607_ _18279_/Q _14599_/X _14606_/X _14602_/X vssd1 vssd1 vccd1 vccd1 _18279_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_33_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18375_ _19637_/CLK _18375_/D vssd1 vssd1 vccd1 vccd1 _18375_/Q sky130_fd_sc_hd__dfxtp_1
X_11819_ _19447_/Q _11814_/X _09079_/X _11815_/X vssd1 vssd1 vccd1 vccd1 _19447_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16853__S _17536_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15587_ _18591_/Q vssd1 vssd1 vccd1 vccd1 _15587_/Y sky130_fd_sc_hd__inv_2
XPHY_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12799_ _19238_/Q vssd1 vssd1 vccd1 vccd1 _12799_/Y sky130_fd_sc_hd__inv_2
XFILLER_239_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17326_ _17325_/X _09471_/A _17530_/S vssd1 vssd1 vccd1 vccd1 _17326_/X sky130_fd_sc_hd__mux2_2
XFILLER_175_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14538_ _18319_/Q _14530_/X _14537_/X _14533_/X vssd1 vssd1 vccd1 vccd1 _18319_/D
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_2_2_0_HCLK clkbuf_2_3_0_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_147_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16000__B1 _17503_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17257_ _16583_/Y _19078_/Q _17490_/S vssd1 vssd1 vccd1 vccd1 _17257_/X sky130_fd_sc_hd__mux2_1
X_14469_ _18358_/Q _14463_/X _14415_/X _14465_/X vssd1 vssd1 vccd1 vccd1 _18358_/D
+ sky130_fd_sc_hd__a22o_1
X_16208_ _16208_/A _16212_/B vssd1 vssd1 vccd1 vccd1 _16208_/Y sky130_fd_sc_hd__nor2_1
XFILLER_161_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17188_ _15768_/Y _14200_/Y _17546_/S vssd1 vssd1 vccd1 vccd1 _17188_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17684__S _17696_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16139_ _16134_/Y _15866_/A _16135_/Y _15854_/X _16138_/X vssd1 vssd1 vccd1 vccd1
+ _16139_/X sky130_fd_sc_hd__o221a_1
XFILLER_127_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15993__A _16634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18846__CLK _18866_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08961_ _19864_/Q _08956_/Y _10330_/A _18784_/Q _08960_/X vssd1 vssd1 vccd1 vccd1
+ _08969_/C sky130_fd_sc_hd__o221a_1
XFILLER_69_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19829_ _19842_/CLK _19829_/D repeater271/X vssd1 vssd1 vccd1 vccd1 _19829_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_217_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12628__B1 _12398_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09513_ _19296_/Q vssd1 vssd1 vccd1 vccd1 _09513_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_240_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09444_ _10036_/A _19380_/Q _10036_/A _19380_/Q vssd1 vssd1 vccd1 vccd1 _09444_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_212_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_197_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17319__A0 _17486_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09375_ _19386_/Q vssd1 vssd1 vccd1 vccd1 _09375_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16763__S _17534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16790__A1 _19155_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19621__CLK _19920_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14553__B1 hold330/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17594__S _17600_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10150_ _12257_/A _15883_/A vssd1 vssd1 vccd1 vccd1 _10186_/B sky130_fd_sc_hd__or2_2
XANTENNA__19973__RESET_B repeater244/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11936__A _11936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10081_ _10101_/A _10081_/B _10081_/C vssd1 vssd1 vccd1 vccd1 _10099_/A sky130_fd_sc_hd__or3_1
XFILLER_58_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_248_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_199_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19902__RESET_B repeater195/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16938__S _16946_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_235_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13840_ _19223_/Q vssd1 vssd1 vccd1 vccd1 _13840_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12619__B1 _12382_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15281__A1 _15205_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_244_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13771_ _18740_/Q _18741_/Q _13772_/S vssd1 vssd1 vccd1 vccd1 _18741_/D sky130_fd_sc_hd__mux2_1
XFILLER_216_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10983_ _10983_/A vssd1 vssd1 vccd1 vccd1 _10984_/B sky130_fd_sc_hd__inv_2
XFILLER_74_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16239__A _16634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_215_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15510_ _15518_/C vssd1 vssd1 vccd1 vccd1 _15510_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12722_ _18955_/Q vssd1 vssd1 vccd1 vccd1 _14812_/A sky130_fd_sc_hd__clkbuf_2
X_16490_ _20049_/Q vssd1 vssd1 vccd1 vccd1 _16490_/Y sky130_fd_sc_hd__inv_2
XFILLER_243_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15441_ _15443_/A _15441_/B vssd1 vssd1 vccd1 vccd1 _18549_/D sky130_fd_sc_hd__nor2_1
XPHY_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12653_ _18997_/Q _12650_/X _12602_/X _12651_/X vssd1 vssd1 vccd1 vccd1 _18997_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11604_ _19567_/Q _11603_/Y _11592_/X _11581_/B vssd1 vssd1 vccd1 vccd1 _19567_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18160_ _18198_/CLK _18160_/D vssd1 vssd1 vccd1 vccd1 _18160_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__18855__RESET_B repeater231/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15372_ _19788_/Q _10648_/B _10649_/B vssd1 vssd1 vccd1 vccd1 _15372_/X sky130_fd_sc_hd__a21bo_1
XPHY_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14792__B1 _14791_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12584_ _12600_/A vssd1 vssd1 vccd1 vccd1 _12584_/X sky130_fd_sc_hd__clkbuf_2
XPHY_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17111_ _17110_/X _13075_/A _17488_/S vssd1 vssd1 vccd1 vccd1 _17111_/X sky130_fd_sc_hd__mux2_1
XPHY_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14323_ _18439_/Q _14318_/X _14279_/X _14320_/X vssd1 vssd1 vccd1 vccd1 _18439_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11535_ _11535_/A vssd1 vssd1 vccd1 vccd1 _11535_/Y sky130_fd_sc_hd__inv_2
X_18091_ _18260_/CLK _18091_/D vssd1 vssd1 vccd1 vccd1 _18091_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_183_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17042_ _17473_/A0 _16658_/Y _17042_/S vssd1 vssd1 vccd1 vccd1 _17042_/X sky130_fd_sc_hd__mux2_1
X_14254_ _18474_/Q _14250_/X _13682_/X _14252_/X vssd1 vssd1 vccd1 vccd1 _18474_/D
+ sky130_fd_sc_hd__a22o_1
X_11466_ _11466_/A _11532_/A vssd1 vssd1 vccd1 vccd1 _11467_/B sky130_fd_sc_hd__or2_2
XFILLER_183_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13205_ _18894_/Q _13204_/Y _13180_/A _13205_/C1 vssd1 vssd1 vccd1 vccd1 _18894_/D
+ sky130_fd_sc_hd__o211a_1
X_10417_ _10419_/A vssd1 vssd1 vccd1 vccd1 _10417_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_152_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14185_ _19124_/Q vssd1 vssd1 vccd1 vccd1 _14185_/Y sky130_fd_sc_hd__inv_2
X_11397_ _19554_/Q vssd1 vssd1 vccd1 vccd1 _11624_/A sky130_fd_sc_hd__inv_2
XFILLER_152_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13136_ _19183_/Q vssd1 vssd1 vccd1 vccd1 _13136_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10348_ _10348_/A vssd1 vssd1 vccd1 vccd1 _10349_/B sky130_fd_sc_hd__inv_2
XFILLER_225_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18993_ _19608_/CLK _18993_/D hold355/X vssd1 vssd1 vccd1 vccd1 _18993_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_151_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17009__S _17546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15318__A _15318_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11846__A _12558_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10279_ _19642_/Q _19641_/Q _14301_/B vssd1 vssd1 vccd1 vccd1 _10279_/Y sky130_fd_sc_hd__o21ai_1
X_17944_ _18465_/CLK _17944_/D vssd1 vssd1 vccd1 vccd1 _17944_/Q sky130_fd_sc_hd__dfxtp_1
X_13067_ _13067_/A _13204_/A vssd1 vssd1 vccd1 vccd1 _13068_/B sky130_fd_sc_hd__or2_2
XFILLER_239_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19643__RESET_B repeater261/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater206 repeater207/X vssd1 vssd1 vccd1 vccd1 repeater206/X sky130_fd_sc_hd__buf_6
Xrepeater217 repeater234/X vssd1 vssd1 vccd1 vccd1 repeater217/X sky130_fd_sc_hd__buf_8
X_12018_ _19352_/Q _12016_/X hold314/X _12017_/X vssd1 vssd1 vccd1 vccd1 _19352_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_239_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrepeater228 repeater229/X vssd1 vssd1 vccd1 vccd1 repeater228/X sky130_fd_sc_hd__buf_6
X_17875_ _16097_/Y _16098_/Y _16099_/Y _16100_/Y _17908_/S0 _18759_/Q vssd1 vssd1
+ vccd1 vccd1 _17875_/X sky130_fd_sc_hd__mux4_1
XANTENNA__16848__S _17546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xrepeater239 repeater240/X vssd1 vssd1 vccd1 vccd1 repeater239/X sky130_fd_sc_hd__buf_6
XFILLER_239_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19614_ _20006_/CLK _19614_/D repeater191/X vssd1 vssd1 vccd1 vccd1 _19614_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17892__S0 _17913_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16826_ _16825_/X _09671_/Y _17523_/S vssd1 vssd1 vccd1 vccd1 _16826_/X sky130_fd_sc_hd__mux2_1
XFILLER_81_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_242_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19545_ _19545_/CLK _19545_/D repeater221/X vssd1 vssd1 vccd1 vccd1 _19545_/Q sky130_fd_sc_hd__dfrtp_2
X_16757_ vssd1 vssd1 vccd1 vccd1 _16757_/HI _16757_/LO sky130_fd_sc_hd__conb_1
XANTENNA__17549__A0 _15860_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13969_ _13964_/A _13964_/B _13964_/C vssd1 vssd1 vccd1 vccd1 _13970_/B sky130_fd_sc_hd__o21a_1
XFILLER_222_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_179_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15708_ _15715_/B vssd1 vssd1 vccd1 vccd1 _15713_/B sky130_fd_sc_hd__clkbuf_2
X_19476_ _19506_/CLK hold185/X repeater256/X vssd1 vssd1 vccd1 vccd1 _19476_/Q sky130_fd_sc_hd__dfrtp_1
X_16688_ _16688_/A vssd1 vssd1 vccd1 vccd1 _16688_/X sky130_fd_sc_hd__buf_1
XFILLER_62_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17679__S _17683_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09051__A hold294/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18427_ _19873_/CLK _18427_/D vssd1 vssd1 vccd1 vccd1 _18427_/Q sky130_fd_sc_hd__dfxtp_1
X_15639_ _18604_/Q vssd1 vssd1 vccd1 vccd1 _15642_/A sky130_fd_sc_hd__inv_2
XFILLER_210_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_203_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09160_ _09156_/A _09156_/B _20082_/Q _09159_/X vssd1 vssd1 vccd1 vccd1 _20082_/D
+ sky130_fd_sc_hd__o22a_1
XANTENNA__18596__RESET_B repeater267/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18358_ _19849_/CLK _18358_/D vssd1 vssd1 vccd1 vccd1 _18358_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14783__B1 _14782_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_187_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17309_ _16437_/Y _09313_/Y _19498_/Q vssd1 vssd1 vccd1 vccd1 _17309_/X sky130_fd_sc_hd__mux2_1
X_09091_ _20096_/Q _09084_/X _09090_/X _09087_/X vssd1 vssd1 vccd1 vccd1 _20096_/D
+ sky130_fd_sc_hd__a22o_1
X_18289_ _18435_/CLK _18289_/D vssd1 vssd1 vccd1 vccd1 _18289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09993_ _19946_/Q _09992_/Y _09968_/A _09856_/B vssd1 vssd1 vccd1 vccd1 _19946_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_135_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08944_ _19861_/Q vssd1 vssd1 vccd1 vccd1 _10327_/A sky130_fd_sc_hd__inv_2
XANTENNA__10660__A _10660_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17883__S0 _17913_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_217_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_226_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12077__A1 _19323_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_231_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_hold149_A HWRITE vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17589__S _17600_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09427_ _09425_/Y _19397_/Q _19937_/Q _09426_/Y vssd1 vssd1 vccd1 vccd1 _09427_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__15898__A _16634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09358_ _20019_/Q vssd1 vssd1 vccd1 vccd1 _09479_/A sky130_fd_sc_hd__inv_2
XANTENNA__14774__B1 _14745_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold316_A HWDATA[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09289_ _20048_/Q _09285_/X _09079_/X _09287_/X vssd1 vssd1 vccd1 vccd1 _20048_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_165_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11320_ _18990_/Q vssd1 vssd1 vccd1 vccd1 _11320_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14526__B1 _14513_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11251_ _19594_/Q _19008_/Q _11474_/A _11250_/Y vssd1 vssd1 vccd1 vccd1 _11261_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_109_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_181_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_181_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10202_ _19830_/Q _19657_/Q _10200_/Y _10957_/A vssd1 vssd1 vccd1 vccd1 _10209_/B
+ sky130_fd_sc_hd__o22a_1
X_11182_ _17708_/X _11176_/X _19623_/Q _11178_/X vssd1 vssd1 vccd1 vccd1 _19623_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_79_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10133_ _10133_/A _10133_/B _10133_/C vssd1 vssd1 vccd1 vccd1 _10133_/X sky130_fd_sc_hd__and3_1
XFILLER_192_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15990_ _17498_/X vssd1 vssd1 vccd1 vccd1 _15990_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10064_ _10044_/A _10044_/B _10032_/A _10062_/Y vssd1 vssd1 vccd1 vccd1 _19928_/D
+ sky130_fd_sc_hd__a211oi_2
XANTENNA_input34_A HRESETn vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14941_ _14941_/A vssd1 vssd1 vccd1 vccd1 _14941_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_248_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_82_HCLK clkbuf_4_13_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19282_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_94_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19054__RESET_B repeater267/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14977__A hold248/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17660_ _15595_/X _19029_/Q _17664_/S vssd1 vssd1 vccd1 vccd1 _18592_/D sky130_fd_sc_hd__mux2_1
XANTENNA__17874__S0 _19633_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14872_ _14872_/A vssd1 vssd1 vccd1 vccd1 _14873_/A sky130_fd_sc_hd__inv_2
XFILLER_36_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16611_ _16815_/X _16573_/X _16821_/X _16574_/X _16610_/X vssd1 vssd1 vccd1 vccd1
+ _16614_/B sky130_fd_sc_hd__o221a_4
XFILLER_91_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13823_ _13909_/B _13823_/B vssd1 vssd1 vccd1 vccd1 _13929_/A sky130_fd_sc_hd__or2_1
X_17591_ _15355_/X _19712_/Q _17600_/S vssd1 vssd1 vccd1 vccd1 _17591_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19330_ _19513_/CLK _19330_/D repeater259/X vssd1 vssd1 vccd1 vccd1 _19330_/Q sky130_fd_sc_hd__dfrtp_1
X_16542_ _16542_/A _16544_/B vssd1 vssd1 vccd1 vccd1 _16542_/Y sky130_fd_sc_hd__nor2_1
XFILLER_141_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13754_ _13749_/Y _17763_/S _13753_/Y vssd1 vssd1 vccd1 vccd1 _13756_/A sky130_fd_sc_hd__o21ai_1
XFILLER_232_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10966_ _10966_/A _10975_/A vssd1 vssd1 vccd1 vccd1 _10973_/A sky130_fd_sc_hd__or2_2
XFILLER_189_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12705_ _18961_/Q _12677_/A _12541_/X _12678_/A vssd1 vssd1 vccd1 vccd1 _18961_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17499__S _17564_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19261_ _20035_/CLK _19261_/D repeater242/X vssd1 vssd1 vccd1 vccd1 _19261_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_189_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16473_ _19447_/Q _17517_/S vssd1 vssd1 vccd1 vccd1 _16473_/Y sky130_fd_sc_hd__nand2_1
XFILLER_71_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13685_ _13686_/A vssd1 vssd1 vccd1 vccd1 _13685_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_repeater173_A _17524_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10897_ _19691_/Q _10893_/X _10882_/X _10895_/X vssd1 vssd1 vccd1 vccd1 _19691_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_231_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18212_ _18333_/CLK _18212_/D vssd1 vssd1 vccd1 vccd1 _18212_/Q sky130_fd_sc_hd__dfxtp_1
X_15424_ _19615_/Q _11160_/B _11161_/B vssd1 vssd1 vccd1 vccd1 _15424_/X sky130_fd_sc_hd__a21bo_1
XPHY_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12636_ _12650_/A vssd1 vssd1 vccd1 vccd1 _12636_/X sky130_fd_sc_hd__clkbuf_2
X_19192_ _20035_/CLK _19192_/D repeater242/X vssd1 vssd1 vccd1 vccd1 _19192_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18143_ _18145_/CLK _18143_/D vssd1 vssd1 vccd1 vccd1 _18143_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15355_ _18499_/Q _14229_/B _14230_/B vssd1 vssd1 vccd1 vccd1 _15355_/X sky130_fd_sc_hd__a21bo_1
XFILLER_184_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12567_ _19053_/Q _12560_/X _12384_/X _12563_/X vssd1 vssd1 vccd1 vccd1 _19053_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14306_ _18449_/Q _14303_/X _14273_/X _14305_/X vssd1 vssd1 vccd1 vccd1 _18449_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11518_ _19593_/Q _11517_/Y _11504_/X _11474_/B vssd1 vssd1 vccd1 vccd1 _19593_/D
+ sky130_fd_sc_hd__o211a_1
X_18074_ _18198_/CLK _18074_/D vssd1 vssd1 vccd1 vccd1 _18074_/Q sky130_fd_sc_hd__dfxtp_1
X_15286_ _18629_/Q _15286_/B vssd1 vssd1 vccd1 vccd1 _15287_/C sky130_fd_sc_hd__nand2_1
XFILLER_172_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12498_ _12505_/A vssd1 vssd1 vccd1 vccd1 _12498_/X sky130_fd_sc_hd__clkbuf_2
Xhold208 hold208/A vssd1 vssd1 vccd1 vccd1 hold208/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19895__RESET_B repeater205/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold219 hold219/A vssd1 vssd1 vccd1 vccd1 hold219/X sky130_fd_sc_hd__dlygate4sd3_1
X_17025_ _16471_/Y _19374_/Q _17413_/S vssd1 vssd1 vccd1 vccd1 _17025_/X sky130_fd_sc_hd__mux2_1
XFILLER_236_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14237_ _18670_/Q _14236_/X _18669_/Q _17600_/S vssd1 vssd1 vccd1 vccd1 _18670_/D
+ sky130_fd_sc_hd__a22o_1
X_11449_ _19548_/Q _11444_/Y _19575_/Q _11445_/Y _11448_/X vssd1 vssd1 vccd1 vccd1
+ _11456_/C sky130_fd_sc_hd__o221a_1
XFILLER_113_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20024__CLK _20091_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14168_ _19096_/Q vssd1 vssd1 vccd1 vccd1 _14168_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13119_ _19186_/Q vssd1 vssd1 vccd1 vccd1 _13119_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18071__CLK _18169_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18976_ _19597_/CLK _18976_/D repeater282/X vssd1 vssd1 vccd1 vccd1 _18976_/Q sky130_fd_sc_hd__dfrtp_1
X_14099_ _14118_/A vssd1 vssd1 vccd1 vccd1 _14135_/B sky130_fd_sc_hd__buf_2
XFILLER_112_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17927_ _19462_/CLK _19399_/Q vssd1 vssd1 vccd1 vccd1 _17927_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09172__B2 _09165_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17865__S0 _17908_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17858_ _16287_/Y _16288_/Y _16289_/Y _16290_/Y _17908_/S0 _18759_/Q vssd1 vssd1
+ vccd1 vccd1 _17858_/X sky130_fd_sc_hd__mux4_2
XFILLER_38_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_208_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16809_ _16808_/X _13554_/A _17536_/S vssd1 vssd1 vccd1 vccd1 _16809_/X sky130_fd_sc_hd__mux2_1
XFILLER_81_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_139_HCLK_A clkbuf_4_3_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17789_ _17785_/X _17786_/X _17787_/X _17788_/X _19647_/Q _19648_/Q vssd1 vssd1 vccd1
+ vccd1 _17789_/X sky130_fd_sc_hd__mux4_2
XFILLER_35_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19528_ _19771_/CLK _19528_/D repeater189/X vssd1 vssd1 vccd1 vccd1 _19528_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_34_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19459_ _19462_/CLK _19459_/D repeater272/X vssd1 vssd1 vccd1 vccd1 _19459_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_22_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_222_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16745__B2 _19627_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17202__S _17536_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09212_ _18649_/Q _09212_/B vssd1 vssd1 vccd1 vccd1 _09213_/A sky130_fd_sc_hd__nand2_1
XFILLER_139_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14756__B1 _14691_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_210_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09143_ _15322_/B _09141_/Y _15322_/A _09140_/Y vssd1 vssd1 vccd1 vccd1 _20086_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_108_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_175_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09074_ hold251/X vssd1 vssd1 vccd1 vccd1 hold250/A sky130_fd_sc_hd__buf_4
XFILLER_162_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_190_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09976_ _19956_/Q _09975_/Y _09865_/B _09964_/X vssd1 vssd1 vccd1 vccd1 _19956_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_162_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08927_ _19867_/Q vssd1 vssd1 vccd1 vccd1 _08927_/Y sky130_fd_sc_hd__inv_2
X_20096_ _20107_/CLK _20096_/D repeater233/X vssd1 vssd1 vccd1 vccd1 _20096_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_58_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_218_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17856__S0 _17908_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11933__B _12372_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13247__B1 _12533_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20052__RESET_B repeater207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10820_ _12257_/A _15845_/D vssd1 vssd1 vccd1 vccd1 _10841_/A sky130_fd_sc_hd__or2_2
XANTENNA__14995__B1 _14992_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_214_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_232_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10751_ _19756_/Q _10742_/A _10427_/X _10743_/A vssd1 vssd1 vccd1 vccd1 _19756_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11273__A2 _19003_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_201_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17112__S _17547_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_240_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13470_ _13470_/A _13470_/B vssd1 vssd1 vccd1 vccd1 _13470_/Y sky130_fd_sc_hd__nor2_1
XFILLER_231_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10682_ _17743_/X _10676_/X _19782_/Q _10677_/X vssd1 vssd1 vccd1 vccd1 _19782_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_200_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12421_ _12428_/A vssd1 vssd1 vccd1 vccd1 _12421_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_200_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10233__B1 _19832_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15140_ _17965_/Q _15134_/X _10698_/X _15136_/X vssd1 vssd1 vccd1 vccd1 _17965_/D
+ sky130_fd_sc_hd__a22o_1
X_12352_ _12361_/A vssd1 vssd1 vccd1 vccd1 _12352_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_127_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11303_ _19605_/Q _11300_/Y _11472_/A _18974_/Q _11302_/X vssd1 vssd1 vccd1 vccd1
+ _11303_/X sky130_fd_sc_hd__a221o_1
X_15071_ _15072_/A vssd1 vssd1 vccd1 vccd1 _15071_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__12780__A _19247_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12283_ _12298_/A vssd1 vssd1 vccd1 vccd1 _12283_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_181_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14022_ _14022_/A _14022_/B vssd1 vssd1 vccd1 vccd1 _14115_/A sky130_fd_sc_hd__or2_1
XANTENNA__13722__A1 _18757_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11234_ _11471_/A _19005_/Q _11462_/A _18995_/Q vssd1 vssd1 vccd1 vccd1 _11234_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_106_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18830_ _19255_/CLK _18830_/D repeater239/X vssd1 vssd1 vccd1 vccd1 _18830_/Q sky130_fd_sc_hd__dfrtp_1
X_11165_ _19620_/Q _11165_/B vssd1 vssd1 vccd1 vccd1 _11166_/B sky130_fd_sc_hd__or2_1
XFILLER_96_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10116_ _18563_/Q _15470_/A vssd1 vssd1 vccd1 vccd1 _15474_/A sky130_fd_sc_hd__or2_2
XANTENNA_output140_A _19672_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15973_ _15973_/A vssd1 vssd1 vccd1 vccd1 _15973_/X sky130_fd_sc_hd__clkbuf_2
X_11096_ _11096_/A vssd1 vssd1 vccd1 vccd1 _15094_/B sky130_fd_sc_hd__buf_1
X_18761_ _20124_/CLK _18761_/D repeater196/X vssd1 vssd1 vccd1 vccd1 _18761_/Q sky130_fd_sc_hd__dfrtp_2
X_17712_ _15428_/X _19765_/Q _18546_/D vssd1 vssd1 vccd1 vccd1 _17712_/X sky130_fd_sc_hd__mux2_1
X_10047_ _10047_/A _10059_/A _10047_/C vssd1 vssd1 vccd1 vccd1 _10055_/A sky130_fd_sc_hd__or3_4
X_14924_ _18097_/Q _14920_/X _14921_/X _14923_/X vssd1 vssd1 vccd1 vccd1 _18097_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_236_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17847__S0 _17908_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18692_ _18701_/CLK _18692_/D hold359/X vssd1 vssd1 vccd1 vccd1 _18692_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_236_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14855_ _18138_/Q _14846_/A _14842_/X _14847_/A vssd1 vssd1 vccd1 vccd1 _18138_/D
+ sky130_fd_sc_hd__a22o_1
X_17643_ _15666_/Y _19046_/Q _17655_/S vssd1 vssd1 vccd1 vccd1 _18609_/D sky130_fd_sc_hd__mux2_1
XANTENNA__16975__A1 _19081_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13806_ _18704_/Q vssd1 vssd1 vccd1 vccd1 _13964_/B sky130_fd_sc_hd__inv_2
X_17574_ _15412_/X _19769_/Q _17584_/S vssd1 vssd1 vccd1 vccd1 _17574_/X sky130_fd_sc_hd__mux2_1
XANTENNA__14986__B1 _14793_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14786_ _14786_/A vssd1 vssd1 vccd1 vccd1 _14787_/A sky130_fd_sc_hd__inv_2
X_11998_ _11998_/A _15769_/A vssd1 vssd1 vccd1 vccd1 _12043_/A sky130_fd_sc_hd__or2_2
XFILLER_91_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19313_ _19314_/CLK _19313_/D repeater214/X vssd1 vssd1 vccd1 vccd1 _19313_/Q sky130_fd_sc_hd__dfrtp_2
X_16525_ _19451_/Q vssd1 vssd1 vccd1 vccd1 _16525_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13737_ _13737_/A _13737_/B vssd1 vssd1 vccd1 vccd1 _13738_/A sky130_fd_sc_hd__or2_1
XFILLER_31_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10949_ _10949_/A vssd1 vssd1 vccd1 vccd1 _10950_/A sky130_fd_sc_hd__inv_2
XANTENNA__12461__A1 _19112_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_189_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17022__S _17543_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16456_ _16452_/Y _15971_/X _15391_/A _15973_/X _16455_/X vssd1 vssd1 vccd1 vccd1
+ _16456_/X sky130_fd_sc_hd__o221a_1
X_19244_ _19282_/CLK _19244_/D repeater214/X vssd1 vssd1 vccd1 vccd1 _19244_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_31_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13668_ _18780_/Q _13664_/X hold259/X _13665_/X vssd1 vssd1 vccd1 vccd1 _18780_/D
+ sky130_fd_sc_hd__a22o_1
X_15407_ _15413_/A _17577_/X vssd1 vssd1 vccd1 vccd1 _18535_/D sky130_fd_sc_hd__and2_1
XPHY_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_176_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12619_ _19021_/Q _12613_/X _12382_/X _12616_/X vssd1 vssd1 vccd1 vccd1 _19021_/D
+ sky130_fd_sc_hd__a22o_1
X_19175_ _19288_/CLK _19175_/D repeater212/X vssd1 vssd1 vccd1 vccd1 _19175_/Q sky130_fd_sc_hd__dfrtp_1
X_16387_ _16384_/Y _15971_/X _15333_/A _15838_/X _16386_/X vssd1 vssd1 vccd1 vccd1
+ _16387_/X sky130_fd_sc_hd__o221a_1
XFILLER_157_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16861__S _17513_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13599_ _13537_/B _13599_/A2 _18813_/Q _13598_/Y _13560_/X vssd1 vssd1 vccd1 vccd1
+ _18813_/D sky130_fd_sc_hd__o221a_1
XFILLER_247_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18126_ _18137_/CLK _18126_/D vssd1 vssd1 vccd1 vccd1 _18126_/Q sky130_fd_sc_hd__dfxtp_1
X_15338_ _15364_/A vssd1 vssd1 vccd1 vccd1 _15347_/A sky130_fd_sc_hd__buf_1
XFILLER_184_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11972__B1 _09075_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18057_ _18169_/CLK _18057_/D vssd1 vssd1 vccd1 vccd1 _18057_/Q sky130_fd_sc_hd__dfxtp_1
X_15269_ _15443_/A _15437_/B _15259_/B _15268_/X vssd1 vssd1 vccd1 vccd1 _18634_/D
+ sky130_fd_sc_hd__o31ai_1
XFILLER_172_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20038__SET_B repeater208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17008_ _17007_/X _15688_/A _17318_/S vssd1 vssd1 vccd1 vccd1 _17008_/X sky130_fd_sc_hd__mux2_1
XFILLER_99_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17692__S _17696_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09830_ _19956_/Q vssd1 vssd1 vccd1 vccd1 _09864_/A sky130_fd_sc_hd__inv_2
XFILLER_59_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14269__A2 _14259_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09761_ _09761_/A vssd1 vssd1 vccd1 vccd1 _09761_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18959_ _18959_/CLK _18959_/D repeater257/X vssd1 vssd1 vccd1 vccd1 _18959_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__09409__A2_N _19395_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18958__RESET_B repeater257/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17838__S0 _17908_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09692_ _19974_/Q _19403_/Q _09635_/B _09691_/Y vssd1 vssd1 vccd1 vccd1 _09692_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_239_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrebuffer12 _13085_/B vssd1 vssd1 vccd1 vccd1 _13171_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XANTENNA__19982__CLK _19992_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer23 _14012_/C vssd1 vssd1 vccd1 vccd1 _14134_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_54_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_215_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrebuffer34 _14005_/B vssd1 vssd1 vccd1 vccd1 _14149_/B1 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer45 _13083_/B vssd1 vssd1 vccd1 vccd1 _13177_/B1 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer56 _13081_/B vssd1 vssd1 vccd1 vccd1 _13178_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer67 _09488_/B vssd1 vssd1 vccd1 vccd1 _09579_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_214_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrebuffer78 _09875_/B vssd1 vssd1 vccd1 vccd1 _09956_/A2 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer89 _09476_/B vssd1 vssd1 vccd1 vccd1 _09600_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_23_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12452__A1 _19119_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14729__B1 _14691_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_195_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_194_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrebuffer102 _09620_/A vssd1 vssd1 vccd1 vccd1 _10025_/A sky130_fd_sc_hd__buf_2
XANTENNA__16771__S _17548_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrebuffer113 _13087_/B vssd1 vssd1 vccd1 vccd1 _13168_/A2 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer124 _09469_/B vssd1 vssd1 vccd1 vccd1 _09616_/C1 sky130_fd_sc_hd__dlygate4sd1_1
X_09126_ _17605_/S _13493_/A vssd1 vssd1 vccd1 vccd1 _09139_/B sky130_fd_sc_hd__or2_1
XANTENNA__19746__RESET_B repeater205/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09057_ hold234/X vssd1 vssd1 vccd1 vccd1 hold233/A sky130_fd_sc_hd__buf_4
XFILLER_136_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11928__B _12309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09959_ _09873_/A _09873_/B _09990_/A _09957_/Y vssd1 vssd1 vccd1 vccd1 _19965_/D
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__17107__S _17535_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20079_ _20079_/CLK _20079_/D repeater205/X vssd1 vssd1 vccd1 vccd1 _20079_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__18699__RESET_B hold351/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17829__S0 _18751_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12970_ _18946_/Q _18945_/Q _12970_/C vssd1 vssd1 vccd1 vccd1 _12970_/X sky130_fd_sc_hd__and3_1
XANTENNA__15209__A1 _15205_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12140__B1 _12076_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_218_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11921_ _19404_/Q _11914_/X _11920_/X _11915_/X vssd1 vssd1 vccd1 vccd1 _19404_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18628__RESET_B repeater221/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16946__S _16946_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_246_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14640_ _18258_/Q _14631_/A _14626_/X _14632_/A vssd1 vssd1 vccd1 vccd1 _18258_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11852_ _19329_/Q vssd1 vssd1 vccd1 vccd1 _11853_/A sky130_fd_sc_hd__clkbuf_2
XPHY_4554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09439__A2 _09374_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_122_HCLK_A clkbuf_4_4_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_112_HCLK clkbuf_opt_0_HCLK/A vssd1 vssd1 vccd1 vccd1 _18701_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_4576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_214_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10803_ _10801_/A _10801_/B _10788_/Y _10801_/Y vssd1 vssd1 vccd1 vccd1 _19734_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_60_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14571_ _14598_/A _14598_/B _14571_/C vssd1 vssd1 vccd1 vccd1 _14573_/A sky130_fd_sc_hd__or3_4
XFILLER_60_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11783_ _11821_/A vssd1 vssd1 vccd1 vccd1 _11800_/A sky130_fd_sc_hd__buf_2
XFILLER_214_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16310_ _16301_/Y _15828_/X _16304_/X _16309_/X vssd1 vssd1 vccd1 vccd1 _16310_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_198_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10454__B1 _10418_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13522_ _15145_/A vssd1 vssd1 vccd1 vccd1 _14857_/A sky130_fd_sc_hd__clkbuf_2
X_10734_ _10734_/A _19530_/Q _10734_/C _19529_/Q vssd1 vssd1 vccd1 vccd1 _10735_/B
+ sky130_fd_sc_hd__or4b_4
XPHY_3886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_186_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17290_ _17289_/X _09475_/A _17414_/S vssd1 vssd1 vccd1 vccd1 _17290_/X sky130_fd_sc_hd__mux2_2
XPHY_3897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_198_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_186_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16241_ _17384_/X _16555_/A _17382_/X _16556_/A vssd1 vssd1 vccd1 vccd1 _16241_/Y
+ sky130_fd_sc_hd__a22oi_4
X_13453_ _13453_/A vssd1 vssd1 vccd1 vccd1 _13453_/Y sky130_fd_sc_hd__inv_2
X_10665_ _17730_/X _10661_/X _19795_/Q _10663_/X vssd1 vssd1 vccd1 vccd1 _19795_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_40_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19487__RESET_B repeater260/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12404_ hold301/X vssd1 vssd1 vccd1 vccd1 _12404_/X sky130_fd_sc_hd__clkbuf_2
X_16172_ _18233_/Q _18232_/Q _18231_/Q _18230_/Q vssd1 vssd1 vccd1 vccd1 _16172_/Y
+ sky130_fd_sc_hd__nor4_2
X_13384_ _20115_/Q _18861_/Q _20115_/Q _18861_/Q vssd1 vssd1 vccd1 vccd1 _13384_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_10596_ _10616_/B _10613_/B vssd1 vssd1 vccd1 vccd1 _15298_/A sky130_fd_sc_hd__or2_1
XANTENNA__11954__B1 _09039_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_182_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15123_ _15123_/A vssd1 vssd1 vccd1 vccd1 _15124_/A sky130_fd_sc_hd__inv_2
XANTENNA__19416__RESET_B repeater210/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12335_ _12335_/A vssd1 vssd1 vccd1 vccd1 _12335_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_182_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19931_ _19933_/CLK _19931_/D repeater236/X vssd1 vssd1 vccd1 vccd1 _19931_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_154_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15054_ _18021_/Q _15047_/X _15002_/X _15049_/X vssd1 vssd1 vccd1 vccd1 _18021_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_5_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12266_ _19222_/Q _12260_/X _12076_/X _12263_/X vssd1 vssd1 vccd1 vccd1 _19222_/D
+ sky130_fd_sc_hd__a22o_1
X_14005_ _14005_/A _14005_/B vssd1 vssd1 vccd1 vccd1 _14145_/A sky130_fd_sc_hd__or2_1
X_11217_ _19013_/Q vssd1 vssd1 vccd1 vccd1 _11217_/Y sky130_fd_sc_hd__inv_2
X_19862_ _19865_/CLK _19862_/D repeater262/X vssd1 vssd1 vccd1 vccd1 _19862_/Q sky130_fd_sc_hd__dfrtp_1
X_12197_ _19254_/Q _12189_/X _12080_/X _12192_/X vssd1 vssd1 vccd1 vccd1 _19254_/D
+ sky130_fd_sc_hd__a22o_1
Xoutput81 _16524_/Y vssd1 vssd1 vccd1 vccd1 HRDATA[11] sky130_fd_sc_hd__clkbuf_2
X_18813_ _19314_/CLK _18813_/D repeater239/X vssd1 vssd1 vccd1 vccd1 _18813_/Q sky130_fd_sc_hd__dfrtp_1
Xoutput92 _16641_/Y vssd1 vssd1 vccd1 vccd1 HRDATA[21] sky130_fd_sc_hd__clkbuf_2
X_11148_ _14598_/B _14301_/B _11053_/B vssd1 vssd1 vccd1 vccd1 _11148_/X sky130_fd_sc_hd__a21bo_1
XFILLER_68_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19793_ _19794_/CLK _19793_/D repeater219/X vssd1 vssd1 vccd1 vccd1 _19793_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_233_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17017__S _17545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18744_ _20066_/CLK _18744_/D repeater209/X vssd1 vssd1 vccd1 vccd1 _18744_/Q sky130_fd_sc_hd__dfrtp_1
X_11079_ _15858_/A _15858_/B _15190_/A _15899_/A vssd1 vssd1 vccd1 vccd1 _15318_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_83_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15956_ _18768_/Q vssd1 vssd1 vccd1 vccd1 _15956_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14907_ _15109_/A _15145_/B _15157_/C vssd1 vssd1 vccd1 vccd1 _14909_/A sky130_fd_sc_hd__or3_4
X_18675_ _18686_/CLK _18675_/D repeater252/X vssd1 vssd1 vccd1 vccd1 _18675_/Q sky130_fd_sc_hd__dfrtp_2
X_15887_ _16238_/A vssd1 vssd1 vccd1 vccd1 _15887_/X sky130_fd_sc_hd__buf_2
XANTENNA__16856__S _17524_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17626_ _19893_/Q _19746_/Q _17630_/S vssd1 vssd1 vccd1 vccd1 _17626_/X sky130_fd_sc_hd__mux2_1
X_14838_ _18150_/Q _14832_/X _14810_/X _14834_/X vssd1 vssd1 vccd1 vccd1 _18150_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_17_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14769_ _18186_/Q _14760_/A _14693_/X _14761_/A vssd1 vssd1 vccd1 vccd1 _18186_/D
+ sky130_fd_sc_hd__a22o_1
X_17557_ _17556_/X _19874_/Q _19497_/Q vssd1 vssd1 vccd1 vccd1 _17557_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12434__B2 _12402_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12685__A _12699_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10445__B1 _09079_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_44_HCLK_A clkbuf_opt_2_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_232_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16508_ _16638_/A vssd1 vssd1 vccd1 vccd1 _16508_/X sky130_fd_sc_hd__buf_1
X_17488_ _17487_/X _13061_/A _17488_/S vssd1 vssd1 vccd1 vccd1 _17488_/X sky130_fd_sc_hd__mux2_1
XANTENNA__17373__A1 _17859_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19227_ _19320_/CLK _19227_/D repeater237/X vssd1 vssd1 vccd1 vccd1 _19227_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__17687__S _17696_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16439_ _19032_/Q vssd1 vssd1 vccd1 vccd1 _16439_/Y sky130_fd_sc_hd__inv_2
XFILLER_176_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19158_ _19293_/CLK _19158_/D repeater212/X vssd1 vssd1 vccd1 vccd1 _19158_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_145_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11945__B1 hold288/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18109_ _18765_/CLK _18109_/D vssd1 vssd1 vccd1 vccd1 _18109_/Q sky130_fd_sc_hd__dfxtp_1
X_19089_ _19609_/CLK _19089_/D hold357/X vssd1 vssd1 vccd1 vccd1 _19089_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__14405__A _14405_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20002_ _20003_/CLK _20002_/D repeater185/X vssd1 vssd1 vccd1 vccd1 _20002_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_99_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16636__B1 _16875_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09813_ _09813_/A _09813_/B _09813_/C vssd1 vssd1 vccd1 vccd1 _19973_/D sky130_fd_sc_hd__nor3_1
XFILLER_113_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11764__A _11771_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18792__RESET_B repeater261/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09744_ _09744_/A _09744_/B vssd1 vssd1 vccd1 vccd1 _09778_/A sky130_fd_sc_hd__or2_1
XFILLER_67_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_228_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_135_HCLK clkbuf_4_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19997_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_227_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18721__RESET_B repeater253/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09675_ _19999_/Q _09671_/Y _19978_/Q _09672_/Y _09674_/X vssd1 vssd1 vccd1 vccd1
+ _09689_/A sky130_fd_sc_hd__o221a_1
XFILLER_228_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16766__S _17534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_243_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17061__A0 _15768_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_227_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_243_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19998__RESET_B repeater192/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10436__B1 _09058_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_hold131_A HADDR[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17597__S _17600_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18752__CLK _19900_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10450_ _10450_/A vssd1 vssd1 vccd1 vccd1 _10450_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_108_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09109_ _20091_/Q _09041_/A _09108_/X _09043_/A vssd1 vssd1 vccd1 vccd1 _20091_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_108_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10381_ _10381_/A vssd1 vssd1 vccd1 vccd1 _19855_/D sky130_fd_sc_hd__inv_2
XFILLER_164_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12120_ _19301_/Q _12114_/X _11975_/X _12115_/X vssd1 vssd1 vccd1 vccd1 _19301_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13689__B1 _13678_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12051_ _19331_/Q _12016_/A _11926_/X _12017_/A vssd1 vssd1 vccd1 vccd1 _19331_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_89_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11002_ _19659_/Q _11002_/B vssd1 vssd1 vccd1 vccd1 _11002_/Y sky130_fd_sc_hd__nor2_1
XFILLER_120_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18809__RESET_B repeater217/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18132__CLK _18198_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14102__A1 _18701_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_237_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15810_ _18130_/Q vssd1 vssd1 vccd1 vccd1 _15810_/Y sky130_fd_sc_hd__inv_2
X_16790_ _16789_/X _19155_/Q _17548_/S vssd1 vssd1 vccd1 vccd1 _16790_/X sky130_fd_sc_hd__mux2_1
XFILLER_93_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12113__B1 _12032_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15741_ _18670_/Q _18668_/Q _18669_/Q _15740_/X vssd1 vssd1 vccd1 vccd1 _18487_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12953_ _12952_/Y _18942_/Q _19285_/Q _12967_/C vssd1 vssd1 vccd1 vccd1 _12953_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_218_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17052__A0 _17473_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11904_ _19413_/Q _11898_/X _09067_/X _11899_/X vssd1 vssd1 vccd1 vccd1 _19413_/D
+ sky130_fd_sc_hd__a22o_1
X_15672_ _18611_/Q vssd1 vssd1 vccd1 vccd1 _15672_/Y sky130_fd_sc_hd__inv_2
X_18460_ _18460_/CLK _18460_/D vssd1 vssd1 vccd1 vccd1 _18460_/Q sky130_fd_sc_hd__dfxtp_1
X_12884_ _12967_/C _12978_/A vssd1 vssd1 vccd1 vccd1 _12885_/B sky130_fd_sc_hd__or2_2
XPHY_4340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14623_ _18269_/Q _14616_/X _09180_/X _14618_/X vssd1 vssd1 vccd1 vccd1 _18269_/D
+ sky130_fd_sc_hd__a22o_1
X_17411_ _17410_/X _09851_/A _17518_/S vssd1 vssd1 vccd1 vccd1 _17411_/X sky130_fd_sc_hd__mux2_1
XPHY_4373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18391_ _18441_/CLK _18391_/D vssd1 vssd1 vccd1 vccd1 _18391_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11835_ _19437_/Q vssd1 vssd1 vccd1 vccd1 _15643_/A sky130_fd_sc_hd__clkbuf_2
XPHY_4384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output103_A _16743_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19668__RESET_B repeater270/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17342_ _16364_/X _18778_/Q _17566_/S vssd1 vssd1 vccd1 vccd1 _17342_/X sky130_fd_sc_hd__mux2_1
XFILLER_214_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14554_ _18308_/Q _14547_/A _14513_/X _14548_/A vssd1 vssd1 vccd1 vccd1 _18308_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_198_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11766_ hold177/X _11764_/X _19480_/Q _11765_/X vssd1 vssd1 vccd1 vccd1 hold179/A
+ sky130_fd_sc_hd__o22a_1
XPHY_3694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_201_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13505_ _14696_/B vssd1 vssd1 vccd1 vccd1 _13506_/A sky130_fd_sc_hd__clkbuf_2
X_10717_ _10842_/A vssd1 vssd1 vccd1 vccd1 _15971_/A sky130_fd_sc_hd__clkbuf_2
XPHY_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17273_ _15768_/Y _11282_/Y _17546_/S vssd1 vssd1 vccd1 vccd1 _17273_/X sky130_fd_sc_hd__mux2_1
XPHY_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14485_ _18349_/Q _14478_/X _12726_/X _14480_/X vssd1 vssd1 vccd1 vccd1 _18349_/D
+ sky130_fd_sc_hd__a22o_1
X_11697_ _19524_/Q _11690_/X _10863_/X _11692_/X vssd1 vssd1 vccd1 vccd1 _19524_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_158_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15905__A2 _16506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17300__S _17535_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16224_ _16219_/Y _16053_/X _16220_/Y _15828_/A _16223_/X vssd1 vssd1 vccd1 vccd1
+ _16224_/X sky130_fd_sc_hd__o221a_1
X_19012_ _19597_/CLK _19012_/D repeater281/X vssd1 vssd1 vccd1 vccd1 _19012_/Q sky130_fd_sc_hd__dfrtp_2
X_13436_ _18864_/Q _13352_/C _13361_/Y _13351_/A _13421_/X vssd1 vssd1 vccd1 vccd1
+ _18864_/D sky130_fd_sc_hd__o221a_1
XFILLER_173_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17107__A1 _20105_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10648_ _19788_/Q _10648_/B vssd1 vssd1 vccd1 vccd1 _10649_/B sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_16_HCLK clkbuf_4_3_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _18333_/CLK sky130_fd_sc_hd__clkbuf_16
Xrebuffer3 _13089_/B vssd1 vssd1 vccd1 vccd1 _13167_/C1 sky130_fd_sc_hd__dlygate4sd1_1
XANTENNA_clkbuf_1_0_0_HCLK_A clkbuf_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11927__B1 _11926_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16155_ _18118_/Q vssd1 vssd1 vccd1 vccd1 _16155_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13367_ _20112_/Q _13428_/A _13366_/Y _18864_/Q vssd1 vssd1 vccd1 vccd1 _13367_/X
+ sky130_fd_sc_hd__o22a_1
X_10579_ _10933_/A _10579_/B vssd1 vssd1 vccd1 vccd1 _15297_/B sky130_fd_sc_hd__nand2_1
X_15106_ _18526_/D vssd1 vssd1 vccd1 vccd1 _15762_/B sky130_fd_sc_hd__inv_2
X_12318_ _12334_/A vssd1 vssd1 vccd1 vccd1 _12318_/X sky130_fd_sc_hd__buf_1
XFILLER_154_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16086_ _18165_/Q vssd1 vssd1 vccd1 vccd1 _16086_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13298_ _18752_/Q _13297_/X _18752_/Q _13297_/X vssd1 vssd1 vccd1 vccd1 _13299_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_244_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19914_ _19971_/CLK _19914_/D repeater191/X vssd1 vssd1 vccd1 vccd1 _19914_/Q sky130_fd_sc_hd__dfrtp_1
X_15037_ _15037_/A vssd1 vssd1 vccd1 vccd1 _15037_/X sky130_fd_sc_hd__clkbuf_2
X_12249_ _12249_/A vssd1 vssd1 vccd1 vccd1 _12556_/A sky130_fd_sc_hd__inv_2
XFILLER_69_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_158_HCLK clkbuf_4_0_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19435_/CLK sky130_fd_sc_hd__clkbuf_16
X_19845_ _19846_/CLK _19845_/D repeater270/X vssd1 vssd1 vccd1 vccd1 _19845_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_122_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10902__A1 _19686_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17291__A0 _17473_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19776_ _20049_/CLK _19776_/D repeater190/X vssd1 vssd1 vccd1 vccd1 _19776_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_56_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_209_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16988_ _16987_/X _11338_/Y _17493_/S vssd1 vssd1 vccd1 vccd1 _16988_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09054__A hold277/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18727_ _18727_/CLK _18727_/D repeater253/X vssd1 vssd1 vccd1 vccd1 _18727_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_110_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15939_ _18243_/Q _16344_/B vssd1 vssd1 vccd1 vccd1 _15939_/Y sky130_fd_sc_hd__nand2_1
XFILLER_225_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_209_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09460_ _19389_/Q vssd1 vssd1 vccd1 vccd1 _09460_/Y sky130_fd_sc_hd__inv_2
XFILLER_52_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_225_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18658_ _20048_/CLK _18658_/D repeater210/X vssd1 vssd1 vccd1 vccd1 _18658_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_92_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_224_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17609_ _10733_/A _11655_/B _19545_/Q vssd1 vssd1 vccd1 vccd1 _17609_/X sky130_fd_sc_hd__mux2_1
X_09391_ _19396_/Q vssd1 vssd1 vccd1 vccd1 _09391_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18589_ _19437_/CLK _18589_/D repeater269/X vssd1 vssd1 vccd1 vccd1 _18589_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_212_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_178_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16149__A2 _16148_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19338__RESET_B repeater245/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16554__C1 _16553_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_177_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17210__S _17459_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09036__B1 hold305/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16857__A0 _15963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12343__B1 _12107_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13693__B _15169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18902__RESET_B repeater245/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_247_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09727_ _09716_/X _09727_/B _09727_/C _09727_/D vssd1 vssd1 vccd1 vccd1 _09728_/D
+ sky130_fd_sc_hd__and4b_1
XFILLER_83_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09658_ _19988_/Q vssd1 vssd1 vccd1 vccd1 _09744_/A sky130_fd_sc_hd__inv_2
XANTENNA_hold346_A hold346/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_243_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09589_ _09589_/A vssd1 vssd1 vccd1 vccd1 _09589_/Y sky130_fd_sc_hd__inv_2
XPHY_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_243_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11620_ _11620_/A _11637_/A vssd1 vssd1 vccd1 vccd1 _11635_/A sky130_fd_sc_hd__or2_2
XPHY_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09275__B1 _09094_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17337__A1 _11328_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_39_HCLK clkbuf_opt_1_HCLK/A vssd1 vssd1 vccd1 vccd1 _19810_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_144_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09814__A2 _09807_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_230_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_211_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11551_ _11625_/A _11624_/A _11551_/C _11626_/A vssd1 vssd1 vccd1 vccd1 _11552_/D
+ sky130_fd_sc_hd__or4_4
XPHY_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17120__S _17513_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10502_ _19533_/Q _10502_/B _10508_/C _10514_/D vssd1 vssd1 vccd1 vccd1 _11649_/A
+ sky130_fd_sc_hd__nor4_2
XANTENNA__19008__RESET_B hold346/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_90_HCLK_A clkbuf_4_12_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14270_ _14270_/A _14270_/B _15192_/A vssd1 vssd1 vccd1 vccd1 _14784_/C sky130_fd_sc_hd__or3_4
XANTENNA_rebuffer37_A _19418_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11482_ _11482_/A _11482_/B vssd1 vssd1 vccd1 vccd1 _11500_/A sky130_fd_sc_hd__or2_1
XPHY_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13221_ _18534_/Q _13221_/B vssd1 vssd1 vccd1 vccd1 _13222_/B sky130_fd_sc_hd__or2_1
XFILLER_7_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10433_ _10450_/A vssd1 vssd1 vccd1 vccd1 _10433_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__16848__A0 _15768_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12582__B1 _12410_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13152_ _19164_/Q vssd1 vssd1 vccd1 vccd1 _13152_/Y sky130_fd_sc_hd__inv_2
X_10364_ _19859_/Q _10364_/B vssd1 vssd1 vccd1 vccd1 _10364_/X sky130_fd_sc_hd__or2_1
XFILLER_98_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12103_ _19312_/Q _12094_/X _12102_/X _12096_/X vssd1 vssd1 vccd1 vccd1 _19312_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_88_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17960_ _20079_/CLK _17960_/D vssd1 vssd1 vccd1 vccd1 _17960_/Q sky130_fd_sc_hd__dfxtp_1
X_13083_ _13083_/A _13083_/B vssd1 vssd1 vccd1 vccd1 _13172_/A sky130_fd_sc_hd__or2_1
XFILLER_3_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10295_ _18589_/Q _18588_/Q vssd1 vssd1 vccd1 vccd1 _15584_/A sky130_fd_sc_hd__or2_2
XFILLER_88_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_239_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16911_ _16910_/X _09681_/Y _17523_/S vssd1 vssd1 vccd1 vccd1 _16911_/X sky130_fd_sc_hd__mux2_1
X_12034_ _12043_/A vssd1 vssd1 vccd1 vccd1 _12034_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_239_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17891_ _16011_/Y _16012_/Y _16013_/Y _16014_/Y _17913_/S0 _19632_/Q vssd1 vssd1
+ vccd1 vccd1 _17891_/X sky130_fd_sc_hd__mux4_2
XANTENNA__17273__A0 _15768_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16076__A1 _15749_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_238_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19630_ _19630_/CLK _19630_/D repeater257/X vssd1 vssd1 vccd1 vccd1 _19630_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__10896__B1 _10877_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16842_ _15768_/Y _11208_/Y _17546_/S vssd1 vssd1 vccd1 vccd1 _16842_/X sky130_fd_sc_hd__mux2_1
XFILLER_66_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19561_ _19561_/CLK _19561_/D repeater269/X vssd1 vssd1 vccd1 vccd1 _19561_/Q sky130_fd_sc_hd__dfrtp_1
X_16773_ _16772_/X _13399_/Y _17385_/S vssd1 vssd1 vccd1 vccd1 _16773_/X sky130_fd_sc_hd__mux2_1
X_13985_ _18689_/Q vssd1 vssd1 vccd1 vccd1 _14019_/A sky130_fd_sc_hd__inv_2
XFILLER_92_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18512_ _18633_/CLK _18512_/D repeater225/X vssd1 vssd1 vccd1 vccd1 _18512_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_19_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19849__RESET_B repeater258/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12936_ _19263_/Q vssd1 vssd1 vccd1 vccd1 _12936_/Y sky130_fd_sc_hd__inv_2
X_15724_ _15724_/A _15725_/B vssd1 vssd1 vccd1 vccd1 _18657_/D sky130_fd_sc_hd__nor2_1
XFILLER_34_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19492_ _19859_/CLK hold132/X repeater262/X vssd1 vssd1 vccd1 vccd1 _19492_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_46_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16379__A2 _15867_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18443_ _19873_/CLK _18443_/D vssd1 vssd1 vccd1 vccd1 _18443_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_233_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15655_ _15668_/B vssd1 vssd1 vccd1 vccd1 _15661_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_61_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12867_ _18927_/Q vssd1 vssd1 vccd1 vccd1 _13006_/A sky130_fd_sc_hd__inv_2
XPHY_4170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18028__CLK _19510_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14606_ _14751_/A vssd1 vssd1 vccd1 vccd1 _14606_/X sky130_fd_sc_hd__buf_2
X_11818_ _19448_/Q _11814_/X _09077_/X _11815_/X vssd1 vssd1 vccd1 vccd1 _19448_/D
+ sky130_fd_sc_hd__a22o_1
X_18374_ _18441_/CLK _18374_/D vssd1 vssd1 vccd1 vccd1 _18374_/Q sky130_fd_sc_hd__dfxtp_1
X_15586_ _15610_/A _15586_/B vssd1 vssd1 vccd1 vccd1 _15586_/Y sky130_fd_sc_hd__nor2_1
X_12798_ _19252_/Q vssd1 vssd1 vccd1 vccd1 _12798_/Y sky130_fd_sc_hd__inv_2
XPHY_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17325_ _17324_/X _09381_/Y _17529_/S vssd1 vssd1 vccd1 vccd1 _17325_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14537_ _14751_/A vssd1 vssd1 vccd1 vccd1 _14537_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_239_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_187_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11749_ hold142/X _10948_/X _19491_/Q _10951_/X vssd1 vssd1 vccd1 vccd1 hold144/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_175_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16000__A1 _17494_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17030__S _17545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16000__B2 _15999_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17256_ _17255_/X _15642_/A _17318_/S vssd1 vssd1 vccd1 vccd1 _17256_/X sky130_fd_sc_hd__mux2_1
X_14468_ _18359_/Q _14463_/X _14443_/X _14465_/X vssd1 vssd1 vccd1 vccd1 _18359_/D
+ sky130_fd_sc_hd__a22o_1
X_13419_ _13419_/A vssd1 vssd1 vccd1 vccd1 _13528_/B sky130_fd_sc_hd__inv_2
X_16207_ _16721_/B vssd1 vssd1 vccd1 vccd1 _16212_/B sky130_fd_sc_hd__buf_4
XFILLER_146_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17187_ _17186_/X _13851_/Y _17545_/S vssd1 vssd1 vccd1 vccd1 _17187_/X sky130_fd_sc_hd__mux2_1
X_14399_ _18399_/Q _14394_/X _14359_/X _14396_/X vssd1 vssd1 vccd1 vccd1 _18399_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_128_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12573__B1 _12394_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16138_ _16136_/Y _16053_/X _16137_/Y _16055_/X vssd1 vssd1 vccd1 vccd1 _16138_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09049__A hold310/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08960_ _10322_/A _18776_/Q _19856_/Q _08959_/Y vssd1 vssd1 vccd1 vccd1 _08960_/X
+ sky130_fd_sc_hd__o22a_1
X_16069_ _16634_/A vssd1 vssd1 vccd1 vccd1 _16069_/X sky130_fd_sc_hd__buf_1
XANTENNA__12325__B1 _12078_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17264__A0 _15963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10887__B1 _10861_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19828_ _19846_/CLK _19828_/D repeater270/X vssd1 vssd1 vccd1 vccd1 _19828_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_204_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19759_ _19772_/CLK _19759_/D repeater228/X vssd1 vssd1 vccd1 vccd1 _19759_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_72_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17205__S _17482_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09512_ _09512_/A _09512_/B _09512_/C _09512_/D vssd1 vssd1 vccd1 vccd1 _09565_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_17_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17567__A1 _11153_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_225_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09443_ _19920_/Q vssd1 vssd1 vccd1 vccd1 _10036_/A sky130_fd_sc_hd__inv_2
XFILLER_240_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_225_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09374_ _19392_/Q vssd1 vssd1 vccd1 vccd1 _09374_/Y sky130_fd_sc_hd__inv_4
XFILLER_33_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_221_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10811__B1 _19732_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20077__RESET_B repeater196/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12564__B1 _12375_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_245_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10080_ _10034_/A _10034_/B _10077_/Y _10107_/C vssd1 vssd1 vccd1 vccd1 _19918_/D
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__11936__B _15897_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17255__A0 _17473_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12619__A1 _19021_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_235_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_235_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17007__A0 _17473_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17115__S _17512_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19942__RESET_B repeater244/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13770_ _18741_/Q _18742_/Q _13772_/S vssd1 vssd1 vccd1 vccd1 _18742_/D sky130_fd_sc_hd__mux2_1
X_10982_ _10982_/A vssd1 vssd1 vccd1 vccd1 _19665_/D sky130_fd_sc_hd__inv_2
X_12721_ _14810_/A _12709_/X _12720_/X _12711_/X vssd1 vssd1 vccd1 vccd1 _18956_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_215_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_215_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15440_ _15285_/A _15243_/Y _15263_/Y _15259_/A _15242_/Y vssd1 vssd1 vccd1 vccd1
+ _15441_/B sky130_fd_sc_hd__o32a_1
XPHY_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12652_ _18998_/Q _12650_/X _12599_/X _12651_/X vssd1 vssd1 vccd1 vccd1 _18998_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11603_ _11603_/A vssd1 vssd1 vccd1 vccd1 _11603_/Y sky130_fd_sc_hd__inv_2
XPHY_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15371_ _19787_/Q _10647_/B _10648_/B vssd1 vssd1 vccd1 vccd1 _15371_/X sky130_fd_sc_hd__a21bo_1
XPHY_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12583_ _12598_/A vssd1 vssd1 vccd1 vccd1 _12583_/X sky130_fd_sc_hd__clkbuf_2
XPHY_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14322_ _18440_/Q _14318_/X _14277_/X _14320_/X vssd1 vssd1 vccd1 vccd1 _18440_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17110_ _17109_/X _12905_/Y _17487_/S vssd1 vssd1 vccd1 vccd1 _17110_/X sky130_fd_sc_hd__mux2_1
XPHY_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11534_ _11465_/A _11465_/B _11523_/X _11532_/Y vssd1 vssd1 vccd1 vccd1 _19584_/D
+ sky130_fd_sc_hd__a211oi_2
X_18090_ _18260_/CLK _18090_/D vssd1 vssd1 vccd1 vccd1 _18090_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17041_ _17040_/X _11386_/Y _17548_/S vssd1 vssd1 vccd1 vccd1 _17041_/X sky130_fd_sc_hd__mux2_1
XPHY_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14253_ _18475_/Q _14250_/X _13680_/X _14252_/X vssd1 vssd1 vccd1 vccd1 _18475_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_183_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11465_ _11465_/A _11465_/B vssd1 vssd1 vccd1 vccd1 _11532_/A sky130_fd_sc_hd__or2_1
XFILLER_143_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13204_ _13204_/A vssd1 vssd1 vccd1 vccd1 _13204_/Y sky130_fd_sc_hd__inv_2
X_10416_ _14681_/A _16434_/B vssd1 vssd1 vccd1 vccd1 _10419_/A sky130_fd_sc_hd__or2_1
XANTENNA__18824__RESET_B repeater217/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14184_ _14184_/A _14184_/B _14184_/C _14184_/D vssd1 vssd1 vccd1 vccd1 _14184_/X
+ sky130_fd_sc_hd__and4_1
X_11396_ _19134_/Q vssd1 vssd1 vccd1 vccd1 _11396_/Y sky130_fd_sc_hd__inv_2
XFILLER_180_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13135_ _19158_/Q vssd1 vssd1 vccd1 vccd1 _13135_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10347_ _10347_/A vssd1 vssd1 vccd1 vccd1 _19864_/D sky130_fd_sc_hd__inv_2
X_18992_ _19608_/CLK _18992_/D hold355/X vssd1 vssd1 vccd1 vccd1 _18992_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_98_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12307__B1 _12238_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17943_ _18465_/CLK _17943_/D vssd1 vssd1 vccd1 vccd1 _17943_/Q sky130_fd_sc_hd__dfxtp_1
X_13066_ _13066_/A _13066_/B vssd1 vssd1 vccd1 vccd1 _13204_/A sky130_fd_sc_hd__or2_1
XANTENNA__11846__B _15774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10278_ _14334_/A _14316_/B vssd1 vssd1 vccd1 vccd1 _14301_/B sky130_fd_sc_hd__or2_2
X_12017_ _12017_/A vssd1 vssd1 vccd1 vccd1 _12017_/X sky130_fd_sc_hd__buf_1
XANTENNA__10869__B1 _10868_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater207 repeater208/X vssd1 vssd1 vccd1 vccd1 repeater207/X sky130_fd_sc_hd__buf_8
Xrepeater218 repeater219/X vssd1 vssd1 vccd1 vccd1 repeater218/X sky130_fd_sc_hd__buf_6
X_17874_ _17870_/X _17871_/X _17872_/X _17873_/X _19633_/Q _19634_/Q vssd1 vssd1 vccd1
+ vccd1 _17874_/X sky130_fd_sc_hd__mux4_2
Xrepeater229 repeater230/X vssd1 vssd1 vccd1 vccd1 repeater229/X sky130_fd_sc_hd__buf_6
XFILLER_239_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19613_ _20006_/CLK _19613_/D repeater191/X vssd1 vssd1 vccd1 vccd1 _19613_/Q sky130_fd_sc_hd__dfrtp_1
X_16825_ _17473_/A0 _09935_/Y _17522_/S vssd1 vssd1 vccd1 vccd1 _16825_/X sky130_fd_sc_hd__mux2_1
XFILLER_241_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17892__S1 _19632_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17025__S _17413_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19544_ _19544_/CLK _19544_/D repeater221/X vssd1 vssd1 vccd1 vccd1 _19544_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__19683__RESET_B repeater219/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16756_ vssd1 vssd1 vccd1 vccd1 _16756_/HI _16756_/LO sky130_fd_sc_hd__conb_1
X_13968_ _13802_/B _13967_/A _18706_/Q _13970_/A _13901_/X vssd1 vssd1 vccd1 vccd1
+ _18706_/D sky130_fd_sc_hd__o221a_1
X_15707_ _18788_/Q _11861_/B _13630_/A _15233_/B vssd1 vssd1 vccd1 vccd1 _18641_/D
+ sky130_fd_sc_hd__o31a_4
XFILLER_46_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_222_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19475_ _19515_/CLK hold198/X repeater259/X vssd1 vssd1 vccd1 vccd1 _19475_/Q sky130_fd_sc_hd__dfrtp_1
X_12919_ _19271_/Q vssd1 vssd1 vccd1 vccd1 _12919_/Y sky130_fd_sc_hd__inv_2
XFILLER_234_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16687_ _16687_/A vssd1 vssd1 vccd1 vccd1 _16687_/X sky130_fd_sc_hd__buf_1
X_13899_ _13899_/A vssd1 vssd1 vccd1 vccd1 _14003_/B sky130_fd_sc_hd__inv_2
XANTENNA__16864__S _17522_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18426_ _19873_/CLK _18426_/D vssd1 vssd1 vccd1 vccd1 _18426_/Q sky130_fd_sc_hd__dfxtp_1
X_15638_ _15642_/B _15637_/X _15614_/X vssd1 vssd1 vccd1 vccd1 _15638_/X sky130_fd_sc_hd__o21a_1
XFILLER_62_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_210_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18357_ _19849_/CLK _18357_/D vssd1 vssd1 vccd1 vccd1 _18357_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_203_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15569_ _18586_/Q vssd1 vssd1 vccd1 vccd1 _15569_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17308_ _16484_/X _10198_/Y _17566_/S vssd1 vssd1 vccd1 vccd1 _17308_/X sky130_fd_sc_hd__mux2_1
XFILLER_119_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09090_ _10451_/A vssd1 vssd1 vccd1 vccd1 _09090_/X sky130_fd_sc_hd__buf_4
X_18288_ _18431_/CLK _18288_/D vssd1 vssd1 vccd1 vccd1 _18288_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__19939__CLK _19976_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17695__S _17696_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17239_ _17238_/X _11304_/Y _17493_/S vssd1 vssd1 vccd1 vccd1 _17239_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12546__B1 _17614_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09992_ _09992_/A vssd1 vssd1 vccd1 vccd1 _09992_/Y sky130_fd_sc_hd__inv_2
XFILLER_130_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08943_ _08935_/X _08943_/B _08943_/C _08943_/D vssd1 vssd1 vccd1 vccd1 _08970_/C
+ sky130_fd_sc_hd__and4b_1
XANTENNA__10660__B _18508_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_215_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_229_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17883__S1 _19632_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11772__A _11772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14471__B1 _14419_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_3_0_HCLK_A clkbuf_2_3_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19353__RESET_B hold371/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16774__S _17386_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_212_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09426_ _19397_/Q vssd1 vssd1 vccd1 vccd1 _09426_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13026__A1 _13021_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_212_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_240_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09357_ _20020_/Q vssd1 vssd1 vccd1 vccd1 _09480_/A sky130_fd_sc_hd__inv_2
XFILLER_40_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09288_ _20049_/Q _09285_/X _09077_/X _09287_/X vssd1 vssd1 vccd1 vccd1 _20049_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_hold211_A HTRANS[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold309_A HWDATA[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_193_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12537__B1 _12536_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11250_ _19008_/Q vssd1 vssd1 vccd1 vccd1 _11250_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_181_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10201_ _19657_/Q vssd1 vssd1 vccd1 vccd1 _10957_/A sky130_fd_sc_hd__inv_2
XANTENNA__15419__A _15419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11181_ _17707_/X _11176_/X _19624_/Q _11178_/X vssd1 vssd1 vccd1 vccd1 _19624_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_69_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10132_ _20123_/Q _10132_/B vssd1 vssd1 vccd1 vccd1 _13283_/C sky130_fd_sc_hd__nor2_2
XFILLER_122_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16949__S _16950_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17228__A0 _17486_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_9_HCLK_A clkbuf_4_2_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10063_ _19929_/Q _10062_/Y _10057_/X _10046_/B vssd1 vssd1 vccd1 vccd1 _19929_/D
+ sky130_fd_sc_hd__o211a_1
X_14940_ _14940_/A vssd1 vssd1 vccd1 vccd1 _14941_/A sky130_fd_sc_hd__inv_2
XANTENNA__10315__A2 _10314_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09181__A2 _09164_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14871_ _14872_/A vssd1 vssd1 vccd1 vccd1 _14871_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__17874__S1 _19634_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16610_ _16853_/X _16394_/X _16859_/X _15898_/X vssd1 vssd1 vccd1 vccd1 _16610_/X
+ sky130_fd_sc_hd__o22a_2
X_13822_ _13910_/C _13932_/A vssd1 vssd1 vccd1 vccd1 _13823_/B sky130_fd_sc_hd__or2_2
X_17590_ _15357_/X _19713_/Q _17600_/S vssd1 vssd1 vccd1 vccd1 _17590_/X sky130_fd_sc_hd__mux2_1
XFILLER_91_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19094__RESET_B hold359/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_232_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16541_ _15199_/A _16536_/X _16538_/X _16540_/X vssd1 vssd1 vccd1 vccd1 _16541_/Y
+ sky130_fd_sc_hd__o211ai_4
X_13753_ _18745_/Q _13753_/B vssd1 vssd1 vccd1 vccd1 _13753_/Y sky130_fd_sc_hd__nand2_1
XFILLER_44_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10965_ _10965_/A _10979_/A vssd1 vssd1 vccd1 vccd1 _10975_/A sky130_fd_sc_hd__or2_1
XFILLER_141_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_189_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12704_ _18962_/Q _12698_/X _12538_/X _12699_/X vssd1 vssd1 vccd1 vccd1 _18962_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_16_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19260_ _20013_/CLK _19260_/D repeater241/X vssd1 vssd1 vccd1 vccd1 _19260_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_31_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13684_ _16434_/B _15169_/A vssd1 vssd1 vccd1 vccd1 _13686_/A sky130_fd_sc_hd__or2_1
X_16472_ _16472_/A _16544_/B vssd1 vssd1 vccd1 vccd1 _16472_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__18836__CLK _19900_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10896_ _19692_/Q _10893_/X _10877_/X _10895_/X vssd1 vssd1 vccd1 vccd1 _19692_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_43_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08991__A _19517_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_231_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18211_ _18333_/CLK _18211_/D vssd1 vssd1 vccd1 vccd1 _18211_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_231_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15423_ _19614_/Q _11159_/B _11160_/B vssd1 vssd1 vccd1 vccd1 _15423_/X sky130_fd_sc_hd__a21bo_1
XPHY_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12635_ _19009_/Q _12629_/X _12410_/X _12630_/X vssd1 vssd1 vccd1 vccd1 _19009_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_169_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19191_ _20035_/CLK _19191_/D repeater242/X vssd1 vssd1 vccd1 vccd1 _19191_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_197_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_repeater166_A _17543_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15354_ _15358_/A _17592_/X vssd1 vssd1 vccd1 vccd1 _18498_/D sky130_fd_sc_hd__and2_1
X_18142_ _18142_/CLK _18142_/D vssd1 vssd1 vccd1 vccd1 _18142_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12566_ _19054_/Q _12560_/X _12382_/X _12563_/X vssd1 vssd1 vccd1 vccd1 _19054_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17703__A1 _19757_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11517_ _11517_/A vssd1 vssd1 vccd1 vccd1 _11517_/Y sky130_fd_sc_hd__inv_2
X_14305_ _14305_/A vssd1 vssd1 vccd1 vccd1 _14305_/X sky130_fd_sc_hd__clkbuf_2
XPHY_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15285_ _15285_/A _15285_/B vssd1 vssd1 vccd1 vccd1 _15443_/B sky130_fd_sc_hd__or2_1
XFILLER_157_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18073_ _18169_/CLK _18073_/D vssd1 vssd1 vccd1 vccd1 _18073_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12497_ _19088_/Q _12489_/X _12386_/X _12492_/X vssd1 vssd1 vccd1 vccd1 _19088_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_7_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14236_ _14236_/A vssd1 vssd1 vccd1 vccd1 _14236_/X sky130_fd_sc_hd__clkbuf_2
Xhold209 hold209/A vssd1 vssd1 vccd1 vccd1 hold209/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_output95_A _16678_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17024_ _17023_/X _13082_/A _17542_/S vssd1 vssd1 vccd1 vccd1 _17024_/X sky130_fd_sc_hd__mux2_2
X_11448_ _19574_/Q _11446_/Y _11621_/A _19131_/Q vssd1 vssd1 vccd1 vccd1 _11448_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_160_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14167_ _19114_/Q vssd1 vssd1 vccd1 vccd1 _14167_/Y sky130_fd_sc_hd__inv_2
X_11379_ _19133_/Q vssd1 vssd1 vccd1 vccd1 _11379_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13118_ _19177_/Q vssd1 vssd1 vccd1 vccd1 _13118_/Y sky130_fd_sc_hd__inv_2
XFILLER_3_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18975_ _19576_/CLK _18975_/D repeater282/X vssd1 vssd1 vccd1 vccd1 _18975_/Q sky130_fd_sc_hd__dfrtp_1
X_14098_ _14116_/A vssd1 vssd1 vccd1 vccd1 _14118_/A sky130_fd_sc_hd__inv_2
XANTENNA__16859__S _17482_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17219__A0 _15963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14150__C1 _14112_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17926_ _19814_/CLK _19814_/Q vssd1 vssd1 vccd1 vccd1 _17926_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__19864__RESET_B repeater267/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13049_ _18897_/Q vssd1 vssd1 vccd1 vccd1 _13069_/A sky130_fd_sc_hd__inv_2
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12700__B1 _12599_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17857_ _16283_/Y _16284_/Y _16285_/Y _16286_/Y _17908_/S0 _18759_/Q vssd1 vssd1
+ vccd1 vccd1 _17857_/X sky130_fd_sc_hd__mux4_1
XANTENNA__17865__S1 _18759_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_226_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16808_ _16807_/X _13366_/Y _17535_/S vssd1 vssd1 vccd1 vccd1 _16808_/X sky130_fd_sc_hd__mux2_1
XFILLER_93_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_226_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17788_ _18294_/Q _18286_/Q _18278_/Q _18446_/Q _17923_/S0 _19646_/Q vssd1 vssd1
+ vccd1 vccd1 _17788_/X sky130_fd_sc_hd__mux4_2
XFILLER_53_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19527_ _19771_/CLK _19527_/D repeater189/X vssd1 vssd1 vccd1 vccd1 _19527_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_53_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16739_ _16834_/X _16493_/A _16881_/X _16512_/A vssd1 vssd1 vccd1 vccd1 _16739_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_35_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15999__A _15999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19458_ _19462_/CLK _19458_/D repeater272/X vssd1 vssd1 vccd1 vccd1 _19458_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__16607__B _16607_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09211_ _09211_/A vssd1 vssd1 vccd1 vccd1 _09212_/B sky130_fd_sc_hd__inv_2
XFILLER_50_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18409_ _18473_/CLK _18409_/D vssd1 vssd1 vccd1 vccd1 _18409_/Q sky130_fd_sc_hd__dfxtp_1
X_19389_ _20091_/CLK _19389_/D repeater235/X vssd1 vssd1 vccd1 vccd1 _19389_/Q sky130_fd_sc_hd__dfrtp_1
X_09142_ _15322_/B _09141_/Y _15321_/A _09140_/Y vssd1 vssd1 vccd1 vccd1 _20087_/D
+ sky130_fd_sc_hd__o22a_1
X_09073_ _20102_/Q _09069_/X _09071_/X _09072_/X vssd1 vssd1 vccd1 vccd1 _20102_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__15705__B1 _15673_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17458__A0 _15768_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09975_ _09975_/A vssd1 vssd1 vccd1 vccd1 _09975_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16769__S _17546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08926_ _08921_/X _18773_/Q _19865_/Q _08922_/Y _08925_/X vssd1 vssd1 vccd1 vccd1
+ _08970_/A sky130_fd_sc_hd__o221a_1
XANTENNA__14141__C1 _14106_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20095_ _20107_/CLK _20095_/D repeater234/X vssd1 vssd1 vccd1 vccd1 _20095_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__14692__B1 _14691_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19534__RESET_B repeater221/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12598__A _12598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17856__S1 _18759_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18859__CLK _18866_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_214_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10750_ _19757_/Q _10742_/A _10425_/X _10743_/A vssd1 vssd1 vccd1 vccd1 _19757_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_26_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_198_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09409_ _19935_/Q _19395_/Q _19935_/Q _19395_/Q vssd1 vssd1 vccd1 vccd1 _09416_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_41_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_186_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_201_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10681_ _17742_/X _10676_/X _19783_/Q _10677_/X vssd1 vssd1 vccd1 vccd1 _19783_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_9_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_240_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12420_ _12427_/A vssd1 vssd1 vccd1 vccd1 _12420_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__18642__SET_B repeater219/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_224_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12351_ _19170_/Q _12341_/X hold270/X _12342_/X vssd1 vssd1 vccd1 vccd1 _19170_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_181_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11302_ _11487_/A _18989_/Q _19602_/Q _11301_/Y vssd1 vssd1 vccd1 vccd1 _11302_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17792__S0 _17923_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10784__A2 _19741_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15070_ _15070_/A _19643_/Q _15070_/C vssd1 vssd1 vccd1 vccd1 _15072_/A sky130_fd_sc_hd__or3_4
X_12282_ _19210_/Q _12276_/X _12104_/X _12277_/X vssd1 vssd1 vccd1 vccd1 _19210_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_153_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17449__A0 _15963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14021_ _14021_/A _14120_/A vssd1 vssd1 vccd1 vccd1 _14022_/B sky130_fd_sc_hd__or2_2
X_11233_ _19581_/Q vssd1 vssd1 vccd1 vccd1 _11462_/A sky130_fd_sc_hd__inv_2
XFILLER_107_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_145_HCLK_A clkbuf_4_1_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11164_ _19619_/Q _11164_/B vssd1 vssd1 vccd1 vccd1 _11165_/B sky130_fd_sc_hd__or2_1
XFILLER_95_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19634__CLK _19851_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10115_ _18562_/Q _15466_/A vssd1 vssd1 vccd1 vccd1 _15470_/A sky130_fd_sc_hd__or2_1
XFILLER_110_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18760_ _18765_/CLK _18760_/D repeater196/X vssd1 vssd1 vccd1 vccd1 _18760_/Q sky130_fd_sc_hd__dfrtp_2
X_15972_ _19694_/Q vssd1 vssd1 vccd1 vccd1 _15972_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11095_ _14378_/B _11064_/B _14489_/B _19631_/Q _11094_/Y vssd1 vssd1 vccd1 vccd1
+ _11103_/B sky130_fd_sc_hd__a221o_1
XFILLER_96_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17711_ _15429_/X _19766_/Q _18546_/D vssd1 vssd1 vccd1 vccd1 _17711_/X sky130_fd_sc_hd__mux2_1
X_10046_ _10046_/A _10046_/B vssd1 vssd1 vccd1 vccd1 _10059_/A sky130_fd_sc_hd__or2_2
X_14923_ _14923_/A vssd1 vssd1 vccd1 vccd1 _14923_/X sky130_fd_sc_hd__clkbuf_2
X_18691_ _18701_/CLK _18691_/D hold359/X vssd1 vssd1 vccd1 vccd1 _18691_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA_output133_A _20038_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17847__S1 _18759_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_208_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17642_ _15671_/X _19047_/Q _17655_/S vssd1 vssd1 vccd1 vccd1 _18610_/D sky130_fd_sc_hd__mux2_1
XFILLER_91_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14854_ _18139_/Q _14846_/A _14816_/X _14847_/A vssd1 vssd1 vccd1 vccd1 _18139_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_35_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13805_ _18709_/Q vssd1 vssd1 vccd1 vccd1 _13946_/A sky130_fd_sc_hd__inv_2
X_17573_ _15414_/X _19770_/Q _17584_/S vssd1 vssd1 vccd1 vccd1 _17573_/X sky130_fd_sc_hd__mux2_1
XANTENNA__20109__RESET_B repeater217/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14785_ _14786_/A vssd1 vssd1 vccd1 vccd1 _14785_/X sky130_fd_sc_hd__clkbuf_2
X_11997_ _12187_/B vssd1 vssd1 vccd1 vccd1 _15769_/A sky130_fd_sc_hd__buf_2
XANTENNA__16708__A _19429_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19312_ _19314_/CLK _19312_/D repeater214/X vssd1 vssd1 vccd1 vccd1 _19312_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__17303__S _17523_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16524_ _16504_/X _16519_/X _16521_/X _16523_/X vssd1 vssd1 vccd1 vccd1 _16524_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_16_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10948_ _11771_/A vssd1 vssd1 vccd1 vccd1 _10948_/X sky130_fd_sc_hd__clkbuf_2
X_13736_ _17764_/X vssd1 vssd1 vccd1 vccd1 _13737_/A sky130_fd_sc_hd__inv_2
XFILLER_232_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_232_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19243_ _19314_/CLK _19243_/D repeater237/X vssd1 vssd1 vccd1 vccd1 _19243_/Q sky130_fd_sc_hd__dfrtp_4
X_16455_ _16453_/Y _15831_/A _16454_/Y _15976_/X vssd1 vssd1 vccd1 vccd1 _16455_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_204_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10879_ _10879_/A vssd1 vssd1 vccd1 vccd1 _10879_/X sky130_fd_sc_hd__clkbuf_2
X_13667_ _18781_/Q _13664_/X hold267/X _13665_/X vssd1 vssd1 vccd1 vccd1 _18781_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13132__A _19170_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15406_ _18535_/Q _13222_/B _13223_/B vssd1 vssd1 vccd1 vccd1 _15406_/X sky130_fd_sc_hd__a21bo_1
XPHY_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12618_ _19022_/Q _12613_/X _12380_/X _12616_/X vssd1 vssd1 vccd1 vccd1 _19022_/D
+ sky130_fd_sc_hd__a22o_1
X_19174_ _19214_/CLK _19174_/D hold367/X vssd1 vssd1 vccd1 vccd1 _19174_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16386_ _15254_/Y _15840_/A _16385_/Y _15842_/X vssd1 vssd1 vccd1 vccd1 _16386_/X
+ sky130_fd_sc_hd__o22a_1
X_13598_ _13598_/A vssd1 vssd1 vccd1 vccd1 _13598_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08968__A2 _08962_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18125_ _18765_/CLK _18125_/D vssd1 vssd1 vccd1 vccd1 _18125_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_247_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15337_ _18491_/Q _18490_/Q _14222_/B vssd1 vssd1 vccd1 vccd1 _15337_/X sky130_fd_sc_hd__a21bo_1
X_12549_ _15222_/A _12247_/B _12556_/B _11086_/A _12548_/Y vssd1 vssd1 vccd1 vccd1
+ _12550_/A sky130_fd_sc_hd__o32a_1
XFILLER_145_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17783__S0 _17923_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18056_ _18169_/CLK _18056_/D vssd1 vssd1 vccd1 vccd1 _18056_/Q sky130_fd_sc_hd__dfxtp_1
X_15268_ _15268_/A _15311_/A _15268_/C vssd1 vssd1 vccd1 vccd1 _15268_/X sky130_fd_sc_hd__or3_4
XANTENNA__15163__B2 _15160_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17007_ _17473_/A0 _16693_/Y _17547_/S vssd1 vssd1 vccd1 vccd1 _17007_/X sky130_fd_sc_hd__mux2_1
X_14219_ _14193_/X _14219_/B _14219_/C _14219_/D vssd1 vssd1 vccd1 vccd1 _14219_/X
+ sky130_fd_sc_hd__and4b_1
X_15199_ _15199_/A vssd1 vssd1 vccd1 vccd1 _17566_/S sky130_fd_sc_hd__clkinv_16
XFILLER_99_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09760_ _20000_/Q _09758_/X _09759_/X _09755_/A vssd1 vssd1 vccd1 vccd1 _20000_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA_clkbuf_leaf_67_HCLK_A clkbuf_opt_3_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18958_ _18959_/CLK _18958_/D repeater257/X vssd1 vssd1 vccd1 vccd1 _18958_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_100_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09145__A2 _17605_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17909_ _17905_/X _17906_/X _17907_/X _17908_/X _18760_/Q _18761_/Q vssd1 vssd1 vccd1
+ vccd1 _17909_/X sky130_fd_sc_hd__mux4_2
X_09691_ _19403_/Q vssd1 vssd1 vccd1 vccd1 _09691_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18889_ _19964_/CLK _18889_/D hold372/X vssd1 vssd1 vccd1 vccd1 _18889_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17838__S1 _18759_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrebuffer13 _13899_/A vssd1 vssd1 vccd1 vccd1 _13903_/A sky130_fd_sc_hd__dlygate4sd1_1
XANTENNA__10160__B1 _09094_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrebuffer24 _14007_/B vssd1 vssd1 vccd1 vccd1 _14146_/C1 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_212_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrebuffer35 _14005_/B vssd1 vssd1 vccd1 vccd1 _14147_/A2 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer46 _13083_/B vssd1 vssd1 vccd1 vccd1 _13174_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_81_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrebuffer57 _19388_/Q vssd1 vssd1 vccd1 vccd1 _09388_/B2 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer68 _14016_/B vssd1 vssd1 vccd1 vccd1 _14130_/C1 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer79 _14032_/B vssd1 vssd1 vccd1 vccd1 _14102_/C1 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17213__S _17523_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_194_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19507__CLK _19510_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18580__RESET_B hold348/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrebuffer103 _10025_/A vssd1 vssd1 vccd1 vccd1 _10053_/A sky130_fd_sc_hd__buf_2
XFILLER_148_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_72_HCLK clkbuf_opt_4_HCLK/A vssd1 vssd1 vccd1 vccd1 _18866_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_194_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09125_ _09154_/A _09149_/A _09144_/C _09125_/D vssd1 vssd1 vccd1 vccd1 _13493_/A
+ sky130_fd_sc_hd__or4_4
Xrebuffer114 _14022_/B vssd1 vssd1 vccd1 vccd1 _14121_/C1 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer125 _13549_/B vssd1 vssd1 vccd1 vccd1 _13576_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_157_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_191_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17774__S0 _19647_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09056_ _20107_/Q _09053_/X hold276/X _09055_/X vssd1 vssd1 vccd1 vccd1 _20107_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_124_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19786__RESET_B repeater203/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_237_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11715__A1 _19516_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11715__B2 _16950_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16654__A1 _17076_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14114__C1 _14135_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09958_ _19966_/Q _09957_/Y _09950_/X _09958_/C1 vssd1 vssd1 vccd1 vccd1 _19966_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_103_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14665__B1 _14567_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20078_ _20079_/CLK _20078_/D repeater205/X vssd1 vssd1 vccd1 vccd1 _20078_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_46_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17829__S1 _18752_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09889_ _19968_/Q _16721_/A _09871_/A _19355_/Q vssd1 vssd1 vccd1 vccd1 _09889_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_57_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11920_ _12234_/A vssd1 vssd1 vccd1 vccd1 _11920_/X sky130_fd_sc_hd__buf_2
XFILLER_246_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12121__A _12121_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11851_ _11851_/A _11867_/A vssd1 vssd1 vccd1 vccd1 _11856_/A sky130_fd_sc_hd__or2_1
XPHY_4544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15090__B1 _14793_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10802_ _19735_/Q _10801_/Y _10793_/B _10797_/A vssd1 vssd1 vccd1 vccd1 _19735_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__17123__S _17545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14570_ _18298_/Q _14559_/A hold320/X _14560_/A vssd1 vssd1 vccd1 vccd1 _18298_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_214_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11782_ _15772_/A _11933_/A vssd1 vssd1 vccd1 vccd1 _11821_/A sky130_fd_sc_hd__or2_4
XPHY_4588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_0_0_HCLK clkbuf_4_1_0_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_0_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XPHY_3865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10733_ _10733_/A vssd1 vssd1 vccd1 vccd1 _10733_/Y sky130_fd_sc_hd__inv_2
XFILLER_214_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13521_ _18765_/Q vssd1 vssd1 vccd1 vccd1 _15145_/A sky130_fd_sc_hd__inv_2
XPHY_3887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_201_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16962__S _17536_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13452_ _13429_/A _13342_/B _13450_/Y _13445_/X vssd1 vssd1 vccd1 vccd1 _18855_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_15_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16240_ _16637_/A vssd1 vssd1 vccd1 vccd1 _16556_/A sky130_fd_sc_hd__inv_2
X_10664_ _17729_/X _10661_/X _19796_/Q _10663_/X vssd1 vssd1 vccd1 vccd1 _19796_/D
+ sky130_fd_sc_hd__a22o_1
X_12403_ _19147_/Q _12400_/X _12401_/X _12402_/X vssd1 vssd1 vccd1 vccd1 _19147_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_40_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13383_ _20098_/Q vssd1 vssd1 vccd1 vccd1 _13383_/Y sky130_fd_sc_hd__inv_2
X_16171_ _19652_/Q _16095_/Y _16024_/Y _16169_/Y vssd1 vssd1 vccd1 vccd1 _16171_/X
+ sky130_fd_sc_hd__a22o_1
X_10595_ _10595_/A _10595_/B _19801_/Q _10595_/D vssd1 vssd1 vccd1 vccd1 _10613_/B
+ sky130_fd_sc_hd__nor4_2
XFILLER_154_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17765__S0 _17923_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12334_ _12334_/A vssd1 vssd1 vccd1 vccd1 _12334_/X sky130_fd_sc_hd__clkbuf_2
X_15122_ _15123_/A vssd1 vssd1 vccd1 vccd1 _15122_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_182_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19930_ _19933_/CLK _19930_/D repeater236/X vssd1 vssd1 vccd1 vccd1 _19930_/Q sky130_fd_sc_hd__dfrtp_1
X_15053_ _18022_/Q _15047_/X _15000_/X _15049_/X vssd1 vssd1 vccd1 vccd1 _18022_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_182_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12265_ _19223_/Q _12260_/X _12074_/X _12263_/X vssd1 vssd1 vccd1 vccd1 _19223_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_141_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14004_ _14004_/A _14148_/A vssd1 vssd1 vccd1 vccd1 _14005_/B sky130_fd_sc_hd__or2_2
XANTENNA_clkbuf_3_6_0_HCLK_A clkbuf_3_7_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11216_ _19601_/Q _11211_/Y _11481_/A _19015_/Q _11215_/X vssd1 vssd1 vccd1 vccd1
+ _11223_/C sky130_fd_sc_hd__o221a_1
XANTENNA__19456__RESET_B repeater272/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19861_ _19867_/CLK _19861_/D repeater263/X vssd1 vssd1 vccd1 vccd1 _19861_/Q sky130_fd_sc_hd__dfrtp_4
X_12196_ _19255_/Q _12189_/X _12078_/X _12192_/X vssd1 vssd1 vccd1 vccd1 _19255_/D
+ sky130_fd_sc_hd__a22o_1
X_18812_ _20115_/CLK _18812_/D repeater238/X vssd1 vssd1 vccd1 vccd1 _18812_/Q sky130_fd_sc_hd__dfrtp_1
Xoutput82 _16533_/Y vssd1 vssd1 vccd1 vccd1 HRDATA[12] sky130_fd_sc_hd__clkbuf_2
Xoutput93 _16656_/X vssd1 vssd1 vccd1 vccd1 HRDATA[22] sky130_fd_sc_hd__clkbuf_2
X_11147_ _11147_/A vssd1 vssd1 vccd1 vccd1 _14598_/B sky130_fd_sc_hd__buf_1
X_19792_ _19794_/CLK _19792_/D repeater219/X vssd1 vssd1 vccd1 vccd1 _19792_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__14511__A hold331/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18743_ _20066_/CLK _18743_/D repeater209/X vssd1 vssd1 vccd1 vccd1 _18743_/Q sky130_fd_sc_hd__dfrtp_1
X_11078_ _18624_/Q vssd1 vssd1 vccd1 vccd1 _15858_/B sky130_fd_sc_hd__inv_2
X_15955_ _18107_/Q vssd1 vssd1 vccd1 vccd1 _15955_/Y sky130_fd_sc_hd__inv_2
X_10029_ _19327_/Q _10029_/B vssd1 vssd1 vccd1 vccd1 _10030_/A sky130_fd_sc_hd__or2_1
XFILLER_37_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14906_ _18106_/Q _14897_/A _14868_/X _14898_/A vssd1 vssd1 vccd1 vccd1 _18106_/D
+ sky130_fd_sc_hd__a22o_1
X_18674_ _18718_/CLK _18674_/D repeater252/X vssd1 vssd1 vccd1 vccd1 _18674_/Q sky130_fd_sc_hd__dfrtp_1
X_15886_ _15882_/Y _15884_/X _15885_/Y _15858_/D vssd1 vssd1 vccd1 vccd1 _15918_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_91_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17625_ _19894_/Q _19747_/Q _17630_/S vssd1 vssd1 vccd1 vccd1 _17625_/X sky130_fd_sc_hd__mux2_1
X_14837_ _18151_/Q _14832_/X _14808_/X _14834_/X vssd1 vssd1 vccd1 vccd1 _18151_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11890__B1 _09039_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15081__B1 _14782_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17033__S _17543_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17556_ _17555_/X _19878_/Q _19498_/Q vssd1 vssd1 vccd1 vccd1 _17556_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12434__A2 _12400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14768_ _18187_/Q _14760_/A _14691_/X _14761_/A vssd1 vssd1 vccd1 vccd1 _18187_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_44_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_95_HCLK clkbuf_4_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19352_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_32_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16507_ _17215_/X _16505_/X _17222_/X _16506_/X vssd1 vssd1 vccd1 vccd1 _16507_/X
+ sky130_fd_sc_hd__o22a_1
X_13719_ _18760_/Q _13710_/B _14857_/A _14642_/A _13706_/B vssd1 vssd1 vccd1 vccd1
+ _13719_/X sky130_fd_sc_hd__a32o_1
XANTENNA__16872__S _17536_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17487_ _17486_/X _12936_/Y _17487_/S vssd1 vssd1 vccd1 vccd1 _17487_/X sky130_fd_sc_hd__mux2_1
XFILLER_204_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14699_ _14699_/A vssd1 vssd1 vccd1 vccd1 _14699_/X sky130_fd_sc_hd__clkbuf_2
X_19226_ _19630_/CLK _19226_/D repeater257/X vssd1 vssd1 vccd1 vccd1 _19226_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_176_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16438_ _19446_/Q vssd1 vssd1 vccd1 vccd1 _16438_/Y sky130_fd_sc_hd__inv_2
XFILLER_176_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13797__A _19125_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_192_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19157_ _19157_/CLK _19157_/D repeater268/X vssd1 vssd1 vccd1 vccd1 _19157_/Q sky130_fd_sc_hd__dfrtp_1
X_16369_ _19445_/Q vssd1 vssd1 vccd1 vccd1 _16369_/Y sky130_fd_sc_hd__inv_2
XFILLER_191_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11945__A1 _19395_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18108_ _18260_/CLK _18108_/D vssd1 vssd1 vccd1 vccd1 _18108_/Q sky130_fd_sc_hd__dfxtp_1
X_19088_ _19609_/CLK _19088_/D hold357/X vssd1 vssd1 vccd1 vccd1 _19088_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_106_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_1_HCLK clkbuf_4_0_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _18169_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_160_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18039_ _19851_/CLK _18039_/D vssd1 vssd1 vccd1 vccd1 _18039_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16620__B _16621_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20001_ _20003_/CLK _20001_/D repeater192/X vssd1 vssd1 vccd1 vccd1 _20001_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17208__S _17414_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19126__RESET_B hold348/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09812_ _09807_/A _09807_/B _09807_/C vssd1 vssd1 vccd1 vccd1 _09813_/B sky130_fd_sc_hd__o21a_1
XFILLER_59_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09743_ _09743_/A _09781_/A vssd1 vssd1 vccd1 vccd1 _09744_/B sky130_fd_sc_hd__or2_2
XFILLER_223_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09674_ _19997_/Q _09673_/Y _09753_/A _19426_/Q vssd1 vssd1 vccd1 vccd1 _09674_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_228_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_227_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_243_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_227_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11881__B1 hold288/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_243_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18761__RESET_B repeater196/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16782__S _17522_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19967__RESET_B repeater274/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09108_ _11926_/A vssd1 vssd1 vccd1 vccd1 _09108_/X sky130_fd_sc_hd__buf_4
XANTENNA__13500__A _18760_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10380_ _10376_/B _10379_/X _10320_/X _10354_/A _10321_/D vssd1 vssd1 vccd1 vccd1
+ _10381_/A sky130_fd_sc_hd__o32a_1
XFILLER_164_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_191_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09039_ hold298/X vssd1 vssd1 vccd1 vccd1 _09039_/X sky130_fd_sc_hd__buf_4
XFILLER_151_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14886__B1 _14802_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12050_ _19332_/Q _12016_/A _11924_/X _12017_/A vssd1 vssd1 vccd1 vccd1 _19332_/D
+ sky130_fd_sc_hd__a22o_1
Xhold370 hold370/A vssd1 vssd1 vccd1 vccd1 hold370/X sky130_fd_sc_hd__dlygate4sd3_1
X_11001_ _11001_/A vssd1 vssd1 vccd1 vccd1 _11002_/B sky130_fd_sc_hd__inv_2
XFILLER_89_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09762__C1 _09759_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17118__S _17542_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_237_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_50_HCLK_A clkbuf_opt_1_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15740_ _18670_/Q _18668_/Q vssd1 vssd1 vccd1 vccd1 _15740_/X sky130_fd_sc_hd__or2_1
XFILLER_19_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18849__RESET_B repeater232/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12952_ _19285_/Q vssd1 vssd1 vccd1 vccd1 _12952_/Y sky130_fd_sc_hd__inv_2
XFILLER_245_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_233_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11903_ _19414_/Q _11898_/X _09064_/X _11899_/X vssd1 vssd1 vccd1 vccd1 _19414_/D
+ sky130_fd_sc_hd__a22o_1
X_15671_ _15669_/Y _15670_/X _15643_/X vssd1 vssd1 vccd1 vccd1 _15671_/X sky130_fd_sc_hd__o21a_1
XPHY_4330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12883_ _12967_/B _12883_/B vssd1 vssd1 vccd1 vccd1 _12978_/A sky130_fd_sc_hd__or2_1
XPHY_4341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17410_ _17409_/X _16120_/Y _17517_/S vssd1 vssd1 vccd1 vccd1 _17410_/X sky130_fd_sc_hd__mux2_1
X_14622_ _18270_/Q _14616_/X _09177_/X _14618_/X vssd1 vssd1 vccd1 vccd1 _18270_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18390_ _18441_/CLK _18390_/D vssd1 vssd1 vccd1 vccd1 _18390_/Q sky130_fd_sc_hd__dfxtp_1
X_11834_ _10147_/X _19438_/Q _11834_/S vssd1 vssd1 vccd1 vccd1 _19438_/D sky130_fd_sc_hd__mux2_1
XPHY_4374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17341_ _16365_/Y _17849_/X _17568_/S vssd1 vssd1 vccd1 vccd1 _17341_/X sky130_fd_sc_hd__mux2_2
X_11765_ _11772_/A vssd1 vssd1 vccd1 vccd1 _11765_/X sky130_fd_sc_hd__clkbuf_2
X_14553_ _18309_/Q _14546_/X hold330/X _14548_/X vssd1 vssd1 vccd1 vccd1 _18309_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_3673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10716_ _10715_/X _19773_/Q _10716_/S vssd1 vssd1 vccd1 vccd1 _19773_/D sky130_fd_sc_hd__mux2_1
XPHY_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13504_ _14628_/A _13511_/A vssd1 vssd1 vccd1 vccd1 _14696_/B sky130_fd_sc_hd__or2_1
XFILLER_158_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17272_ _17271_/X _09858_/A _17488_/S vssd1 vssd1 vccd1 vccd1 _17272_/X sky130_fd_sc_hd__mux2_1
XFILLER_201_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11696_ _19525_/Q _11690_/X _10861_/X _11692_/X vssd1 vssd1 vccd1 vccd1 _19525_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14484_ _18350_/Q _14478_/X _12723_/X _14480_/X vssd1 vssd1 vccd1 vccd1 _18350_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_186_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19011_ _19597_/CLK _19011_/D repeater281/X vssd1 vssd1 vccd1 vccd1 _19011_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__16705__B _16705_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16223_ _16221_/Y _16303_/A _16222_/Y _16055_/A vssd1 vssd1 vccd1 vccd1 _16223_/X
+ sky130_fd_sc_hd__o22a_1
X_13435_ _13435_/A _13489_/C _13435_/C vssd1 vssd1 vccd1 vccd1 _18865_/D sky130_fd_sc_hd__nor3_1
X_10647_ _19787_/Q _10647_/B vssd1 vssd1 vccd1 vccd1 _10648_/B sky130_fd_sc_hd__or2_1
XANTENNA__18623__D _18623_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrebuffer4 _13089_/B vssd1 vssd1 vccd1 vccd1 _13165_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XANTENNA__11927__B2 _11892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13366_ _20118_/Q vssd1 vssd1 vccd1 vccd1 _13366_/Y sky130_fd_sc_hd__inv_2
X_16154_ _18030_/Q vssd1 vssd1 vccd1 vccd1 _16154_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19637__RESET_B repeater258/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10578_ _10592_/B _19803_/Q _19804_/Q vssd1 vssd1 vccd1 vccd1 _10579_/B sky130_fd_sc_hd__or3b_4
XFILLER_6_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19972__CLK _19976_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13129__B1 _19173_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15105_ _17986_/Q _15096_/A _18952_/Q _15097_/A vssd1 vssd1 vccd1 vccd1 _17986_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_142_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12317_ _12361_/A vssd1 vssd1 vccd1 vccd1 _12334_/A sky130_fd_sc_hd__buf_2
X_16085_ _18053_/Q vssd1 vssd1 vccd1 vccd1 _16085_/Y sky130_fd_sc_hd__inv_2
X_13297_ _14819_/A _13293_/X _18756_/Q _13293_/X vssd1 vssd1 vccd1 vccd1 _13297_/X
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__12026__A hold233/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19913_ _19971_/CLK _19913_/D repeater191/X vssd1 vssd1 vccd1 vccd1 _19913_/Q sky130_fd_sc_hd__dfrtp_1
X_15036_ _15036_/A vssd1 vssd1 vccd1 vccd1 _15037_/A sky130_fd_sc_hd__inv_2
X_12248_ _19226_/Q _19225_/Q vssd1 vssd1 vccd1 vccd1 _12249_/A sky130_fd_sc_hd__or2_2
XANTENNA__17028__S _17518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19844_ _19846_/CLK _19844_/D repeater270/X vssd1 vssd1 vccd1 vccd1 _19844_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_123_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_229_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12179_ _19262_/Q _12150_/A _11926_/X _12151_/A vssd1 vssd1 vccd1 vccd1 _19262_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17910__S0 _17913_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19775_ _20049_/CLK _19775_/D repeater190/X vssd1 vssd1 vccd1 vccd1 _19775_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_56_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16867__S _17546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16987_ _15768_/Y _11211_/Y _17546_/S vssd1 vssd1 vccd1 vccd1 _16987_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20124__RESET_B repeater196/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_237_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18726_ _18727_/CLK _18726_/D repeater253/X vssd1 vssd1 vccd1 vccd1 _18726_/Q sky130_fd_sc_hd__dfrtp_1
X_15938_ _16483_/B vssd1 vssd1 vccd1 vccd1 _16344_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_225_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18657_ _20048_/CLK _18657_/D repeater210/X vssd1 vssd1 vccd1 vccd1 _18657_/Q sky130_fd_sc_hd__dfrtp_1
X_15869_ _19192_/Q _15878_/B vssd1 vssd1 vccd1 vccd1 _15869_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__15054__B1 _15002_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_225_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16251__C1 _16250_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17608_ _10531_/B _11655_/B _19545_/Q vssd1 vssd1 vccd1 vccd1 _17608_/X sky130_fd_sc_hd__mux2_1
XANTENNA__15072__A _15072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09390_ _19936_/Q vssd1 vssd1 vccd1 vccd1 _10023_/A sky130_fd_sc_hd__inv_2
X_18588_ _19437_/CLK _18588_/D repeater269/X vssd1 vssd1 vccd1 vccd1 _18588_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_51_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17539_ _17538_/X _15865_/Y _17539_/S vssd1 vssd1 vccd1 vccd1 _17539_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_193_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_177_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16554__B1 _17132_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16615__B _16615_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19209_ _19214_/CLK _19209_/D hold367/X vssd1 vssd1 vccd1 vccd1 _19209_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_193_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09036__A1 _20115_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19378__RESET_B repeater230/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12040__B1 _11909_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14135__B _14135_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_102_HCLK clkbuf_4_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19288_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_99_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14151__A _19122_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17901__S0 _17913_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_219_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16777__S _17414_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09726_ _09741_/A _19414_/Q _19985_/Q _09723_/Y _09725_/X vssd1 vssd1 vccd1 vccd1
+ _09727_/D sky130_fd_sc_hd__o221a_1
XFILLER_67_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_227_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_215_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09657_ _19991_/Q vssd1 vssd1 vccd1 vccd1 _09747_/A sky130_fd_sc_hd__inv_2
XANTENNA__15045__B1 _15020_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16242__C1 _16241_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_243_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09588_ _09484_/A _09484_/B _09584_/Y _09587_/X vssd1 vssd1 vccd1 vccd1 _20024_/D
+ sky130_fd_sc_hd__a211oi_2
XANTENNA_hold241_A HWDATA[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16793__A0 _16792_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold339_A sda_i_S5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17401__S _17565_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11550_ _11623_/A _11622_/A _11621_/A _11639_/A vssd1 vssd1 vccd1 vccd1 _11552_/C
+ sky130_fd_sc_hd__or4_4
XPHY_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10501_ _19542_/Q _19541_/Q _10501_/C _11654_/B vssd1 vssd1 vccd1 vccd1 _10514_/D
+ sky130_fd_sc_hd__or4_4
XPHY_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11481_ _11481_/A _11503_/A vssd1 vssd1 vccd1 vccd1 _11482_/B sky130_fd_sc_hd__or2_2
XPHY_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10854__A _15823_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_183_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14326__A hold331/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13220_ _18533_/Q _13220_/B vssd1 vssd1 vccd1 vccd1 _13221_/B sky130_fd_sc_hd__or2_1
X_10432_ _14681_/A _15199_/A vssd1 vssd1 vccd1 vccd1 _10450_/A sky130_fd_sc_hd__or2_2
XFILLER_171_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12031__B1 _12030_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13151_ _13148_/Y _18908_/Q _13149_/Y _18896_/Q _13150_/X vssd1 vssd1 vccd1 vccd1
+ _13159_/B sky130_fd_sc_hd__o221a_1
X_10363_ _10363_/A vssd1 vssd1 vccd1 vccd1 _19860_/D sky130_fd_sc_hd__inv_2
XFILLER_191_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12102_ hold310/X vssd1 vssd1 vccd1 vccd1 _12102_/X sky130_fd_sc_hd__clkbuf_4
X_13082_ _13082_/A _13175_/A vssd1 vssd1 vccd1 vccd1 _13083_/B sky130_fd_sc_hd__or2_2
X_10294_ _18613_/Q _18612_/Q vssd1 vssd1 vccd1 vccd1 _10310_/C sky130_fd_sc_hd__or2_1
XFILLER_88_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16910_ _17473_/A0 _09912_/Y _17522_/S vssd1 vssd1 vccd1 vccd1 _16910_/X sky130_fd_sc_hd__mux2_1
X_12033_ _19343_/Q _12023_/X _12032_/X _12024_/X vssd1 vssd1 vccd1 vccd1 _19343_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_88_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17890_ _16007_/Y _16008_/Y _16009_/Y _16010_/Y _17913_/S0 _19632_/Q vssd1 vssd1
+ vccd1 vccd1 _17890_/X sky130_fd_sc_hd__mux4_2
XFILLER_104_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_239_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16841_ _16840_/X _15559_/Y _17474_/S vssd1 vssd1 vccd1 vccd1 _16841_/X sky130_fd_sc_hd__mux2_1
XFILLER_144_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19560_ _19561_/CLK _19560_/D repeater269/X vssd1 vssd1 vccd1 vccd1 _19560_/Q sky130_fd_sc_hd__dfrtp_1
X_16772_ _15963_/X _12765_/Y _17534_/S vssd1 vssd1 vccd1 vccd1 _16772_/X sky130_fd_sc_hd__mux2_1
XANTENNA__18683__RESET_B repeater252/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13984_ _18690_/Q vssd1 vssd1 vccd1 vccd1 _14020_/A sky130_fd_sc_hd__inv_2
XANTENNA__08994__A _18620_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18511_ _19780_/CLK _18511_/D repeater226/X vssd1 vssd1 vccd1 vccd1 _18511_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_207_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15723_ _15723_/A _15725_/B vssd1 vssd1 vccd1 vccd1 _18656_/D sky130_fd_sc_hd__nor2_1
X_19491_ _19515_/CLK hold144/X repeater260/X vssd1 vssd1 vccd1 vccd1 _19491_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_37_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12935_ _19265_/Q _12859_/A _12933_/Y _18925_/Q _12934_/X vssd1 vssd1 vccd1 vccd1
+ _12941_/C sky130_fd_sc_hd__o221a_1
XFILLER_18_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_207_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18442_ _19859_/CLK _18442_/D vssd1 vssd1 vccd1 vccd1 _18442_/Q sky130_fd_sc_hd__dfxtp_1
X_15654_ _18607_/Q _15654_/B vssd1 vssd1 vccd1 vccd1 _15668_/B sky130_fd_sc_hd__or2_1
XFILLER_221_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12866_ _18928_/Q vssd1 vssd1 vccd1 vccd1 _13007_/A sky130_fd_sc_hd__clkinv_1
XPHY_4171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14605_ _18280_/Q _14599_/X _14604_/X _14602_/X vssd1 vssd1 vccd1 vccd1 _18280_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18373_ _18441_/CLK _18373_/D vssd1 vssd1 vccd1 vccd1 _18373_/Q sky130_fd_sc_hd__dfxtp_1
X_11817_ _19449_/Q _11814_/X _09075_/X _11815_/X vssd1 vssd1 vccd1 vccd1 _19449_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_199_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15585_ _18590_/Q _15584_/A _15583_/Y _15584_/Y vssd1 vssd1 vccd1 vccd1 _15586_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_199_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12797_ _19227_/Q vssd1 vssd1 vccd1 vccd1 _12797_/Y sky130_fd_sc_hd__inv_2
XPHY_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17324_ _15963_/X _09525_/Y _17534_/S vssd1 vssd1 vccd1 vccd1 _17324_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17311__S _17568_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14536_ _18320_/Q _14530_/X _14535_/X _14533_/X vssd1 vssd1 vccd1 vccd1 _18320_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_175_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11748_ hold130/X _10948_/X _19492_/Q _10951_/X vssd1 vssd1 vccd1 vccd1 hold132/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_239_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17255_ _17473_/A0 _16570_/Y _17547_/S vssd1 vssd1 vccd1 vccd1 _17255_/X sky130_fd_sc_hd__mux2_1
X_14467_ _18360_/Q _14463_/X _14441_/X _14465_/X vssd1 vssd1 vccd1 vccd1 _18360_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14236__A _14236_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11679_ _11671_/X _11672_/Y _18625_/Q _19538_/Q _11666_/X vssd1 vssd1 vccd1 vccd1
+ _19538_/D sky130_fd_sc_hd__a32o_1
X_16206_ _16437_/A _18741_/Q vssd1 vssd1 vccd1 vccd1 _16206_/Y sky130_fd_sc_hd__nand2_1
X_13418_ _13418_/A _13418_/B _13418_/C _13418_/D vssd1 vssd1 vccd1 vccd1 _13419_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__19471__RESET_B repeater260/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12022__B1 _09051_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_125_HCLK clkbuf_4_4_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19041_/CLK sky130_fd_sc_hd__clkbuf_16
X_17186_ _17185_/X _14054_/Y _17544_/S vssd1 vssd1 vccd1 vccd1 _17186_/X sky130_fd_sc_hd__mux2_1
XFILLER_127_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14398_ _18400_/Q _14394_/X _14356_/X _14396_/X vssd1 vssd1 vccd1 vccd1 _18400_/D
+ sky130_fd_sc_hd__a22o_1
X_16137_ _19818_/Q vssd1 vssd1 vccd1 vccd1 _16137_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13349_ _13433_/A _13439_/A vssd1 vssd1 vccd1 vccd1 _13350_/B sky130_fd_sc_hd__or2_2
XFILLER_142_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16068_ _16066_/Y _15884_/X _16067_/Y _15915_/X vssd1 vssd1 vccd1 vccd1 _16068_/X
+ sky130_fd_sc_hd__o22a_1
X_15019_ _18043_/Q _15011_/A _15006_/X _15012_/A vssd1 vssd1 vccd1 vccd1 _18043_/D
+ sky130_fd_sc_hd__a22o_1
X_19827_ _19842_/CLK _19827_/D repeater271/X vssd1 vssd1 vccd1 vccd1 _19827_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_96_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_204_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12089__B1 _12088_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19758_ _19772_/CLK _19758_/D repeater189/X vssd1 vssd1 vccd1 vccd1 _19758_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_84_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_209_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09511_ _09472_/A _19301_/Q _20009_/Q _09508_/Y _09510_/X vssd1 vssd1 vccd1 vccd1
+ _09512_/D sky130_fd_sc_hd__o221a_1
X_18709_ _19224_/CLK _18709_/D repeater186/X vssd1 vssd1 vccd1 vccd1 _18709_/Q sky130_fd_sc_hd__dfrtp_1
X_19689_ _19720_/CLK _19689_/D repeater201/X vssd1 vssd1 vccd1 vccd1 _19689_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__15027__B1 _14996_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09442_ _19378_/Q vssd1 vssd1 vccd1 vccd1 _09442_/Y sky130_fd_sc_hd__inv_2
XFILLER_92_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16775__A0 _15963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09373_ _20004_/Q vssd1 vssd1 vccd1 vccd1 _09465_/A sky130_fd_sc_hd__inv_2
XFILLER_197_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17221__S _17386_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_4_9_0_HCLK_A clkbuf_4_9_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19559__RESET_B hold348/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_177_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12013__B1 hold305/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_229_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19141__RESET_B repeater274/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09965__C1 _09964_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_4_0_HCLK clkbuf_3_5_0_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_9_0_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_133_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_hold191_A HADDR[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09709_ _09748_/A _19421_/Q _09753_/C _19427_/Q _09708_/Y vssd1 vssd1 vccd1 vccd1
+ _09713_/C sky130_fd_sc_hd__o221a_1
XANTENNA__11827__B1 _10866_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10981_ _10976_/B _10978_/X _10980_/Y _10408_/X _10965_/A vssd1 vssd1 vccd1 vccd1
+ _10982_/A sky130_fd_sc_hd__o32a_1
XFILLER_74_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15018__B1 _15004_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12720_ _14808_/A vssd1 vssd1 vccd1 vccd1 _12720_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__16766__A0 _15963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_230_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12651_ _12651_/A vssd1 vssd1 vccd1 vccd1 _12651_/X sky130_fd_sc_hd__clkbuf_2
XPHY_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19982__RESET_B repeater192/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17131__S _17545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11602_ _11581_/A _11581_/B _11569_/A _11600_/Y vssd1 vssd1 vccd1 vccd1 _19568_/D
+ sky130_fd_sc_hd__a211oi_2
XPHY_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15370_ _19786_/Q _10646_/B _10647_/B vssd1 vssd1 vccd1 vccd1 _15370_/X sky130_fd_sc_hd__a21bo_1
XFILLER_157_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12582_ _19042_/Q _12576_/X _12410_/X _12577_/X vssd1 vssd1 vccd1 vccd1 _19042_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_148_HCLK clkbuf_4_1_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19865_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14321_ _18441_/Q _14318_/X _14273_/X _14320_/X vssd1 vssd1 vccd1 vccd1 _18441_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17191__A0 _15768_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11533_ _19585_/Q _11532_/Y _11521_/X _11533_/C1 vssd1 vssd1 vccd1 vccd1 _19585_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16970__S _17523_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17040_ _17039_/X _11332_/Y _17493_/S vssd1 vssd1 vccd1 vccd1 _17040_/X sky130_fd_sc_hd__mux2_1
XPHY_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11464_ _11464_/A _11535_/A vssd1 vssd1 vccd1 vccd1 _11465_/B sky130_fd_sc_hd__or2_1
XANTENNA__12004__B1 _09016_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14252_ _14252_/A vssd1 vssd1 vccd1 vccd1 _14252_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_183_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10415_ _14680_/A _15826_/A vssd1 vssd1 vccd1 vccd1 _16434_/B sky130_fd_sc_hd__or2_4
X_13203_ _13068_/A _13203_/A2 _13200_/Y _13202_/X vssd1 vssd1 vccd1 vccd1 _18895_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_137_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14183_ _14180_/Y _18697_/Q _16467_/A _18680_/Q _14182_/X vssd1 vssd1 vccd1 vccd1
+ _14184_/D sky130_fd_sc_hd__o221a_1
X_11395_ _11572_/A _19139_/Q _19559_/Q _11391_/Y _11394_/X vssd1 vssd1 vccd1 vccd1
+ _11412_/A sky130_fd_sc_hd__o221a_1
XFILLER_124_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10346_ _10341_/B _10320_/X _10344_/Y _10345_/X _10330_/A vssd1 vssd1 vccd1 vccd1
+ _10347_/A sky130_fd_sc_hd__o32a_1
X_13134_ _13131_/Y _18892_/Q _19161_/Q _13063_/A _13133_/X vssd1 vssd1 vccd1 vccd1
+ _13144_/B sky130_fd_sc_hd__o221a_1
X_18991_ _19115_/CLK _18991_/D hold273/X vssd1 vssd1 vccd1 vccd1 _18991_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_140_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17942_ _19842_/CLK _17942_/D vssd1 vssd1 vccd1 vccd1 _17942_/Q sky130_fd_sc_hd__dfxtp_1
X_13065_ _13065_/A _13207_/A vssd1 vssd1 vccd1 vccd1 _13066_/B sky130_fd_sc_hd__or2_1
XANTENNA__18864__RESET_B repeater231/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10277_ _19642_/Q vssd1 vssd1 vccd1 vccd1 _14334_/A sky130_fd_sc_hd__inv_2
XANTENNA_repeater209_A repeater210/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_238_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12016_ _12016_/A vssd1 vssd1 vccd1 vccd1 _12016_/X sky130_fd_sc_hd__clkbuf_2
Xrepeater208 repeater210/X vssd1 vssd1 vccd1 vccd1 repeater208/X sky130_fd_sc_hd__buf_8
X_17873_ _16164_/Y _16165_/Y _16166_/Y _16167_/Y _17913_/S0 _19632_/Q vssd1 vssd1
+ vccd1 vccd1 _17873_/X sky130_fd_sc_hd__mux4_2
Xrepeater219 repeater226/X vssd1 vssd1 vccd1 vccd1 repeater219/X sky130_fd_sc_hd__clkbuf_8
X_16824_ _16823_/X _09491_/A _17482_/S vssd1 vssd1 vccd1 vccd1 _16824_/X sky130_fd_sc_hd__mux2_1
X_19612_ _20048_/CLK _19612_/D repeater191/X vssd1 vssd1 vccd1 vccd1 _19612_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__17306__S _17544_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_247_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19543_ _19544_/CLK _19543_/D repeater221/X vssd1 vssd1 vccd1 vccd1 _19543_/Q sky130_fd_sc_hd__dfrtp_1
X_16755_ vssd1 vssd1 vccd1 vccd1 _16755_/HI _16755_/LO sky130_fd_sc_hd__conb_1
XANTENNA__11818__B1 _09077_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13967_ _13967_/A vssd1 vssd1 vccd1 vccd1 _13970_/A sky130_fd_sc_hd__inv_2
XFILLER_34_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15706_ _19897_/Q _10133_/B _08982_/A vssd1 vssd1 vccd1 vccd1 _18642_/D sky130_fd_sc_hd__a21o_2
XFILLER_234_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19474_ _19513_/CLK hold208/X repeater259/X vssd1 vssd1 vccd1 vccd1 _19474_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_62_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12918_ _12917_/Y _18937_/Q _19280_/Q _12965_/B vssd1 vssd1 vccd1 vccd1 _12924_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_61_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16686_ _17017_/X _16683_/X _17035_/X _16684_/X _16685_/X vssd1 vssd1 vccd1 vccd1
+ _16691_/B sky130_fd_sc_hd__o221a_4
X_13898_ _13850_/X _13898_/B _13898_/C _13898_/D vssd1 vssd1 vccd1 vccd1 _13899_/A
+ sky130_fd_sc_hd__and4b_1
XFILLER_222_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18425_ _18441_/CLK _18425_/D vssd1 vssd1 vccd1 vccd1 _18425_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_179_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15637_ _18602_/Q _15629_/A _18603_/Q vssd1 vssd1 vccd1 vccd1 _15637_/X sky130_fd_sc_hd__o21a_1
XFILLER_222_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12849_ _18935_/Q vssd1 vssd1 vccd1 vccd1 _12877_/A sky130_fd_sc_hd__inv_2
XFILLER_61_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_210_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17041__S _17548_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18356_ _18416_/CLK _18356_/D vssd1 vssd1 vccd1 vccd1 _18356_/Q sky130_fd_sc_hd__dfxtp_1
X_15568_ _15566_/Y _15567_/X _15542_/X vssd1 vssd1 vccd1 vccd1 _15568_/X sky130_fd_sc_hd__o21a_1
XFILLER_202_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12794__A1 _19250_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17307_ _17306_/X _13845_/Y _17545_/S vssd1 vssd1 vccd1 vccd1 _17307_/X sky130_fd_sc_hd__mux2_1
XFILLER_175_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14519_ _14519_/A vssd1 vssd1 vccd1 vccd1 _14520_/A sky130_fd_sc_hd__inv_2
XANTENNA__17182__A0 _15768_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16880__S _17413_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18287_ _18435_/CLK _18287_/D vssd1 vssd1 vccd1 vccd1 _18287_/Q sky130_fd_sc_hd__dfxtp_1
X_15499_ _18568_/Q _15490_/A _18569_/Q vssd1 vssd1 vccd1 vccd1 _15499_/X sky130_fd_sc_hd__o21a_1
X_17238_ _15768_/Y _11200_/Y _17546_/S vssd1 vssd1 vccd1 vccd1 _17238_/X sky130_fd_sc_hd__mux2_1
XFILLER_162_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11349__A2 _18968_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12546__A1 hold242/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17169_ _17168_/X _15635_/Y _17318_/S vssd1 vssd1 vccd1 vccd1 _17169_/X sky130_fd_sc_hd__mux2_2
XFILLER_143_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17485__A1 _13529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09991_ _09856_/A _09856_/B _09988_/Y _09990_/X vssd1 vssd1 vccd1 vccd1 _19947_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_88_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08942_ _10321_/C _18774_/Q _19854_/Q _08941_/Y vssd1 vssd1 vccd1 vccd1 _08943_/D
+ sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_29_HCLK clkbuf_4_9_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20089_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_85_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17216__S _17543_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_217_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11809__B1 hold276/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10669__A _10676_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_231_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_225_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12482__B1 _12232_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09425_ _19937_/Q vssd1 vssd1 vccd1 vccd1 _09425_/Y sky130_fd_sc_hd__inv_2
XFILLER_212_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_212_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_185_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09356_ _20021_/Q vssd1 vssd1 vccd1 vccd1 _09481_/A sky130_fd_sc_hd__inv_2
XFILLER_139_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_240_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17173__A0 _17486_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09287_ _09294_/A vssd1 vssd1 vccd1 vccd1 _09287_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__16790__S _17548_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16920__A0 _17473_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14526__A2 _14519_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_193_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10200_ _19830_/Q vssd1 vssd1 vccd1 vccd1 _10200_/Y sky130_fd_sc_hd__inv_2
XFILLER_107_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_180_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11180_ _17706_/X _11176_/X _19625_/Q _11178_/X vssd1 vssd1 vccd1 vccd1 _19625_/D
+ sky130_fd_sc_hd__a22o_1
X_10131_ _19905_/Q _10130_/X _10109_/Y vssd1 vssd1 vccd1 vccd1 _19905_/D sky130_fd_sc_hd__o21a_1
XANTENNA__09166__B1 hold344/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10062_ _10062_/A vssd1 vssd1 vccd1 vccd1 _10062_/Y sky130_fd_sc_hd__inv_2
XFILLER_236_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11963__A _11979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17126__S _17318_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18665__SET_B repeater222/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16987__A0 _15768_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14870_ _15121_/A _15109_/B _15145_/C vssd1 vssd1 vccd1 vccd1 _14872_/A sky130_fd_sc_hd__or3_4
XFILLER_236_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18168__CLK _18169_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_229_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16451__A2 _15867_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13821_ _13910_/A _13821_/B vssd1 vssd1 vccd1 vccd1 _13932_/A sky130_fd_sc_hd__or2_1
XFILLER_63_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16965__S _17474_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16540_ _17152_/X _16512_/X _17135_/X _16513_/X _16539_/X vssd1 vssd1 vccd1 vccd1
+ _16540_/X sky130_fd_sc_hd__o221a_4
XFILLER_244_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12473__B1 _12353_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13752_ _13749_/Y _13751_/A _18746_/Q _13750_/A vssd1 vssd1 vccd1 vccd1 _13753_/B
+ sky130_fd_sc_hd__o22a_1
X_10964_ _10964_/A _10983_/A vssd1 vssd1 vccd1 vccd1 _10979_/A sky130_fd_sc_hd__or2_1
XFILLER_232_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12703_ _18963_/Q _12698_/X _12536_/X _12699_/X vssd1 vssd1 vccd1 vccd1 _18963_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_105_HCLK_A clkbuf_4_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16471_ _16471_/A _16544_/B vssd1 vssd1 vccd1 vccd1 _16471_/Y sky130_fd_sc_hd__nor2_1
X_13683_ _18772_/Q _13671_/A _13682_/X _13672_/A vssd1 vssd1 vccd1 vccd1 _18772_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_188_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10895_ _10895_/A vssd1 vssd1 vccd1 vccd1 _10895_/X sky130_fd_sc_hd__clkbuf_2
X_18210_ _18333_/CLK _18210_/D vssd1 vssd1 vccd1 vccd1 _18210_/Q sky130_fd_sc_hd__dfxtp_1
X_15422_ _19613_/Q _11158_/B _11159_/B vssd1 vssd1 vccd1 vccd1 _15422_/X sky130_fd_sc_hd__a21bo_1
XFILLER_31_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12634_ _19010_/Q _12629_/X _12408_/X _12630_/X vssd1 vssd1 vccd1 vccd1 _19010_/D
+ sky130_fd_sc_hd__a22o_1
X_19190_ _19952_/CLK _19190_/D repeater244/X vssd1 vssd1 vccd1 vccd1 _19190_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_231_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18141_ _19510_/CLK _18141_/D vssd1 vssd1 vccd1 vccd1 _18141_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17164__A0 _15963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15353_ _18498_/Q _14228_/B _14229_/B vssd1 vssd1 vccd1 vccd1 _15353_/X sky130_fd_sc_hd__a21bo_1
XPHY_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12565_ _19055_/Q _12560_/X _12380_/X _12563_/X vssd1 vssd1 vccd1 vccd1 _19055_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_repeater159_A _17490_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14304_ _14304_/A vssd1 vssd1 vccd1 vccd1 _14305_/A sky130_fd_sc_hd__inv_2
XPHY_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11516_ _11474_/A _11474_/B _11506_/X _11514_/Y vssd1 vssd1 vccd1 vccd1 _19594_/D
+ sky130_fd_sc_hd__a211oi_2
XPHY_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18072_ _18169_/CLK _18072_/D vssd1 vssd1 vccd1 vccd1 _18072_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15284_ _15254_/Y _15436_/A _18630_/Q vssd1 vssd1 vccd1 vccd1 _15285_/B sky130_fd_sc_hd__a21oi_1
XPHY_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12496_ _19089_/Q _12489_/X _12384_/X _12492_/X vssd1 vssd1 vccd1 vccd1 _19089_/D
+ sky130_fd_sc_hd__a22o_1
X_17023_ _17022_/X _12952_/Y _17541_/S vssd1 vssd1 vccd1 vccd1 _17023_/X sky130_fd_sc_hd__mux2_1
X_14235_ _14235_/A vssd1 vssd1 vccd1 vccd1 _17600_/S sky130_fd_sc_hd__buf_8
X_11447_ _19551_/Q vssd1 vssd1 vccd1 vccd1 _11621_/A sky130_fd_sc_hd__inv_2
XFILLER_124_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output88_A _16607_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14166_ _14166_/A _14166_/B _14166_/C _14166_/D vssd1 vssd1 vccd1 vccd1 _14166_/X
+ sky130_fd_sc_hd__and4_1
X_11378_ _19553_/Q vssd1 vssd1 vccd1 vccd1 _11623_/A sky130_fd_sc_hd__inv_2
X_10329_ _10329_/A _10348_/A vssd1 vssd1 vccd1 vccd1 _10343_/A sky130_fd_sc_hd__or2_1
X_13117_ _13114_/Y _18917_/Q _19188_/Q _13089_/A _13116_/X vssd1 vssd1 vccd1 vccd1
+ _13127_/B sky130_fd_sc_hd__o221a_1
X_14097_ _18703_/Q _14033_/Y _14034_/Y _14033_/A _14096_/X vssd1 vssd1 vccd1 vccd1
+ _18703_/D sky130_fd_sc_hd__o221a_1
X_18974_ _19576_/CLK _18974_/D repeater282/X vssd1 vssd1 vccd1 vccd1 _18974_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_113_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17925_ _19544_/CLK _19672_/Q vssd1 vssd1 vccd1 vccd1 _17925_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13048_ _18898_/Q vssd1 vssd1 vccd1 vccd1 _13070_/A sky130_fd_sc_hd__inv_2
XFILLER_39_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11873__A _15772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17856_ _16279_/Y _16280_/Y _16281_/Y _16282_/Y _17908_/S0 _18759_/Q vssd1 vssd1
+ vccd1 vccd1 _17856_/X sky130_fd_sc_hd__mux4_2
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16807_ _15963_/X _12746_/Y _17534_/S vssd1 vssd1 vccd1 vccd1 _16807_/X sky130_fd_sc_hd__mux2_1
XFILLER_226_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17787_ _18326_/Q _18006_/Q _18310_/Q _18302_/Q _17923_/S0 _19646_/Q vssd1 vssd1
+ vccd1 vccd1 _17787_/X sky130_fd_sc_hd__mux4_2
XANTENNA__16875__S _17542_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14999_ _18055_/Q _14991_/X _14998_/X _14994_/X vssd1 vssd1 vccd1 vccd1 _18055_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19526_ _19771_/CLK _19526_/D repeater189/X vssd1 vssd1 vccd1 vccd1 _19526_/Q sky130_fd_sc_hd__dfstp_1
X_16738_ _19056_/Q vssd1 vssd1 vccd1 vccd1 _16738_/Y sky130_fd_sc_hd__inv_2
XFILLER_47_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_241_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_234_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20070__CLK _20070_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19457_ _19462_/CLK _19457_/D repeater272/X vssd1 vssd1 vccd1 vccd1 _19457_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_34_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16669_ _16669_/A vssd1 vssd1 vccd1 vccd1 _16718_/B sky130_fd_sc_hd__buf_4
XFILLER_61_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09210_ _18648_/Q _09238_/A vssd1 vssd1 vccd1 vccd1 _09211_/A sky130_fd_sc_hd__nand2_1
XANTENNA__12216__B1 _12028_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18408_ _18473_/CLK _18408_/D vssd1 vssd1 vccd1 vccd1 _18408_/Q sky130_fd_sc_hd__dfxtp_1
X_19388_ _19933_/CLK _19388_/D repeater235/X vssd1 vssd1 vccd1 vccd1 _19388_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_194_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_203_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_194_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09141_ _15322_/A _09139_/Y _09140_/Y vssd1 vssd1 vccd1 vccd1 _09141_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA_clkbuf_leaf_27_HCLK_A clkbuf_4_9_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18339_ _18954_/CLK _18339_/D vssd1 vssd1 vccd1 vccd1 _18339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_175_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09072_ _09087_/A vssd1 vssd1 vccd1 vccd1 _09072_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_163_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_190_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18715__RESET_B repeater252/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09974_ _09865_/A _09865_/B _09972_/Y _09970_/X vssd1 vssd1 vccd1 vccd1 _19957_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_104_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08925_ _10329_/A _18783_/Q _19863_/Q _08924_/Y vssd1 vssd1 vccd1 vccd1 _08925_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_76_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20094_ _20107_/CLK _20094_/D repeater234/X vssd1 vssd1 vccd1 vccd1 _20094_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_112_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11783__A _11821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16969__A0 _17473_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_218_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16785__S _17512_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12455__B1 _12396_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold154_A HADDR[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_214_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_198_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_198_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09408_ _10087_/A _19375_/Q _19915_/Q _09407_/Y vssd1 vssd1 vccd1 vccd1 _09416_/A
+ sky130_fd_sc_hd__o22a_1
X_10680_ _17741_/X _10676_/X _19784_/Q _10677_/X vssd1 vssd1 vccd1 vccd1 _19784_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12207__B1 _12095_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_213_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_179_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09339_ _14780_/A vssd1 vssd1 vccd1 vccd1 _09339_/X sky130_fd_sc_hd__buf_2
XFILLER_187_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12350_ hold271/X vssd1 vssd1 vccd1 vccd1 hold270/A sky130_fd_sc_hd__buf_4
XFILLER_166_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_217_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11301_ _18984_/Q vssd1 vssd1 vccd1 vccd1 _11301_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17792__S1 _19646_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12281_ _19211_/Q _12276_/X _12102_/X _12277_/X vssd1 vssd1 vccd1 vccd1 _19211_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_126_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14020_ _14020_/A _14020_/B vssd1 vssd1 vccd1 vccd1 _14120_/A sky130_fd_sc_hd__or2_1
X_11232_ _19591_/Q vssd1 vssd1 vccd1 vccd1 _11471_/A sky130_fd_sc_hd__inv_2
XFILLER_153_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11163_ _19618_/Q _11163_/B vssd1 vssd1 vccd1 vccd1 _11164_/B sky130_fd_sc_hd__or2_1
XFILLER_1_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10114_ _18561_/Q _15462_/A vssd1 vssd1 vccd1 vccd1 _15466_/A sky130_fd_sc_hd__or2_1
XFILLER_49_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15971_ _15971_/A vssd1 vssd1 vccd1 vccd1 _15971_/X sky130_fd_sc_hd__clkbuf_2
X_11094_ _17755_/X vssd1 vssd1 vccd1 vccd1 _11094_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17710_ _15430_/X _19767_/Q _18546_/D vssd1 vssd1 vccd1 vccd1 _17710_/X sky130_fd_sc_hd__mux2_1
X_10045_ _10045_/A _10062_/A vssd1 vssd1 vccd1 vccd1 _10046_/B sky130_fd_sc_hd__or2_2
XFILLER_96_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14922_ _14922_/A vssd1 vssd1 vccd1 vccd1 _14923_/A sky130_fd_sc_hd__inv_2
X_18690_ _18701_/CLK _18690_/D hold359/X vssd1 vssd1 vccd1 vccd1 _18690_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_248_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12694__B1 hold250/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17641_ _15674_/X _19048_/Q _17655_/S vssd1 vssd1 vccd1 vccd1 _18611_/D sky130_fd_sc_hd__mux2_1
XANTENNA__09163__A _09164_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14853_ _18140_/Q _14846_/A _14814_/X _14847_/A vssd1 vssd1 vccd1 vccd1 _18140_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_output126_A _15778_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13804_ _18710_/Q vssd1 vssd1 vccd1 vccd1 _13947_/A sky130_fd_sc_hd__inv_2
XFILLER_91_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17572_ _15416_/X _19771_/Q _17584_/S vssd1 vssd1 vccd1 vccd1 _17572_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12446__B1 _12380_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14784_ _14819_/A _14975_/B _14784_/C vssd1 vssd1 vccd1 vccd1 _14786_/A sky130_fd_sc_hd__or3_4
XFILLER_223_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11996_ _11996_/A _16053_/A vssd1 vssd1 vccd1 vccd1 _12187_/B sky130_fd_sc_hd__or2_4
XFILLER_216_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19311_ _19315_/CLK _19311_/D repeater214/X vssd1 vssd1 vccd1 vccd1 _19311_/Q sky130_fd_sc_hd__dfrtp_2
X_16523_ _17290_/X _16512_/X _17272_/X _16513_/X _16522_/X vssd1 vssd1 vccd1 vccd1
+ _16523_/X sky130_fd_sc_hd__o221a_4
X_13735_ _13733_/A _14286_/B _13733_/Y vssd1 vssd1 vccd1 vccd1 _18753_/D sky130_fd_sc_hd__a21oi_1
XFILLER_188_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10947_ _10949_/A vssd1 vssd1 vccd1 vccd1 _11771_/A sky130_fd_sc_hd__buf_2
XANTENNA__14509__A hold325/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_188_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19242_ _19314_/CLK _19242_/D repeater239/X vssd1 vssd1 vccd1 vccd1 _19242_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_204_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16454_ _19822_/Q vssd1 vssd1 vccd1 vccd1 _16454_/Y sky130_fd_sc_hd__inv_2
XFILLER_149_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13666_ _18782_/Q _13664_/X hold250/X _13665_/X vssd1 vssd1 vccd1 vccd1 _18782_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_32_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10878_ _10878_/A vssd1 vssd1 vccd1 vccd1 _10879_/A sky130_fd_sc_hd__inv_2
X_15405_ _15413_/A _17578_/X vssd1 vssd1 vccd1 vccd1 _18534_/D sky130_fd_sc_hd__and2_1
XPHY_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12617_ _19023_/Q _12613_/X _12375_/X _12616_/X vssd1 vssd1 vccd1 vccd1 _19023_/D
+ sky130_fd_sc_hd__a22o_1
X_19173_ _19208_/CLK _19173_/D hold370/X vssd1 vssd1 vccd1 vccd1 _19173_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16385_ _19821_/Q vssd1 vssd1 vccd1 vccd1 _16385_/Y sky130_fd_sc_hd__inv_2
XPHY_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13597_ _13597_/A _13597_/B _13597_/C vssd1 vssd1 vccd1 vccd1 _18814_/D sky130_fd_sc_hd__nor3_1
XFILLER_157_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18124_ _18765_/CLK _18124_/D vssd1 vssd1 vccd1 vccd1 _18124_/Q sky130_fd_sc_hd__dfxtp_1
X_15336_ _15336_/A _17600_/X vssd1 vssd1 vccd1 vccd1 _18490_/D sky130_fd_sc_hd__nor2_1
X_12548_ _12246_/B _12249_/A _12551_/C vssd1 vssd1 vccd1 vccd1 _12548_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_247_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15699__B1 _15673_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17783__S1 _19646_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18055_ _18142_/CLK _18055_/D vssd1 vssd1 vccd1 vccd1 _18055_/Q sky130_fd_sc_hd__dfxtp_1
X_15267_ _15443_/A _15437_/B _15242_/Y _15266_/X vssd1 vssd1 vccd1 vccd1 _18633_/D
+ sky130_fd_sc_hd__o31ai_1
XANTENNA__15163__A2 _15158_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12479_ _12479_/A vssd1 vssd1 vccd1 vccd1 _12479_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_144_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17006_ _17005_/X _15526_/A _17513_/S vssd1 vssd1 vccd1 vccd1 _17006_/X sky130_fd_sc_hd__mux2_1
X_14218_ _14218_/A _14218_/B _14218_/C _14218_/D vssd1 vssd1 vccd1 vccd1 _14219_/D
+ sky130_fd_sc_hd__and4_1
X_15198_ _16434_/B vssd1 vssd1 vccd1 vccd1 _17565_/S sky130_fd_sc_hd__inv_4
XFILLER_153_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12921__A1 _12919_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14149_ _18673_/Q _14148_/Y _14149_/B1 _14112_/X vssd1 vssd1 vccd1 vccd1 _18673_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_86_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18957_ _18959_/CLK _18957_/D repeater257/X vssd1 vssd1 vccd1 vccd1 _18957_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12699__A _12699_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17908_ _15814_/Y _15815_/Y _15816_/Y _15817_/Y _17908_/S0 _18759_/Q vssd1 vssd1
+ vccd1 vccd1 _17908_/X sky130_fd_sc_hd__mux4_1
X_09690_ _19419_/Q vssd1 vssd1 vccd1 vccd1 _09690_/Y sky130_fd_sc_hd__inv_2
X_18888_ _19222_/CLK _18888_/D repeater188/X vssd1 vssd1 vccd1 vccd1 _18888_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_67_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrebuffer14 _14014_/B vssd1 vssd1 vccd1 vccd1 _14133_/C1 sky130_fd_sc_hd__dlygate4sd1_1
X_17839_ _17835_/X _17836_/X _17837_/X _17838_/X _18760_/Q _18761_/Q vssd1 vssd1 vccd1
+ vccd1 _17839_/X sky130_fd_sc_hd__mux4_2
XFILLER_94_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrebuffer25 _14007_/B vssd1 vssd1 vccd1 vccd1 _14144_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_55_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xrebuffer36 _19418_/Q vssd1 vssd1 vccd1 vccd1 _11897_/A1 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_212_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrebuffer47 _13551_/B vssd1 vssd1 vccd1 vccd1 _13575_/C1 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer58 _09388_/B2 vssd1 vssd1 vccd1 vccd1 _11954_/A1 sky130_fd_sc_hd__dlygate4sd1_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xrebuffer69 _14016_/B vssd1 vssd1 vccd1 vccd1 _14128_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XANTENNA__16618__B _16621_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19509_ _19510_/CLK hold223/X repeater256/X vssd1 vssd1 vccd1 vccd1 _19509_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__10947__A _10949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_151_HCLK_A clkbuf_4_1_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_176_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16634__A _16634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrebuffer104 _10025_/A vssd1 vssd1 vccd1 vccd1 _10057_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_41_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09124_ _20085_/Q vssd1 vssd1 vccd1 vccd1 _09125_/D sky130_fd_sc_hd__inv_2
XFILLER_148_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrebuffer115 _14022_/B vssd1 vssd1 vccd1 vccd1 _14119_/A2 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer126 _13549_/B vssd1 vssd1 vccd1 vccd1 _13578_/C1 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_157_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09055_ _09087_/A vssd1 vssd1 vccd1 vccd1 _09055_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_163_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17774__S1 _19648_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11778__A _12659_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14362__B1 _14326_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_237_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13993__A _18681_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09957_ _09957_/A vssd1 vssd1 vccd1 vccd1 _09957_/Y sky130_fd_sc_hd__inv_2
XFILLER_104_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12676__B1 hold298/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20077_ _20077_/CLK _20077_/D repeater196/X vssd1 vssd1 vccd1 vccd1 _20077_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12402__A _12402_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09888_ _19360_/Q vssd1 vssd1 vccd1 vccd1 _16721_/A sky130_fd_sc_hd__inv_2
XANTENNA_hold369_A scl_i_S4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_245_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_218_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17404__S _17568_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11850_ _19433_/Q vssd1 vssd1 vccd1 vccd1 _11867_/A sky130_fd_sc_hd__inv_2
XFILLER_17_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_233_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10801_ _10801_/A _10801_/B vssd1 vssd1 vccd1 vccd1 _10801_/Y sky130_fd_sc_hd__nor2_2
XPHY_4567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11781_ _12371_/A _16238_/A vssd1 vssd1 vccd1 vccd1 _11933_/A sky130_fd_sc_hd__or2_4
XPHY_4589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13520_ _14695_/A vssd1 vssd1 vccd1 vccd1 _14668_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_241_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10732_ _19542_/Q _10732_/B _10732_/C vssd1 vssd1 vccd1 vccd1 _10733_/A sky130_fd_sc_hd__or3_1
XFILLER_41_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15917__A1 _17513_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_3888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15917__B2 _16505_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13451_ _18856_/Q _13450_/Y _13426_/X _13344_/B vssd1 vssd1 vccd1 vccd1 _18856_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__17119__A0 _17473_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10663_ _10677_/A vssd1 vssd1 vccd1 vccd1 _10663_/X sky130_fd_sc_hd__clkbuf_2
X_12402_ _12402_/A vssd1 vssd1 vccd1 vccd1 _12402_/X sky130_fd_sc_hd__buf_1
XANTENNA_clkbuf_leaf_10_HCLK_A clkbuf_4_2_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16170_ _16024_/Y _16169_/Y _19651_/Q vssd1 vssd1 vccd1 vccd1 _16170_/X sky130_fd_sc_hd__o21a_1
X_10594_ _10594_/A _10594_/B _10594_/C vssd1 vssd1 vccd1 vccd1 _10616_/B sky130_fd_sc_hd__or3_1
X_13382_ _20110_/Q _13429_/C _13380_/Y _18856_/Q _13381_/X vssd1 vssd1 vccd1 vccd1
+ _13386_/C sky130_fd_sc_hd__o221a_1
XANTENNA_clkbuf_leaf_73_HCLK_A clkbuf_opt_4_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17765__S1 _19646_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15121_ _15121_/A _18764_/Q _15121_/C vssd1 vssd1 vccd1 vccd1 _15123_/A sky130_fd_sc_hd__or3_4
X_12333_ _19180_/Q _12327_/X _12092_/X _12328_/X vssd1 vssd1 vccd1 vccd1 _19180_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_182_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15052_ _18023_/Q _15047_/X _14998_/X _15049_/X vssd1 vssd1 vccd1 vccd1 _18023_/D
+ sky130_fd_sc_hd__a22o_1
X_12264_ _19224_/Q _12260_/X _12069_/X _12263_/X vssd1 vssd1 vccd1 vccd1 _19224_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_147_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14003_ _14003_/A _14003_/B vssd1 vssd1 vccd1 vccd1 _14148_/A sky130_fd_sc_hd__or2_1
X_11215_ _11477_/A _19011_/Q _19597_/Q _11214_/Y vssd1 vssd1 vccd1 vccd1 _11215_/X
+ sky130_fd_sc_hd__o22a_1
X_12195_ _19256_/Q _12189_/X _12076_/X _12192_/X vssd1 vssd1 vccd1 vccd1 _19256_/D
+ sky130_fd_sc_hd__a22o_1
X_19860_ _19867_/CLK _19860_/D repeater263/X vssd1 vssd1 vccd1 vccd1 _19860_/Q sky130_fd_sc_hd__dfrtp_1
X_18811_ _20115_/CLK _18811_/D repeater238/X vssd1 vssd1 vccd1 vccd1 _18811_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__19751__CLK _20070_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput83 _16541_/Y vssd1 vssd1 vccd1 vccd1 HRDATA[13] sky130_fd_sc_hd__clkbuf_2
X_11146_ _11144_/A _11139_/A _11144_/Y vssd1 vssd1 vccd1 vccd1 _19628_/D sky130_fd_sc_hd__a21oi_1
X_19791_ _19794_/CLK _19791_/D repeater203/X vssd1 vssd1 vccd1 vccd1 _19791_/Q sky130_fd_sc_hd__dfrtp_1
Xoutput94 _16664_/Y vssd1 vssd1 vccd1 vccd1 HRDATA[23] sky130_fd_sc_hd__clkbuf_2
XFILLER_95_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11077_ _19519_/Q vssd1 vssd1 vccd1 vccd1 _15858_/A sky130_fd_sc_hd__clkbuf_4
X_15954_ _18099_/Q vssd1 vssd1 vccd1 vccd1 _15954_/Y sky130_fd_sc_hd__inv_2
X_18742_ _20066_/CLK _18742_/D repeater209/X vssd1 vssd1 vccd1 vccd1 _18742_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12667__B1 hold289/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_236_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10028_ _10029_/B vssd1 vssd1 vccd1 vccd1 _10032_/A sky130_fd_sc_hd__buf_2
X_14905_ _18107_/Q _14897_/A _14713_/X _14898_/A vssd1 vssd1 vccd1 vccd1 _18107_/D
+ sky130_fd_sc_hd__a22o_1
X_18673_ _18718_/CLK _18673_/D repeater252/X vssd1 vssd1 vccd1 vccd1 _18673_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__19425__RESET_B repeater274/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15885_ _17549_/X vssd1 vssd1 vccd1 vccd1 _15885_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_236_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17314__S _17568_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17624_ _19895_/Q _19748_/Q _17630_/S vssd1 vssd1 vccd1 vccd1 _17624_/X sky130_fd_sc_hd__mux2_1
X_14836_ _18152_/Q _14832_/X _14806_/X _14834_/X vssd1 vssd1 vccd1 vccd1 _18152_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12419__B1 hold270/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11890__A1 _19423_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17555_ _20059_/Q _19868_/Q _19499_/Q vssd1 vssd1 vccd1 vccd1 _17555_/X sky130_fd_sc_hd__mux2_1
X_14767_ _18188_/Q _14760_/A _14727_/X _14761_/A vssd1 vssd1 vccd1 vccd1 _18188_/D
+ sky130_fd_sc_hd__a22o_1
X_11979_ _11979_/A vssd1 vssd1 vccd1 vccd1 _11979_/X sky130_fd_sc_hd__clkbuf_2
X_16506_ _16506_/A vssd1 vssd1 vccd1 vccd1 _16506_/X sky130_fd_sc_hd__buf_1
XFILLER_177_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13718_ _14629_/B _13717_/Y _14629_/B _13717_/Y vssd1 vssd1 vccd1 vccd1 _13721_/C
+ sky130_fd_sc_hd__a2bb2o_1
X_17486_ _17486_/A0 _13156_/Y _17543_/S vssd1 vssd1 vccd1 vccd1 _17486_/X sky130_fd_sc_hd__mux2_1
X_14698_ _14700_/A vssd1 vssd1 vccd1 vccd1 _14698_/X sky130_fd_sc_hd__clkbuf_2
X_19225_ _19849_/CLK _19225_/D repeater257/X vssd1 vssd1 vccd1 vccd1 _19225_/Q sky130_fd_sc_hd__dfrtp_4
X_16437_ _16437_/A _18744_/Q vssd1 vssd1 vccd1 vccd1 _16437_/Y sky130_fd_sc_hd__nand2_1
X_13649_ _16955_/X _13644_/X _18792_/Q _13646_/X vssd1 vssd1 vccd1 vccd1 _18792_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13395__A1 _20095_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19156_ _19576_/CLK _19156_/D repeater268/X vssd1 vssd1 vccd1 vccd1 _19156_/Q sky130_fd_sc_hd__dfrtp_1
X_16368_ _19132_/Q vssd1 vssd1 vccd1 vccd1 _16368_/Y sky130_fd_sc_hd__inv_2
XFILLER_191_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_200_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18107_ _18260_/CLK _18107_/D vssd1 vssd1 vccd1 vccd1 _18107_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_191_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15319_ _15319_/A _15319_/B vssd1 vssd1 vccd1 vccd1 _15319_/X sky130_fd_sc_hd__or2_1
XFILLER_184_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19087_ _19119_/CLK _19087_/D hold351/X vssd1 vssd1 vccd1 vccd1 _19087_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_173_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16299_ _19444_/Q vssd1 vssd1 vccd1 vccd1 _16299_/Y sky130_fd_sc_hd__inv_2
XFILLER_145_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18849__CLK _18866_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14344__B1 _14329_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18038_ _18169_/CLK _18038_/D vssd1 vssd1 vccd1 vccd1 _18038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_20000_ _20003_/CLK _20000_/D repeater192/X vssd1 vssd1 vccd1 vccd1 _20000_/Q sky130_fd_sc_hd__dfrtp_1
X_09811_ _09635_/B _09810_/A _19974_/Q _09813_/A _09759_/X vssd1 vssd1 vccd1 vccd1
+ _19974_/D sky130_fd_sc_hd__o221a_1
XFILLER_86_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_247_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19989_ _19992_/CLK _19989_/D repeater192/X vssd1 vssd1 vccd1 vccd1 _19989_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_98_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09742_ _09742_/A _09742_/B vssd1 vssd1 vccd1 vccd1 _09781_/A sky130_fd_sc_hd__or2_1
XANTENNA__12658__B1 _12543_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09673_ _19426_/Q vssd1 vssd1 vccd1 vccd1 _09673_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17224__S _17544_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_243_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_215_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17349__A0 _17486_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19624__CLK _19920_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14583__B1 _14582_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_176_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_248_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09107_ hold322/X vssd1 vssd1 vccd1 vccd1 _11926_/A sky130_fd_sc_hd__buf_1
XFILLER_184_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09038_ _20114_/Q _09029_/X _09037_/X _09031_/X vssd1 vssd1 vccd1 vccd1 _20114_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_163_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold360 hold360/A vssd1 vssd1 vccd1 vccd1 hold360/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold371 hold371/A vssd1 vssd1 vccd1 vccd1 hold371/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11000_ _10996_/B _10955_/Y _10999_/X _10954_/A _19660_/Q vssd1 vssd1 vccd1 vccd1
+ _19660_/D sky130_fd_sc_hd__a32o_1
XFILLER_219_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12649__B1 _12596_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12132__A _15772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12951_ _19275_/Q vssd1 vssd1 vccd1 vccd1 _12951_/Y sky130_fd_sc_hd__inv_2
XFILLER_19_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11902_ _19415_/Q _11898_/X _09061_/X _11899_/X vssd1 vssd1 vccd1 vccd1 _19415_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17134__S _17413_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15670_ _18609_/Q _15661_/A _15661_/B _18610_/Q vssd1 vssd1 vccd1 vccd1 _15670_/X
+ sky130_fd_sc_hd__o31a_1
XPHY_4320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12882_ _12964_/A _12983_/A vssd1 vssd1 vccd1 vccd1 _12883_/B sky130_fd_sc_hd__or2_2
XFILLER_245_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14621_ _18271_/Q _14616_/X _09174_/X _14618_/X vssd1 vssd1 vccd1 vccd1 _18271_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11833_ _12558_/B _12309_/A vssd1 vssd1 vccd1 vccd1 _11834_/S sky130_fd_sc_hd__or2_1
XPHY_4364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16973__S _17535_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17340_ _16366_/Y _15301_/Y _19498_/Q vssd1 vssd1 vccd1 vccd1 _17340_/X sky130_fd_sc_hd__mux2_1
XPHY_4397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14552_ _18310_/Q _14546_/X _14509_/X _14548_/X vssd1 vssd1 vccd1 vccd1 _18310_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_202_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11764_ _11771_/A vssd1 vssd1 vccd1 vccd1 _11764_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__18818__RESET_B repeater231/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13503_ _18762_/Q vssd1 vssd1 vccd1 vccd1 _13511_/A sky130_fd_sc_hd__inv_2
XFILLER_198_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17271_ _17270_/X _09676_/Y _17523_/S vssd1 vssd1 vccd1 vccd1 _17271_/X sky130_fd_sc_hd__mux2_1
X_10715_ _14793_/A vssd1 vssd1 vccd1 vccd1 _10715_/X sky130_fd_sc_hd__clkbuf_4
XPHY_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14483_ _18351_/Q _14478_/X _12720_/X _14480_/X vssd1 vssd1 vccd1 vccd1 _18351_/D
+ sky130_fd_sc_hd__a22o_1
X_11695_ _19526_/Q _11690_/X _10885_/X _11692_/X vssd1 vssd1 vccd1 vccd1 _19526_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19010_ _19597_/CLK _19010_/D repeater281/X vssd1 vssd1 vccd1 vccd1 _19010_/Q sky130_fd_sc_hd__dfrtp_4
X_16222_ _19677_/Q vssd1 vssd1 vccd1 vccd1 _16222_/Y sky130_fd_sc_hd__inv_2
XPHY_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13434_ _13361_/Y _13350_/A _13433_/X _13387_/Y vssd1 vssd1 vccd1 vccd1 _13435_/C
+ sky130_fd_sc_hd__o31a_1
XFILLER_173_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10646_ _19786_/Q _10646_/B vssd1 vssd1 vccd1 vccd1 _10647_/B sky130_fd_sc_hd__or2_1
XFILLER_201_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11927__A2 _11891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16153_ _18022_/Q vssd1 vssd1 vccd1 vccd1 _16153_/Y sky130_fd_sc_hd__inv_2
Xrebuffer5 _13062_/B vssd1 vssd1 vccd1 vccd1 _13214_/B1 sky130_fd_sc_hd__dlygate4sd1_1
X_13365_ _20091_/Q vssd1 vssd1 vccd1 vccd1 _13365_/Y sky130_fd_sc_hd__inv_2
XFILLER_166_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17512__A0 _17511_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10577_ _19813_/Q _10577_/B _10585_/C vssd1 vssd1 vccd1 vccd1 _10592_/B sky130_fd_sc_hd__or3_4
XFILLER_6_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15104_ _17987_/Q _15096_/A _14816_/A _15097_/A vssd1 vssd1 vccd1 vccd1 _17987_/D
+ sky130_fd_sc_hd__a22o_1
X_12316_ _15769_/A _12316_/B vssd1 vssd1 vccd1 vccd1 _12361_/A sky130_fd_sc_hd__or2_2
X_16084_ _18037_/Q vssd1 vssd1 vccd1 vccd1 _16084_/Y sky130_fd_sc_hd__inv_2
X_13296_ _18756_/Q vssd1 vssd1 vccd1 vccd1 _14819_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_182_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16721__B _16721_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19912_ _20006_/CLK _19912_/D repeater191/X vssd1 vssd1 vccd1 vccd1 _19912_/Q sky130_fd_sc_hd__dfrtp_1
X_15035_ _15036_/A vssd1 vssd1 vccd1 vccd1 _15035_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__17309__S _19498_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12247_ _12247_/A _12247_/B vssd1 vssd1 vccd1 vccd1 _15223_/A sky130_fd_sc_hd__nand2_1
XFILLER_123_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19606__RESET_B hold359/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19843_ _19846_/CLK _19843_/D repeater270/X vssd1 vssd1 vccd1 vccd1 _19843_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_68_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12178_ _19263_/Q _12150_/A _11924_/X _12151_/A vssd1 vssd1 vccd1 vccd1 _19263_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_123_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_229_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17910__S1 _19632_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11129_ _17747_/X _11066_/B _11128_/X vssd1 vssd1 vccd1 vccd1 _19632_/D sky130_fd_sc_hd__a21oi_1
X_19774_ _20049_/CLK _19774_/D repeater190/X vssd1 vssd1 vccd1 vccd1 _19774_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_209_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16986_ _17834_/X _19904_/Q _16986_/S vssd1 vssd1 vccd1 vccd1 _16986_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13381__A1_N _20099_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_62_HCLK clkbuf_opt_3_HCLK/A vssd1 vssd1 vccd1 vccd1 _19933_/CLK sky130_fd_sc_hd__clkbuf_16
X_18725_ _18727_/CLK _18725_/D repeater253/X vssd1 vssd1 vccd1 vccd1 _18725_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_237_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15937_ _16115_/A vssd1 vssd1 vccd1 vccd1 _16483_/B sky130_fd_sc_hd__inv_2
XFILLER_209_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17044__S _17547_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_237_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18656_ _19905_/CLK _18656_/D repeater210/X vssd1 vssd1 vccd1 vccd1 _18656_/Q sky130_fd_sc_hd__dfrtp_1
X_15868_ _15881_/B vssd1 vssd1 vccd1 vccd1 _15878_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_225_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_224_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17607_ _10940_/X _10583_/B _19813_/Q vssd1 vssd1 vccd1 vccd1 _17607_/X sky130_fd_sc_hd__mux2_1
X_14819_ _14819_/A _14975_/B _14975_/C vssd1 vssd1 vccd1 vccd1 _14821_/A sky130_fd_sc_hd__or3_4
XFILLER_24_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15799_ _18226_/Q vssd1 vssd1 vccd1 vccd1 _15799_/Y sky130_fd_sc_hd__inv_2
X_18587_ _19997_/CLK _18587_/D repeater271/X vssd1 vssd1 vccd1 vccd1 _18587_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__16883__S _17523_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_240_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_233_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17538_ _17537_/X _13776_/Y _17548_/S vssd1 vssd1 vccd1 vccd1 _17538_/X sky130_fd_sc_hd__mux2_1
XANTENNA__18559__RESET_B repeater193/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_220_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17469_ _17468_/X _16023_/Y _17565_/S vssd1 vssd1 vccd1 vccd1 _17469_/X sky130_fd_sc_hd__mux2_1
XANTENNA__16554__B2 _15908_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14565__B1 hold330/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19208_ _19208_/CLK _19208_/D hold367/X vssd1 vssd1 vccd1 vccd1 _19208_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_193_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19139_ _19561_/CLK _19139_/D repeater274/X vssd1 vssd1 vccd1 vccd1 _19139_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_218_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17219__S _17534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19347__RESET_B repeater245/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20004__CLK _20091_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17901__S1 _19632_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09725_ _19995_/Q _09724_/Y _09751_/A _19424_/Q vssd1 vssd1 vccd1 vccd1 _09725_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_227_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09656_ _19989_/Q vssd1 vssd1 vccd1 vccd1 _09745_/A sky130_fd_sc_hd__inv_2
XFILLER_227_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16242__B1 _17404_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09261__A _12257_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09587_ _09607_/A vssd1 vssd1 vccd1 vccd1 _09587_/X sky130_fd_sc_hd__buf_2
XFILLER_43_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16793__S _17545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_179_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18911__RESET_B repeater188/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10500_ _19536_/Q _19535_/Q _10514_/C vssd1 vssd1 vccd1 vccd1 _10508_/C sky130_fd_sc_hd__or3_4
XFILLER_195_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14556__B1 _14474_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11480_ _11480_/A _11480_/B vssd1 vssd1 vccd1 vccd1 _11503_/A sky130_fd_sc_hd__or2_1
XPHY_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10854__B _14245_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10431_ _14680_/A _16053_/A vssd1 vssd1 vccd1 vccd1 _15199_/A sky130_fd_sc_hd__or2_4
XFILLER_195_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14308__B1 _14279_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13150_ _19159_/Q _13061_/A _19185_/Q _13086_/A vssd1 vssd1 vccd1 vccd1 _13150_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_152_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10362_ _10358_/B _10368_/A _10361_/X _10354_/X _10361_/A vssd1 vssd1 vccd1 vccd1
+ _10363_/A sky130_fd_sc_hd__o32a_1
XFILLER_124_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12101_ _19313_/Q _12094_/X _12100_/X _12096_/X vssd1 vssd1 vccd1 vccd1 _19313_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11790__B1 hold288/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17129__S _17414_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13081_ _13081_/A _13081_/B vssd1 vssd1 vccd1 vccd1 _13175_/A sky130_fd_sc_hd__or2_1
X_10293_ _19436_/Q vssd1 vssd1 vccd1 vccd1 _10293_/Y sky130_fd_sc_hd__inv_2
XFILLER_88_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12032_ _12032_/A vssd1 vssd1 vccd1 vccd1 _12032_/X sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_85_HCLK clkbuf_4_13_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19314_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold190 input29/X vssd1 vssd1 vccd1 vccd1 hold190/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16968__S _17488_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_238_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16840_ _17473_/A0 _16699_/Y _17042_/S vssd1 vssd1 vccd1 vccd1 _16840_/X sky130_fd_sc_hd__mux2_1
X_16771_ _16770_/X _11425_/Y _17548_/S vssd1 vssd1 vccd1 vccd1 _16771_/X sky130_fd_sc_hd__mux2_1
X_13983_ _18691_/Q vssd1 vssd1 vccd1 vccd1 _14021_/A sky130_fd_sc_hd__inv_2
XFILLER_219_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_219_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18510_ _19780_/CLK _18510_/D repeater226/X vssd1 vssd1 vccd1 vccd1 _18510_/Q sky130_fd_sc_hd__dfrtp_2
X_15722_ _15722_/A _15725_/B vssd1 vssd1 vccd1 vccd1 _18655_/D sky130_fd_sc_hd__nor2_1
X_12934_ _19266_/Q _13002_/A _19290_/Q _12888_/A vssd1 vssd1 vccd1 vccd1 _12934_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_207_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19490_ _19513_/CLK hold173/X repeater260/X vssd1 vssd1 vccd1 vccd1 _19490_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_34_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18441_ _18441_/CLK _18441_/D vssd1 vssd1 vccd1 vccd1 _18441_/Q sky130_fd_sc_hd__dfxtp_1
X_15653_ _18607_/Q vssd1 vssd1 vccd1 vccd1 _15657_/A sky130_fd_sc_hd__inv_2
X_12865_ _13005_/A _13004_/A _13003_/A _13021_/B vssd1 vssd1 vccd1 vccd1 _12871_/C
+ sky130_fd_sc_hd__or4_4
XPHY_4150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_222_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14604_ _14749_/A vssd1 vssd1 vccd1 vccd1 _14604_/X sky130_fd_sc_hd__buf_2
XPHY_4183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18372_ _18795_/CLK _18372_/D vssd1 vssd1 vccd1 vccd1 _18372_/Q sky130_fd_sc_hd__dfxtp_1
X_11816_ _19450_/Q _11814_/X _09071_/X _11815_/X vssd1 vssd1 vccd1 vccd1 _19450_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15584_ _15584_/A vssd1 vssd1 vccd1 vccd1 _15584_/Y sky130_fd_sc_hd__inv_2
XPHY_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12796_ _18830_/Q vssd1 vssd1 vccd1 vccd1 _13553_/A sky130_fd_sc_hd__inv_2
XANTENNA__18652__RESET_B repeater205/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16716__B _16718_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17323_ _17322_/X _09854_/A _17518_/S vssd1 vssd1 vccd1 vccd1 _17323_/X sky130_fd_sc_hd__mux2_1
XFILLER_202_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14535_ _14749_/A vssd1 vssd1 vccd1 vccd1 _14535_/X sky130_fd_sc_hd__clkbuf_2
XPHY_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11747_ hold136/X _10948_/X _19493_/Q _10951_/X vssd1 vssd1 vccd1 vccd1 hold138/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_202_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17254_ _17253_/X _15511_/A _17513_/S vssd1 vssd1 vccd1 vccd1 _17254_/X sky130_fd_sc_hd__mux2_1
XPHY_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14466_ _18361_/Q _14463_/X _14437_/X _14465_/X vssd1 vssd1 vccd1 vccd1 _18361_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11678_ _19539_/Q _11668_/X _10736_/A _11669_/X vssd1 vssd1 vccd1 vccd1 _19539_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_175_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16205_ _20063_/Q _16437_/A vssd1 vssd1 vccd1 vccd1 _16205_/Y sky130_fd_sc_hd__nand2_1
X_13417_ _13405_/X _13417_/B _13417_/C _13417_/D vssd1 vssd1 vccd1 vccd1 _13418_/D
+ sky130_fd_sc_hd__and4b_1
X_10629_ _19804_/Q _10609_/A _10594_/B _10606_/X vssd1 vssd1 vccd1 vccd1 _19804_/D
+ sky130_fd_sc_hd__o22a_1
XANTENNA__19858__RESET_B repeater261/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17185_ _15768_/Y _14212_/Y _17546_/S vssd1 vssd1 vccd1 vccd1 _17185_/X sky130_fd_sc_hd__mux2_1
XFILLER_139_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14397_ _18401_/Q _14394_/X _14351_/X _14396_/X vssd1 vssd1 vccd1 vccd1 _18401_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_139_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16136_ _18875_/Q vssd1 vssd1 vccd1 vccd1 _16136_/Y sky130_fd_sc_hd__inv_2
X_13348_ _13433_/B _13348_/B vssd1 vssd1 vccd1 vccd1 _13439_/A sky130_fd_sc_hd__or2_1
XFILLER_143_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20027__CLK _20115_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17039__S _17546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16067_ _17461_/X vssd1 vssd1 vccd1 vccd1 _16067_/Y sky130_fd_sc_hd__inv_2
X_13279_ _19518_/Q _19517_/Q _13279_/C vssd1 vssd1 vccd1 vccd1 _15909_/A sky130_fd_sc_hd__or3_4
XANTENNA__18074__CLK _18198_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15018_ _18044_/Q _15011_/A _15004_/X _15012_/A vssd1 vssd1 vccd1 vccd1 _18044_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19440__RESET_B repeater193/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16878__S _17482_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19826_ _19841_/CLK _19826_/D repeater271/X vssd1 vssd1 vccd1 vccd1 _19826_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__17895__S0 _17908_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_238_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19757_ _19772_/CLK _19757_/D repeater189/X vssd1 vssd1 vccd1 vccd1 _19757_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_83_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16969_ _17473_/A0 _09921_/Y _17522_/S vssd1 vssd1 vccd1 vccd1 _16969_/X sky130_fd_sc_hd__mux2_1
XFILLER_209_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09510_ _09493_/A _19323_/Q _20011_/Q _09509_/Y vssd1 vssd1 vccd1 vccd1 _09510_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_37_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18708_ _19224_/CLK _18708_/D repeater186/X vssd1 vssd1 vccd1 vccd1 _18708_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_204_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19688_ _19720_/CLK _19688_/D repeater201/X vssd1 vssd1 vccd1 vccd1 _19688_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_64_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09081__A hold248/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09441_ _19918_/Q vssd1 vssd1 vccd1 vccd1 _10034_/A sky130_fd_sc_hd__inv_2
X_18639_ _19810_/CLK _18639_/D repeater224/X vssd1 vssd1 vccd1 vccd1 _18639_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_92_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_197_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17502__S _17567_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_240_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09372_ _20005_/Q vssd1 vssd1 vccd1 vccd1 _09466_/A sky130_fd_sc_hd__inv_2
XFILLER_240_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_178_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_177_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_193_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_opt_1_HCLK_A clkbuf_opt_1_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_229_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09256__A _11936_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16788__S _17474_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_181_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17886__S0 _17908_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold184_A HADDR[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20086__RESET_B repeater205/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16463__B1 _16768_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13277__B1 _18750_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09708_ _09748_/A _19421_/Q _09750_/A _19423_/Q vssd1 vssd1 vccd1 vccd1 _09708_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_114_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_244_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12410__A hold294/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10980_ _19665_/Q _10980_/B vssd1 vssd1 vccd1 vccd1 _10980_/Y sky130_fd_sc_hd__nor2_1
XFILLER_243_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09639_ _19972_/Q vssd1 vssd1 vccd1 vccd1 _09640_/A sky130_fd_sc_hd__inv_2
XFILLER_28_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_204_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17412__S _17534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12650_ _12650_/A vssd1 vssd1 vccd1 vccd1 _12650_/X sky130_fd_sc_hd__clkbuf_2
XPHY_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_247_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_230_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11601_ _19569_/Q _11600_/Y _11592_/X _11583_/B vssd1 vssd1 vccd1 vccd1 _19569_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12581_ _19043_/Q _12576_/X _12408_/X _12577_/X vssd1 vssd1 vccd1 vccd1 _19043_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10865__A hold264/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14320_ _14320_/A vssd1 vssd1 vccd1 vccd1 _14320_/X sky130_fd_sc_hd__clkbuf_2
XPHY_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11532_ _11532_/A vssd1 vssd1 vccd1 vccd1 _11532_/Y sky130_fd_sc_hd__inv_2
XPHY_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17810__S0 _17918_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14251_ _14251_/A vssd1 vssd1 vccd1 vccd1 _14252_/A sky130_fd_sc_hd__inv_2
XFILLER_139_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09405__C1 _09404_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11463_ _11463_/A _11463_/B vssd1 vssd1 vccd1 vccd1 _11535_/A sky130_fd_sc_hd__or2_1
XANTENNA__19951__RESET_B repeater244/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13202_ _13202_/A vssd1 vssd1 vccd1 vccd1 _13202_/X sky130_fd_sc_hd__clkbuf_4
X_10414_ _14245_/A _15821_/B _10430_/A vssd1 vssd1 vccd1 vccd1 _15826_/A sky130_fd_sc_hd__or3_4
X_14182_ _19118_/Q _14027_/A _19112_/Q _14021_/A vssd1 vssd1 vccd1 vccd1 _14182_/X
+ sky130_fd_sc_hd__o22a_1
X_11394_ _11625_/A _19135_/Q _19555_/Q _11393_/Y vssd1 vssd1 vccd1 vccd1 _11394_/X
+ sky130_fd_sc_hd__o22a_1
X_13133_ _19181_/Q _13082_/A _13132_/Y _18899_/Q vssd1 vssd1 vccd1 vccd1 _13133_/X
+ sky130_fd_sc_hd__o22a_1
X_10345_ _10354_/A vssd1 vssd1 vccd1 vccd1 _10345_/X sky130_fd_sc_hd__clkbuf_2
X_18990_ _19115_/CLK _18990_/D hold273/X vssd1 vssd1 vccd1 vccd1 _18990_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_151_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_128_HCLK_A clkbuf_4_4_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17941_ _19842_/CLK _17941_/D vssd1 vssd1 vccd1 vccd1 _17941_/Q sky130_fd_sc_hd__dfxtp_1
X_13064_ _13064_/A _13064_/B vssd1 vssd1 vccd1 vccd1 _13207_/A sky130_fd_sc_hd__or2_1
X_10276_ _14317_/B _10275_/Y _14317_/B _10275_/Y vssd1 vssd1 vccd1 vccd1 _10281_/C
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_78_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12015_ _19353_/Q _12009_/X _09039_/X _12010_/X vssd1 vssd1 vccd1 vccd1 _19353_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_238_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17872_ _16160_/Y _16161_/Y _16162_/Y _16163_/Y _17913_/S0 _19632_/Q vssd1 vssd1
+ vccd1 vccd1 _17872_/X sky130_fd_sc_hd__mux4_1
XANTENNA__17877__S0 _17908_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrepeater209 repeater210/X vssd1 vssd1 vccd1 vccd1 repeater209/X sky130_fd_sc_hd__buf_6
X_19611_ _19771_/CLK _19611_/D repeater190/X vssd1 vssd1 vccd1 vccd1 _19611_/Q sky130_fd_sc_hd__dfrtp_1
X_16823_ _16822_/X _09418_/Y _17529_/S vssd1 vssd1 vccd1 vccd1 _16823_/X sky130_fd_sc_hd__mux2_1
XANTENNA__08931__B2 _08930_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19542_ _19544_/CLK _19542_/D repeater221/X vssd1 vssd1 vccd1 vccd1 _19542_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_171_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16754_ vssd1 vssd1 vccd1 vccd1 _16926_/A1 _16754_/LO sky130_fd_sc_hd__conb_1
X_13966_ _13966_/A _13966_/B _13970_/C vssd1 vssd1 vccd1 vccd1 _18707_/D sky130_fd_sc_hd__nor3_1
XFILLER_0_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15705_ _10314_/B _15704_/X _15673_/X vssd1 vssd1 vccd1 vccd1 _15705_/X sky130_fd_sc_hd__o21a_1
X_12917_ _19280_/Q vssd1 vssd1 vccd1 vccd1 _12917_/Y sky130_fd_sc_hd__inv_1
X_16685_ _16962_/X _16633_/X _16924_/X _16634_/X vssd1 vssd1 vccd1 vccd1 _16685_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_19_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19473_ _19515_/CLK hold201/X repeater260/X vssd1 vssd1 vccd1 vccd1 _19473_/Q sky130_fd_sc_hd__dfrtp_1
X_13897_ _13885_/X _13897_/B _13897_/C _13897_/D vssd1 vssd1 vccd1 vccd1 _13898_/D
+ sky130_fd_sc_hd__and4b_1
XANTENNA__17322__S _17523_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18424_ _18441_/CLK _18424_/D vssd1 vssd1 vccd1 vccd1 _18424_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14768__B1 _14691_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12848_ _18936_/Q vssd1 vssd1 vccd1 vccd1 _12878_/A sky130_fd_sc_hd__inv_2
X_15636_ _15640_/B vssd1 vssd1 vccd1 vccd1 _15642_/B sky130_fd_sc_hd__inv_2
XFILLER_222_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18355_ _18465_/CLK _18355_/D vssd1 vssd1 vccd1 vccd1 _18355_/Q sky130_fd_sc_hd__dfxtp_1
X_15567_ _18584_/Q _15562_/A _18585_/Q vssd1 vssd1 vccd1 vccd1 _15567_/X sky130_fd_sc_hd__o21a_1
X_12779_ _19237_/Q vssd1 vssd1 vccd1 vccd1 _12779_/Y sky130_fd_sc_hd__inv_2
XPHY_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14518_ _14519_/A vssd1 vssd1 vccd1 vccd1 _14518_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_17306_ _17305_/X _14065_/Y _17544_/S vssd1 vssd1 vccd1 vccd1 _17306_/X sky130_fd_sc_hd__mux2_1
XANTENNA__17801__S0 _17918_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18286_ _19847_/CLK _18286_/D vssd1 vssd1 vccd1 vccd1 _18286_/Q sky130_fd_sc_hd__dfxtp_1
X_15498_ _15498_/A vssd1 vssd1 vccd1 vccd1 _15498_/Y sky130_fd_sc_hd__inv_2
XFILLER_159_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17237_ _16590_/Y _15645_/Y _17318_/S vssd1 vssd1 vccd1 vccd1 _17237_/X sky130_fd_sc_hd__mux2_2
X_14449_ _18370_/Q _14438_/A _14405_/X _14439_/A vssd1 vssd1 vccd1 vccd1 _18370_/D
+ sky130_fd_sc_hd__a22o_1
X_17168_ _17473_/A0 _16561_/Y _17547_/S vssd1 vssd1 vccd1 vccd1 _17168_/X sky130_fd_sc_hd__mux2_1
XFILLER_116_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16119_ _19369_/Q vssd1 vssd1 vccd1 vccd1 _16119_/Y sky130_fd_sc_hd__inv_2
XFILLER_115_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17099_ _15963_/X _09509_/Y _17534_/S vssd1 vssd1 vccd1 vccd1 _17099_/X sky130_fd_sc_hd__mux2_1
X_09990_ _09990_/A vssd1 vssd1 vccd1 vccd1 _09990_/X sky130_fd_sc_hd__buf_2
XFILLER_142_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08941_ _18774_/Q vssd1 vssd1 vccd1 vccd1 _08941_/Y sky130_fd_sc_hd__inv_2
XFILLER_170_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09175__B2 _09165_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17868__S0 _17908_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_218_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19809_ _19810_/CLK _19809_/D repeater224/X vssd1 vssd1 vccd1 vccd1 _19809_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__19985__CLK _19992_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18574__RESET_B repeater272/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_225_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16637__A _16637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_225_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17232__S _17459_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09424_ _19377_/Q vssd1 vssd1 vccd1 vccd1 _09424_/Y sky130_fd_sc_hd__inv_2
XFILLER_240_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_213_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_212_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09355_ _20022_/Q vssd1 vssd1 vccd1 vccd1 _09482_/A sky130_fd_sc_hd__inv_2
XFILLER_12_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_212_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10685__A _19500_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09286_ _09293_/A vssd1 vssd1 vccd1 vccd1 _09294_/A sky130_fd_sc_hd__inv_2
XFILLER_139_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_176_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15184__B1 _10446_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19362__RESET_B hold370/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_180_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10130_ _17927_/Q _10130_/B vssd1 vssd1 vccd1 vccd1 _10130_/X sky130_fd_sc_hd__and2_1
XFILLER_79_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10061_ _10046_/A _10046_/B _10032_/A _10059_/Y vssd1 vssd1 vccd1 vccd1 _19930_/D
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__09166__B2 _09165_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17407__S _17517_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17859__S0 _18760_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_197_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12170__B1 _11975_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13820_ _13910_/B _13935_/A vssd1 vssd1 vccd1 vccd1 _13821_/B sky130_fd_sc_hd__or2_2
XFILLER_29_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_115_HCLK clkbuf_opt_0_HCLK/A vssd1 vssd1 vccd1 vccd1 _19115_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_62_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_244_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13751_ _13751_/A vssd1 vssd1 vccd1 vccd1 _17763_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_28_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10963_ _10963_/A _10987_/A vssd1 vssd1 vccd1 vccd1 _10983_/A sky130_fd_sc_hd__or2_1
XFILLER_90_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16739__B2 _16512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13670__B1 _12599_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_244_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_231_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17142__S _17493_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12702_ _18964_/Q _12698_/X _12533_/X _12699_/X vssd1 vssd1 vccd1 vccd1 _18964_/D
+ sky130_fd_sc_hd__a22o_1
X_16470_ _16616_/A vssd1 vssd1 vccd1 vccd1 _16544_/B sky130_fd_sc_hd__buf_4
X_13682_ _14405_/A vssd1 vssd1 vccd1 vccd1 _13682_/X sky130_fd_sc_hd__buf_2
X_10894_ _10894_/A vssd1 vssd1 vccd1 vccd1 _10895_/A sky130_fd_sc_hd__inv_2
XFILLER_71_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15421_ _19612_/Q _19611_/Q _11158_/B vssd1 vssd1 vccd1 vccd1 _15421_/X sky130_fd_sc_hd__a21bo_1
XPHY_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12633_ _19011_/Q _12629_/X _12406_/X _12630_/X vssd1 vssd1 vccd1 vccd1 _19011_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15352_ _15358_/A _17593_/X vssd1 vssd1 vccd1 vccd1 _18497_/D sky130_fd_sc_hd__and2_1
XPHY_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18140_ _19851_/CLK _18140_/D vssd1 vssd1 vccd1 vccd1 _18140_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_196_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12564_ _19056_/Q _12560_/X _12375_/X _12563_/X vssd1 vssd1 vccd1 vccd1 _19056_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11984__B1 _11920_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14303_ _14304_/A vssd1 vssd1 vccd1 vccd1 _14303_/X sky130_fd_sc_hd__clkbuf_2
XPHY_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11515_ _19595_/Q _11514_/Y _11504_/X _11476_/B vssd1 vssd1 vccd1 vccd1 _19595_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18071_ _18169_/CLK _18071_/D vssd1 vssd1 vccd1 vccd1 _18071_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15283_ _15283_/A vssd1 vssd1 vccd1 vccd1 _15439_/A sky130_fd_sc_hd__clkbuf_2
XPHY_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15175__B1 hold244/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12495_ _19090_/Q _12489_/X _12382_/X _12492_/X vssd1 vssd1 vccd1 vccd1 _19090_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_200_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17022_ _17486_/A0 _13097_/Y _17543_/S vssd1 vssd1 vccd1 vccd1 _17022_/X sky130_fd_sc_hd__mux2_1
X_14234_ _14236_/A vssd1 vssd1 vccd1 vccd1 _14235_/A sky130_fd_sc_hd__inv_2
XFILLER_184_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_184_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11446_ _19154_/Q vssd1 vssd1 vccd1 vccd1 _11446_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19032__RESET_B repeater269/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14165_ _19105_/Q _14014_/A _19093_/Q _14003_/A _14164_/X vssd1 vssd1 vccd1 vccd1
+ _14166_/D sky130_fd_sc_hd__o221a_1
X_11377_ _11622_/A _19132_/Q _11584_/C _19152_/Q _11376_/X vssd1 vssd1 vccd1 vccd1
+ _11389_/B sky130_fd_sc_hd__o221a_1
XFILLER_180_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13116_ _13115_/Y _18913_/Q _19169_/Q _13070_/A vssd1 vssd1 vccd1 vccd1 _13116_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_180_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10328_ _10328_/A _10352_/A vssd1 vssd1 vccd1 vccd1 _10348_/A sky130_fd_sc_hd__or2_1
XFILLER_112_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18973_ _19597_/CLK _18973_/D repeater282/X vssd1 vssd1 vccd1 vccd1 _18973_/Q sky130_fd_sc_hd__dfrtp_2
X_14096_ _14112_/A vssd1 vssd1 vccd1 vccd1 _14096_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__17317__S _17473_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17924_ _17920_/X _17921_/X _17922_/X _17923_/X _19647_/Q _19648_/Q vssd1 vssd1 vccd1
+ vccd1 _17924_/X sky130_fd_sc_hd__mux4_2
X_13047_ _18899_/Q vssd1 vssd1 vccd1 vccd1 _13071_/A sky130_fd_sc_hd__inv_2
X_10259_ _11029_/A vssd1 vssd1 vccd1 vccd1 _17753_/S sky130_fd_sc_hd__inv_2
XFILLER_59_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12161__B1 _12028_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11873__B _11998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17855_ _16275_/Y _16276_/Y _16277_/Y _16278_/Y _17908_/S0 _18759_/Q vssd1 vssd1
+ vccd1 vccd1 _17855_/X sky130_fd_sc_hd__mux4_2
XFILLER_38_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16978__A1 _19146_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16806_ _16805_/X _13086_/A _17488_/S vssd1 vssd1 vccd1 vccd1 _16806_/X sky130_fd_sc_hd__mux2_1
XANTENNA__14989__B1 _14782_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_208_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17786_ _18390_/Q _18382_/Q _18374_/Q _18366_/Q _17923_/S0 _19646_/Q vssd1 vssd1
+ vccd1 vccd1 _17786_/X sky130_fd_sc_hd__mux4_2
XFILLER_226_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14998_ _18957_/Q vssd1 vssd1 vccd1 vccd1 _14998_/X sky130_fd_sc_hd__buf_2
XFILLER_82_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19525_ _19771_/CLK _19525_/D repeater190/X vssd1 vssd1 vccd1 vccd1 _19525_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__11267__A2 _19012_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16737_ _19470_/Q vssd1 vssd1 vccd1 vccd1 _16737_/Y sky130_fd_sc_hd__inv_2
XFILLER_241_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13661__B1 _12030_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13949_ _13949_/A _13949_/B vssd1 vssd1 vccd1 vccd1 _13954_/A sky130_fd_sc_hd__or2_1
XFILLER_34_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17052__S _17522_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19456_ _19462_/CLK _19456_/D repeater272/X vssd1 vssd1 vccd1 vccd1 _19456_/Q sky130_fd_sc_hd__dfrtp_1
X_16668_ _16668_/A _16668_/B vssd1 vssd1 vccd1 vccd1 _16668_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__16176__B _16344_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18407_ _18959_/CLK _18407_/D vssd1 vssd1 vccd1 vccd1 _18407_/Q sky130_fd_sc_hd__dfxtp_1
X_15619_ _15622_/B _15618_/Y _15614_/X vssd1 vssd1 vccd1 vccd1 _15619_/X sky130_fd_sc_hd__o21a_1
X_19387_ _19927_/CLK _19387_/D repeater235/X vssd1 vssd1 vccd1 vccd1 _19387_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__16891__S _17545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16599_ _17250_/X _16597_/X _17245_/X _16598_/X vssd1 vssd1 vccd1 vccd1 _16600_/D
+ sky130_fd_sc_hd__a22o_2
X_09140_ _13494_/A _15321_/B hold344/X _17602_/X vssd1 vssd1 vccd1 vccd1 _09140_/Y
+ sky130_fd_sc_hd__a31oi_2
X_18338_ _18954_/CLK _18338_/D vssd1 vssd1 vccd1 vccd1 _18338_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17155__A1 _08930_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09071_ hold239/X vssd1 vssd1 vccd1 vccd1 _09071_/X sky130_fd_sc_hd__buf_4
XANTENNA__16902__A1 _20099_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18269_ _20076_/CLK _18269_/D vssd1 vssd1 vccd1 vccd1 _18269_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13177__C1 _13176_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_190_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12225__A hold260/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09973_ _19958_/Q _09972_/Y _09968_/X _09867_/B vssd1 vssd1 vccd1 vccd1 _19958_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__17227__S _17318_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08924_ _18783_/Q vssd1 vssd1 vccd1 vccd1 _08924_/Y sky130_fd_sc_hd__inv_2
X_20093_ _20107_/CLK _20093_/D repeater233/X vssd1 vssd1 vccd1 vccd1 _20093_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_clkbuf_leaf_111_HCLK_A clkbuf_opt_0_HCLK/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18755__RESET_B repeater195/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12152__B1 _12095_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_138_HCLK clkbuf_4_3_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _20058_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_245_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_233_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_226_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_226_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_241_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_198_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09407_ _19375_/Q vssd1 vssd1 vccd1 vccd1 _09407_/Y sky130_fd_sc_hd__inv_2
XFILLER_71_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13404__B1 _20105_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_201_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_187_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09338_ _17622_/X _13766_/D _20038_/Q _15727_/B vssd1 vssd1 vccd1 vccd1 _20038_/D
+ sky130_fd_sc_hd__o22a_1
XANTENNA__19543__RESET_B repeater221/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_178_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_178_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11966__B1 _09061_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09269_ _09270_/A vssd1 vssd1 vccd1 vccd1 _09269_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_194_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11300_ _18987_/Q vssd1 vssd1 vccd1 vccd1 _11300_/Y sky130_fd_sc_hd__inv_2
XFILLER_153_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12280_ _19212_/Q _12276_/X _12100_/X _12277_/X vssd1 vssd1 vccd1 vccd1 _19212_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_112_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11231_ _19607_/Q vssd1 vssd1 vccd1 vccd1 _11487_/A sky130_fd_sc_hd__inv_2
XFILLER_181_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12391__B1 _12389_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11162_ _19617_/Q _11162_/B vssd1 vssd1 vccd1 vccd1 _11163_/B sky130_fd_sc_hd__or2_1
XFILLER_150_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17137__S _17513_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10113_ _18560_/Q _15457_/A vssd1 vssd1 vccd1 vccd1 _15462_/A sky130_fd_sc_hd__or2_1
XANTENNA__15446__A _15479_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15970_ _19710_/Q vssd1 vssd1 vccd1 vccd1 _15970_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14350__A hold248/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11093_ _19639_/Q vssd1 vssd1 vccd1 vccd1 _11093_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18496__RESET_B repeater203/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10044_ _10044_/A _10044_/B vssd1 vssd1 vccd1 vccd1 _10062_/A sky130_fd_sc_hd__or2_1
X_14921_ _20081_/Q vssd1 vssd1 vccd1 vccd1 _14921_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_102_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16976__S _17545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17082__A0 _17473_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17640_ _15679_/X _19049_/Q _17655_/S vssd1 vssd1 vccd1 vccd1 _18612_/D sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_33_HCLK_A _18641_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14852_ _18141_/Q _14845_/X _14812_/X _14847_/X vssd1 vssd1 vccd1 vccd1 _18141_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_75_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_96_HCLK_A clkbuf_4_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13803_ _18711_/Q vssd1 vssd1 vccd1 vccd1 _13948_/A sky130_fd_sc_hd__inv_2
XFILLER_223_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17571_ _15418_/X _19772_/Q _17584_/S vssd1 vssd1 vccd1 vccd1 _17571_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12446__A1 _19123_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14783_ _18178_/Q _14772_/A _14782_/X _14773_/A vssd1 vssd1 vccd1 vccd1 _18178_/D
+ sky130_fd_sc_hd__a22o_1
X_11995_ _11991_/X _19363_/Q _11995_/S vssd1 vssd1 vccd1 vccd1 _19363_/D sky130_fd_sc_hd__mux2_1
XANTENNA_output119_A _16750_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19310_ _20032_/CLK _19310_/D repeater240/X vssd1 vssd1 vccd1 vccd1 _19310_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_72_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10457__B1 _10425_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13734_ _13733_/A _14392_/A _18754_/Q _13733_/Y vssd1 vssd1 vccd1 vccd1 _18754_/D
+ sky130_fd_sc_hd__o22a_1
X_16522_ _17269_/X _15896_/X _17301_/X _16493_/X vssd1 vssd1 vccd1 vccd1 _16522_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_216_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10946_ hold266/X hold368/A vssd1 vssd1 vccd1 vccd1 _10949_/A sky130_fd_sc_hd__nand2_4
XANTENNA__17385__A1 _20095_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_231_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_188_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19241_ _19314_/CLK _19241_/D repeater239/X vssd1 vssd1 vccd1 vccd1 _19241_/Q sky130_fd_sc_hd__dfrtp_4
X_16453_ _18516_/Q vssd1 vssd1 vccd1 vccd1 _16453_/Y sky130_fd_sc_hd__inv_2
X_13665_ _13672_/A vssd1 vssd1 vccd1 vccd1 _13665_/X sky130_fd_sc_hd__buf_1
XFILLER_188_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_repeater171_A _17482_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10877_ _14273_/A vssd1 vssd1 vccd1 vccd1 _10877_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_176_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17600__S _17600_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15404_ _15404_/A vssd1 vssd1 vccd1 vccd1 _15413_/A sky130_fd_sc_hd__clkbuf_2
X_12616_ _12630_/A vssd1 vssd1 vccd1 vccd1 _12616_/X sky130_fd_sc_hd__buf_1
X_16384_ _19771_/Q vssd1 vssd1 vccd1 vccd1 _16384_/Y sky130_fd_sc_hd__inv_2
X_19172_ _19208_/CLK _19172_/D hold367/X vssd1 vssd1 vccd1 vccd1 _19172_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13596_ _13537_/B _13596_/A2 _13537_/A vssd1 vssd1 vccd1 vccd1 _13597_/C sky130_fd_sc_hd__o21a_1
XPHY_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_19_HCLK clkbuf_4_3_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19900_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11957__B1 hold314/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15335_ _19703_/Q vssd1 vssd1 vccd1 vccd1 _15335_/Y sky130_fd_sc_hd__inv_2
X_18123_ _18260_/CLK _18123_/D vssd1 vssd1 vccd1 vccd1 _18123_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__18642__D _18642_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12547_ _12551_/C vssd1 vssd1 vccd1 vccd1 _12556_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_157_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_177_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15266_ _15311_/A _15266_/B vssd1 vssd1 vccd1 vccd1 _15266_/X sky130_fd_sc_hd__or2_1
X_18054_ _18142_/CLK _18054_/D vssd1 vssd1 vccd1 vccd1 _18054_/Q sky130_fd_sc_hd__dfxtp_1
X_12478_ _12478_/A vssd1 vssd1 vccd1 vccd1 _12478_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_8_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20118__RESET_B repeater217/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14217_ _19110_/Q _14019_/A _16666_/A _18696_/Q _14216_/X vssd1 vssd1 vccd1 vccd1
+ _14218_/D sky130_fd_sc_hd__o221a_1
XFILLER_6_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17005_ _17473_/A0 _16608_/Y _17512_/S vssd1 vssd1 vccd1 vccd1 _17005_/X sky130_fd_sc_hd__mux2_1
XFILLER_160_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11429_ _19140_/Q vssd1 vssd1 vccd1 vccd1 _11429_/Y sky130_fd_sc_hd__inv_2
X_15197_ _15197_/A vssd1 vssd1 vccd1 vccd1 _17567_/S sky130_fd_sc_hd__clkinv_8
XFILLER_98_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14148_ _14148_/A vssd1 vssd1 vccd1 vccd1 _14148_/Y sky130_fd_sc_hd__clkinvlp_2
XANTENNA__17047__S _17490_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11884__A _11891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14079_ _19082_/Q _14023_/A _19078_/Q _14019_/A _14078_/X vssd1 vssd1 vccd1 vccd1
+ _14080_/D sky130_fd_sc_hd__o221a_1
X_18956_ _18959_/CLK _18956_/D repeater257/X vssd1 vssd1 vccd1 vccd1 _18956_/Q sky130_fd_sc_hd__dfrtp_1
X_17907_ _15810_/Y _15811_/Y _15812_/Y _15813_/Y _17908_/S0 _18759_/Q vssd1 vssd1
+ vccd1 vccd1 _17907_/X sky130_fd_sc_hd__mux4_1
XFILLER_239_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16886__S _17513_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18887_ _19288_/CLK _18887_/D repeater212/X vssd1 vssd1 vccd1 vccd1 _18887_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_227_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17838_ _16429_/Y _16430_/Y _16431_/Y _16432_/Y _17908_/S0 _18759_/Q vssd1 vssd1
+ vccd1 vccd1 _17838_/X sky130_fd_sc_hd__mux4_2
Xrebuffer15 _14014_/B vssd1 vssd1 vccd1 vccd1 _14131_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_67_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_208_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrebuffer26 _13061_/B vssd1 vssd1 vccd1 vccd1 _13215_/B1 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_66_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrebuffer37 _19418_/Q vssd1 vssd1 vccd1 vccd1 _17246_/A1 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer48 _13551_/B vssd1 vssd1 vccd1 vccd1 _13572_/A2 sky130_fd_sc_hd__dlygate4sd1_1
X_17769_ _17765_/X _17766_/X _17767_/X _17768_/X _19647_/Q _19648_/Q vssd1 vssd1 vccd1
+ vccd1 _17769_/X sky130_fd_sc_hd__mux4_2
XFILLER_212_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xrebuffer59 _09388_/B2 vssd1 vssd1 vccd1 vccd1 _16963_/A1 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_47_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19508_ _19510_/CLK hold214/X repeater256/X vssd1 vssd1 vccd1 vccd1 _19508_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_81_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_212_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19439_ _20066_/CLK _19439_/D repeater193/X vssd1 vssd1 vccd1 vccd1 _19439_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_223_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_211_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17510__S _17548_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_195_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_176_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09123_ _20084_/Q vssd1 vssd1 vccd1 vccd1 _09144_/C sky130_fd_sc_hd__inv_2
XFILLER_148_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrebuffer105 _13536_/B vssd1 vssd1 vccd1 vccd1 _13602_/C1 sky130_fd_sc_hd__dlygate4sd1_1
XANTENNA__15139__B1 hold244/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrebuffer116 _13532_/B vssd1 vssd1 vccd1 vccd1 _13608_/C1 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer127 _12968_/B vssd1 vssd1 vccd1 vccd1 rebuffer1/A sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_176_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16887__A0 _17473_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09054_ hold277/X vssd1 vssd1 vccd1 vccd1 hold276/A sky130_fd_sc_hd__buf_6
XFILLER_136_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18158__CLK _18198_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_237_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19403__CLK _19984_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11794__A _11801_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09956_ _09875_/A _09956_/A2 _09954_/Y _09987_/B vssd1 vssd1 vccd1 vccd1 _19967_/D
+ sky130_fd_sc_hd__a211oi_4
XANTENNA__12125__B1 _11918_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16796__S _17534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09887_ _19345_/Q vssd1 vssd1 vccd1 vccd1 _16548_/A sky130_fd_sc_hd__inv_2
X_20076_ _20076_/CLK _20076_/D repeater196/X vssd1 vssd1 vccd1 vccd1 _20076_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_245_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19795__RESET_B repeater219/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10800_ _19733_/Q _10800_/B vssd1 vssd1 vccd1 vccd1 _10801_/B sky130_fd_sc_hd__nand2_1
XANTENNA__10439__B1 _09067_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_226_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11780_ _12130_/A _12370_/B _12130_/C vssd1 vssd1 vccd1 vccd1 _16238_/A sky130_fd_sc_hd__or3_4
XPHY_3834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_241_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_213_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10731_ _11651_/A _11651_/B _17608_/X vssd1 vssd1 vccd1 vccd1 _15270_/C sky130_fd_sc_hd__or3b_1
XPHY_3856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15917__A2 _15908_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_241_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17420__S _17488_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13450_ _13450_/A vssd1 vssd1 vccd1 vccd1 _13450_/Y sky130_fd_sc_hd__inv_2
XFILLER_185_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10662_ _10676_/A vssd1 vssd1 vccd1 vccd1 _10677_/A sky130_fd_sc_hd__inv_2
XFILLER_167_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_201_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12401_ hold315/X vssd1 vssd1 vccd1 vccd1 _12401_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__16544__B _16544_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11969__A _11977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13381_ _20099_/Q _18845_/Q _20099_/Q _18845_/Q vssd1 vssd1 vccd1 vccd1 _13381_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_10593_ _19800_/Q _10593_/B _19799_/Q vssd1 vssd1 vccd1 vccd1 _10594_/C sky130_fd_sc_hd__nor3b_2
XANTENNA__10873__A _16053_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15120_ _17977_/Q _15111_/A _14949_/X _15112_/A vssd1 vssd1 vccd1 vccd1 _17977_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_194_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12332_ _19181_/Q _12327_/X _12090_/X _12328_/X vssd1 vssd1 vccd1 vccd1 _19181_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_31_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15051_ _18024_/Q _15047_/X _14996_/X _15049_/X vssd1 vssd1 vccd1 vccd1 _18024_/D
+ sky130_fd_sc_hd__a22o_1
X_12263_ _12277_/A vssd1 vssd1 vccd1 vccd1 _12263_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__18677__RESET_B repeater252/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14002_ _18672_/Q vssd1 vssd1 vccd1 vccd1 _14003_/A sky130_fd_sc_hd__inv_2
XANTENNA__12364__B1 _12302_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_181_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13561__C1 _13560_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11214_ _19011_/Q vssd1 vssd1 vccd1 vccd1 _11214_/Y sky130_fd_sc_hd__inv_2
XFILLER_141_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12194_ _19257_/Q _12189_/X _12074_/X _12192_/X vssd1 vssd1 vccd1 vccd1 _19257_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_134_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18810_ _20115_/CLK _18810_/D repeater217/X vssd1 vssd1 vccd1 vccd1 _18810_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_1_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11145_ _19629_/Q _11144_/Y _11141_/X vssd1 vssd1 vccd1 vccd1 _19629_/D sky130_fd_sc_hd__o21a_1
X_19790_ _20089_/CLK _19790_/D repeater203/X vssd1 vssd1 vccd1 vccd1 _19790_/Q sky130_fd_sc_hd__dfrtp_1
Xoutput84 _16559_/Y vssd1 vssd1 vccd1 vccd1 HRDATA[14] sky130_fd_sc_hd__clkbuf_2
Xoutput95 _16678_/X vssd1 vssd1 vccd1 vccd1 HRDATA[24] sky130_fd_sc_hd__clkbuf_2
XFILLER_89_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12116__B1 _12035_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18741_ _20066_/CLK _18741_/D repeater209/X vssd1 vssd1 vccd1 vccd1 _18741_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__12667__A1 _18989_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11076_ _11076_/A _11076_/B _11076_/C _11103_/A vssd1 vssd1 vccd1 vccd1 _11076_/X
+ sky130_fd_sc_hd__or4b_1
X_15953_ _18083_/Q vssd1 vssd1 vccd1 vccd1 _15953_/Y sky130_fd_sc_hd__inv_2
XFILLER_237_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_236_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10027_ _19937_/Q _10032_/B _09425_/Y _10024_/A _10026_/X vssd1 vssd1 vccd1 vccd1
+ _19937_/D sky130_fd_sc_hd__o221a_1
X_14904_ _18108_/Q _14897_/A _14711_/X _14898_/A vssd1 vssd1 vccd1 vccd1 _18108_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_237_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18672_ _18686_/CLK _18672_/D repeater252/X vssd1 vssd1 vccd1 vccd1 _18672_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_64_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_248_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15884_ _15884_/A vssd1 vssd1 vccd1 vccd1 _15884_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_76_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16719__B _16721_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17623_ _10789_/Y _10786_/Y _18653_/Q vssd1 vssd1 vccd1 vccd1 _18653_/D sky130_fd_sc_hd__mux2_1
X_14835_ _18153_/Q _14832_/X _14802_/X _14834_/X vssd1 vssd1 vccd1 vccd1 _18153_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__15081__A2 _15072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19465__RESET_B repeater274/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17554_ _17553_/X _20058_/Q _17558_/S vssd1 vssd1 vccd1 vccd1 _17554_/X sky130_fd_sc_hd__mux2_1
XFILLER_205_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_189_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14766_ _18189_/Q _14759_/X _14725_/X _14761_/X vssd1 vssd1 vccd1 vccd1 _18189_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_91_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11978_ _14277_/A vssd1 vssd1 vccd1 vccd1 _11978_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__09296__B1 _09098_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13631__A3 _19873_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16505_ _16505_/A vssd1 vssd1 vccd1 vccd1 _16505_/X sky130_fd_sc_hd__clkbuf_2
X_10929_ _17725_/X _10923_/X _19676_/Q _10924_/X vssd1 vssd1 vccd1 vccd1 _19676_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_60_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13717_ _18760_/Q _13710_/B _13706_/B vssd1 vssd1 vccd1 vccd1 _13717_/Y sky130_fd_sc_hd__o21ai_1
X_17485_ _17484_/X _13529_/A _17536_/S vssd1 vssd1 vccd1 vccd1 _17485_/X sky130_fd_sc_hd__mux2_4
X_14697_ _15121_/A _15145_/B _15121_/C vssd1 vssd1 vccd1 vccd1 _14700_/A sky130_fd_sc_hd__or3_4
XFILLER_32_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17330__S _17543_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19224_ _19224_/CLK _19224_/D repeater186/X vssd1 vssd1 vccd1 vccd1 _19224_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__09048__B1 hold317/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10850__B1 _10421_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16436_ _20066_/Q _16436_/B vssd1 vssd1 vccd1 vccd1 _16436_/Y sky130_fd_sc_hd__nand2_1
XFILLER_158_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14041__B1 _19084_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13648_ _16956_/X _13644_/X _18793_/Q _13646_/X vssd1 vssd1 vccd1 vccd1 _18793_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_13_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19155_ _19577_/CLK _19155_/D repeater268/X vssd1 vssd1 vccd1 vccd1 _19155_/Q sky130_fd_sc_hd__dfrtp_2
X_13579_ _13547_/A _13547_/B _13571_/X _13577_/Y vssd1 vssd1 vccd1 vccd1 _18824_/D
+ sky130_fd_sc_hd__a211oi_2
X_16367_ _16437_/A _18743_/Q vssd1 vssd1 vccd1 vccd1 _16367_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__10783__A _20036_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18106_ _18260_/CLK _18106_/D vssd1 vssd1 vccd1 vccd1 _18106_/Q sky130_fd_sc_hd__dfxtp_1
X_15318_ _15318_/A _15318_/B vssd1 vssd1 vccd1 vccd1 _15318_/Y sky130_fd_sc_hd__nor2_1
XFILLER_157_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19086_ _19119_/CLK _19086_/D hold351/X vssd1 vssd1 vccd1 vccd1 _19086_/Q sky130_fd_sc_hd__dfrtp_2
X_16298_ _16437_/A _18742_/Q vssd1 vssd1 vccd1 vccd1 _16298_/Y sky130_fd_sc_hd__nand2_1
XFILLER_184_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18037_ _19851_/CLK _18037_/D vssd1 vssd1 vccd1 vccd1 _18037_/Q sky130_fd_sc_hd__dfxtp_1
X_15249_ _18519_/Q vssd1 vssd1 vccd1 vccd1 _15437_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__12355__B1 _12353_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17294__A0 _17486_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09810_ _09810_/A vssd1 vssd1 vccd1 vccd1 _09813_/A sky130_fd_sc_hd__inv_2
X_19988_ _19992_/CLK _19988_/D repeater192/X vssd1 vssd1 vccd1 vccd1 _19988_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_140_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09084__A _09084_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09741_ _09741_/A _09784_/A vssd1 vssd1 vccd1 vccd1 _09742_/B sky130_fd_sc_hd__or2_2
X_18939_ _19325_/CLK _18939_/D repeater213/X vssd1 vssd1 vccd1 vccd1 _18939_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_98_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17046__A0 _15768_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17505__S _17565_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09672_ _19407_/Q vssd1 vssd1 vccd1 vccd1 _09672_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11330__B2 _11328_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16629__B _16629_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_199_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_242_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14280__B1 _14279_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_223_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_211_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17240__S _17548_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10693__A _10704_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09106_ _20092_/Q _09041_/A _09105_/X _09043_/A vssd1 vssd1 vccd1 vccd1 _20092_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12594__B1 hold267/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_184_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09037_ hold296/X vssd1 vssd1 vccd1 vccd1 _09037_/X sky130_fd_sc_hd__buf_4
XANTENNA__18770__RESET_B repeater271/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold350 hold350/A vssd1 vssd1 vccd1 vccd1 hold367/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold361 hold361/A vssd1 vssd1 vccd1 vccd1 hold361/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17285__A0 _15768_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold372 hold372/A vssd1 vssd1 vccd1 vccd1 hold372/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12413__A hold277/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09939_ _19356_/Q vssd1 vssd1 vccd1 vccd1 _09939_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19976__RESET_B repeater244/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_219_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12132__B _12316_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17415__S _17534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12950_ _19277_/Q _12876_/A _12948_/Y _18934_/Q _12949_/Y vssd1 vssd1 vccd1 vccd1
+ _12955_/C sky130_fd_sc_hd__o221a_1
XFILLER_219_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20059_ _20059_/CLK _20059_/D repeater197/X vssd1 vssd1 vccd1 vccd1 _20059_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_218_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11901_ _19416_/Q _11898_/X _09058_/X _11899_/X vssd1 vssd1 vccd1 vccd1 _19416_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_45_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_206_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12881_ _12964_/B _12881_/B vssd1 vssd1 vccd1 vccd1 _12983_/A sky130_fd_sc_hd__or2_1
XPHY_4310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_245_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14620_ _18272_/Q _14616_/X _09171_/X _14618_/X vssd1 vssd1 vccd1 vccd1 _18272_/D
+ sky130_fd_sc_hd__a22o_1
X_11832_ _15823_/A _11832_/B _11832_/C _19503_/Q vssd1 vssd1 vccd1 vccd1 _12309_/A
+ sky130_fd_sc_hd__or4b_4
XANTENNA__09278__B1 _09105_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_221_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_4376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14551_ _18311_/Q _14546_/X _14537_/X _14548_/X vssd1 vssd1 vccd1 vccd1 _18311_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_54_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11763_ hold168/X _11757_/X _19481_/Q _11758_/X vssd1 vssd1 vccd1 vccd1 hold170/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_42_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17150__S _17534_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10714_ _10714_/A vssd1 vssd1 vccd1 vccd1 _19774_/D sky130_fd_sc_hd__inv_2
XPHY_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13502_ _18763_/Q vssd1 vssd1 vccd1 vccd1 _14628_/A sky130_fd_sc_hd__inv_2
XPHY_3697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14482_ _18352_/Q _14478_/X _12717_/X _14480_/X vssd1 vssd1 vccd1 vccd1 _18352_/D
+ sky130_fd_sc_hd__a22o_1
X_17270_ _17473_/A0 _09901_/Y _17522_/S vssd1 vssd1 vccd1 vccd1 _17270_/X sky130_fd_sc_hd__mux2_1
X_11694_ _19527_/Q _11690_/X _10882_/X _11692_/X vssd1 vssd1 vccd1 vccd1 _19527_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17760__A1 _13491_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13433_ _13433_/A _13433_/B _13433_/C _13432_/X vssd1 vssd1 vccd1 vccd1 _13433_/X
+ sky130_fd_sc_hd__or4b_4
X_16221_ _19705_/Q vssd1 vssd1 vccd1 vccd1 _16221_/Y sky130_fd_sc_hd__inv_2
XPHY_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10645_ _19785_/Q _10645_/B vssd1 vssd1 vccd1 vccd1 _10646_/B sky130_fd_sc_hd__or2_1
XPHY_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18858__RESET_B repeater231/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12585__B1 _12413_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16152_ _18142_/Q vssd1 vssd1 vccd1 vccd1 _16152_/Y sky130_fd_sc_hd__inv_2
X_13364_ _20118_/Q _13361_/Y _20097_/Q _13466_/A _13363_/X vssd1 vssd1 vccd1 vccd1
+ _13372_/B sky130_fd_sc_hd__o221a_1
X_10576_ _19802_/Q _19801_/Q _10576_/C vssd1 vssd1 vccd1 vccd1 _10585_/C sky130_fd_sc_hd__or3_1
Xrebuffer6 _13062_/B vssd1 vssd1 vccd1 vccd1 _13212_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_166_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15103_ _17988_/Q _15096_/A _14814_/A _15097_/A vssd1 vssd1 vccd1 vccd1 _17988_/D
+ sky130_fd_sc_hd__a22o_1
X_12315_ _12313_/X _19190_/Q _12315_/S vssd1 vssd1 vccd1 vccd1 _19190_/D sky130_fd_sc_hd__mux2_1
X_16083_ _18069_/Q vssd1 vssd1 vccd1 vccd1 _16083_/Y sky130_fd_sc_hd__inv_2
XFILLER_181_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13295_ _13256_/X _13294_/Y _13256_/X _13294_/Y vssd1 vssd1 vccd1 vccd1 _13299_/C
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_108_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12337__B1 _12098_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19911_ _20006_/CLK _19911_/D repeater191/X vssd1 vssd1 vccd1 vccd1 _19911_/Q sky130_fd_sc_hd__dfrtp_1
X_15034_ _15094_/A _15034_/B _15034_/C vssd1 vssd1 vccd1 vccd1 _15036_/A sky130_fd_sc_hd__or3_4
XFILLER_181_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12246_ _19060_/Q _12246_/B vssd1 vssd1 vccd1 vccd1 _12247_/B sky130_fd_sc_hd__or2_1
XFILLER_108_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10899__B1 _10861_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19842_ _19842_/CLK _19842_/D repeater270/X vssd1 vssd1 vccd1 vccd1 _19842_/Q sky130_fd_sc_hd__dfrtp_1
X_12177_ _19264_/Q _12171_/X _11922_/X _12172_/X vssd1 vssd1 vccd1 vccd1 _19264_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_111_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11128_ _11123_/A _11064_/B _11064_/A vssd1 vssd1 vccd1 vccd1 _11128_/X sky130_fd_sc_hd__o21a_1
X_19773_ _20049_/CLK _19773_/D repeater190/X vssd1 vssd1 vccd1 vccd1 _19773_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__13837__B1 _19222_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16985_ _17829_/X _19903_/Q _16986_/S vssd1 vssd1 vccd1 vccd1 _16985_/X sky130_fd_sc_hd__mux2_1
XFILLER_209_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17325__S _17529_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18724_ _18727_/CLK _18724_/D repeater253/X vssd1 vssd1 vccd1 vccd1 _18724_/Q sky130_fd_sc_hd__dfrtp_1
X_15936_ _18227_/Q vssd1 vssd1 vccd1 vccd1 _15936_/Y sky130_fd_sc_hd__inv_2
X_11059_ _19640_/Q vssd1 vssd1 vccd1 vccd1 _11059_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_237_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18655_ _19905_/CLK _18655_/D repeater210/X vssd1 vssd1 vccd1 vccd1 _18655_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_237_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15867_ _15867_/A _15867_/B vssd1 vssd1 vccd1 vccd1 _17539_/S sky130_fd_sc_hd__nor2_8
XFILLER_92_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17606_ _10552_/B _10583_/B _19813_/Q vssd1 vssd1 vccd1 vccd1 _17606_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14818_ _18162_/Q _14803_/A _14268_/X _14804_/A vssd1 vssd1 vccd1 vccd1 _18162_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_240_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18586_ _19470_/CLK _18586_/D repeater272/X vssd1 vssd1 vccd1 vccd1 _18586_/Q sky130_fd_sc_hd__dfrtp_1
X_15798_ _19842_/Q vssd1 vssd1 vccd1 vccd1 _16747_/A sky130_fd_sc_hd__inv_2
XFILLER_224_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_205_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17537_ _15869_/Y _13021_/A _17537_/S vssd1 vssd1 vccd1 vccd1 _17537_/X sky130_fd_sc_hd__mux2_1
X_14749_ _14749_/A vssd1 vssd1 vccd1 vccd1 _14749_/X sky130_fd_sc_hd__buf_2
XFILLER_233_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_205_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17200__A0 _15963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17060__S _17386_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_177_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17468_ _16025_/Y _16024_/Y _17564_/S vssd1 vssd1 vccd1 vccd1 _17468_/X sky130_fd_sc_hd__mux2_1
X_19207_ _19208_/CLK _19207_/D hold367/X vssd1 vssd1 vccd1 vccd1 _19207_/Q sky130_fd_sc_hd__dfrtp_2
X_16419_ _17952_/Q vssd1 vssd1 vccd1 vccd1 _16419_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18599__RESET_B repeater267/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17399_ _17398_/X _17869_/X _17568_/S vssd1 vssd1 vccd1 vccd1 _17399_/X sky130_fd_sc_hd__mux2_2
X_19138_ _19470_/CLK _19138_/D repeater274/X vssd1 vssd1 vccd1 vccd1 _19138_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__09079__A hold260/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17503__A1 _17899_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_218_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19069_ _19610_/CLK _19069_/D hold361/X vssd1 vssd1 vccd1 vccd1 _19069_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_173_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17267__A0 _17486_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_234_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17990__CLK _18169_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_248_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17019__A0 _15963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09724_ _19424_/Q vssd1 vssd1 vccd1 vccd1 _09724_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17235__S _17541_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11303__B2 _18974_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12500__B1 _12389_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09655_ _19990_/Q vssd1 vssd1 vccd1 vccd1 _09746_/A sky130_fd_sc_hd__inv_2
XFILLER_227_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_242_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_227_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09261__B _15914_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09586_ _20025_/Q _09584_/Y _09585_/X _09486_/B vssd1 vssd1 vccd1 vccd1 _20025_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_83_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_242_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14253__B1 _13680_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_203_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_230_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_223_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19741__CLK _20051_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_195_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12408__A hold310/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12567__B1 _12384_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10430_ _10430_/A _16492_/A vssd1 vssd1 vccd1 vccd1 _16053_/A sky130_fd_sc_hd__or2_4
XFILLER_148_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_192_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10361_ _10361_/A _10361_/B vssd1 vssd1 vccd1 vccd1 _10361_/X sky130_fd_sc_hd__and2_1
XFILLER_128_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16702__C1 _16701_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12100_ hold318/X vssd1 vssd1 vccd1 vccd1 _12100_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_124_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13080_ _13080_/A _13179_/A vssd1 vssd1 vccd1 vccd1 _13081_/B sky130_fd_sc_hd__or2_2
X_10292_ _10771_/A _10291_/X _19871_/Q vssd1 vssd1 vccd1 vccd1 _19871_/D sky130_fd_sc_hd__mux2_1
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12031_ _19344_/Q _12023_/X _12030_/X _12024_/X vssd1 vssd1 vccd1 vccd1 _19344_/D
+ sky130_fd_sc_hd__a22o_1
Xhold180 input31/X vssd1 vssd1 vccd1 vccd1 hold180/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold191 HADDR[6] vssd1 vssd1 vccd1 vccd1 input29/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_160_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17145__S _17529_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16770_ _16769_/X _11320_/Y _17493_/S vssd1 vssd1 vccd1 vccd1 _16770_/X sky130_fd_sc_hd__mux2_1
XFILLER_219_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13982_ _18692_/Q vssd1 vssd1 vccd1 vccd1 _14022_/A sky130_fd_sc_hd__inv_2
X_15721_ _15721_/A _15725_/B vssd1 vssd1 vccd1 vccd1 _18654_/D sky130_fd_sc_hd__nor2_1
XFILLER_234_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19057__RESET_B repeater257/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12933_ _19268_/Q vssd1 vssd1 vccd1 vccd1 _12933_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16233__A1 _15253_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18440_ _18795_/CLK _18440_/D vssd1 vssd1 vccd1 vccd1 _18440_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15652_ _15657_/B _15651_/X _15643_/X vssd1 vssd1 vccd1 vccd1 _15652_/X sky130_fd_sc_hd__o21a_1
XFILLER_222_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12864_ _12864_/A vssd1 vssd1 vccd1 vccd1 _13021_/B sky130_fd_sc_hd__clkbuf_2
XPHY_4151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14603_ _18281_/Q _14599_/X _14600_/X _14602_/X vssd1 vssd1 vccd1 vccd1 _18281_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_4173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18371_ _19647_/CLK _18371_/D vssd1 vssd1 vccd1 vccd1 _18371_/Q sky130_fd_sc_hd__dfxtp_1
X_11815_ _11822_/A vssd1 vssd1 vccd1 vccd1 _11815_/X sky130_fd_sc_hd__clkbuf_2
XPHY_4184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12795_ _12790_/Y _18809_/Q _19230_/Q _13531_/A _12794_/X vssd1 vssd1 vccd1 vccd1
+ _12808_/B sky130_fd_sc_hd__o221a_1
XANTENNA_output101_A _16077_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15583_ _18590_/Q vssd1 vssd1 vccd1 vccd1 _15583_/Y sky130_fd_sc_hd__inv_2
XPHY_4195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_215_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_230_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17322_ _17321_/X _09672_/Y _17523_/S vssd1 vssd1 vccd1 vccd1 _17322_/X sky130_fd_sc_hd__mux2_1
X_14534_ _18321_/Q _14530_/X _14531_/X _14533_/X vssd1 vssd1 vccd1 vccd1 _18321_/D
+ sky130_fd_sc_hd__a22o_1
X_11746_ hold139/X _10948_/X _19494_/Q _10951_/X vssd1 vssd1 vccd1 vccd1 hold141/A
+ sky130_fd_sc_hd__o22a_1
XPHY_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17253_ _17473_/A0 _16569_/Y _17512_/S vssd1 vssd1 vccd1 vccd1 _17253_/X sky130_fd_sc_hd__mux2_1
XPHY_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11677_ _10491_/B _11674_/X _10493_/B _11675_/X vssd1 vssd1 vccd1 vccd1 _19540_/D
+ sky130_fd_sc_hd__o22ai_1
XFILLER_169_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14465_ _14465_/A vssd1 vssd1 vccd1 vccd1 _14465_/X sky130_fd_sc_hd__clkbuf_2
XPHY_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18692__RESET_B hold359/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12318__A _12334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16204_ _16204_/A vssd1 vssd1 vccd1 vccd1 _16437_/A sky130_fd_sc_hd__clkbuf_2
X_10628_ _10558_/B _10618_/X _10579_/B _10608_/A vssd1 vssd1 vccd1 vccd1 _19805_/D
+ sky130_fd_sc_hd__o22ai_1
X_13416_ _13413_/Y _18850_/Q _20104_/Q _13428_/C _13415_/X vssd1 vssd1 vccd1 vccd1
+ _13417_/D sky130_fd_sc_hd__o221a_1
X_14396_ _14396_/A vssd1 vssd1 vccd1 vccd1 _14396_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_17184_ _17183_/X _13864_/Y _17545_/S vssd1 vssd1 vccd1 vccd1 _17184_/X sky130_fd_sc_hd__mux2_1
XFILLER_190_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13347_ _13431_/C _13442_/A vssd1 vssd1 vccd1 vccd1 _13348_/B sky130_fd_sc_hd__or2_2
X_16135_ _19773_/Q vssd1 vssd1 vccd1 vccd1 _16135_/Y sky130_fd_sc_hd__inv_2
XFILLER_143_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10559_ _19806_/Q _19805_/Q _10559_/C vssd1 vssd1 vccd1 vccd1 _10572_/B sky130_fd_sc_hd__or3_1
XFILLER_155_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_185_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13278_ _13278_/A _13278_/B _13278_/C _13299_/A vssd1 vssd1 vccd1 vccd1 _13278_/X
+ sky130_fd_sc_hd__or4b_1
X_16066_ _17462_/X vssd1 vssd1 vccd1 vccd1 _16066_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19898__RESET_B repeater195/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12229_ _12229_/A vssd1 vssd1 vccd1 vccd1 _12229_/X sky130_fd_sc_hd__clkbuf_2
X_15017_ _18045_/Q _15010_/X _15002_/X _15012_/X vssd1 vssd1 vccd1 vccd1 _18045_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19827__RESET_B repeater271/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19825_ _19825_/CLK _19825_/D repeater229/X vssd1 vssd1 vccd1 vccd1 _19825_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_110_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17895__S1 _18759_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11892__A _11892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15364__A _15364_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17055__S _17541_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19756_ _19772_/CLK _19756_/D repeater189/X vssd1 vssd1 vccd1 vccd1 _19756_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_110_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16968_ _16967_/X _19963_/Q _17488_/S vssd1 vssd1 vccd1 vccd1 _16968_/X sky130_fd_sc_hd__mux2_1
XFILLER_111_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_204_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18707_ _19224_/CLK _18707_/D repeater186/X vssd1 vssd1 vccd1 vccd1 _18707_/Q sky130_fd_sc_hd__dfrtp_1
X_15919_ _18139_/Q vssd1 vssd1 vccd1 vccd1 _15919_/Y sky130_fd_sc_hd__inv_2
XFILLER_209_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19687_ _19720_/CLK _19687_/D repeater202/X vssd1 vssd1 vccd1 vccd1 _19687_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__16894__S _17488_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16899_ _16898_/X _09875_/A _17513_/S vssd1 vssd1 vccd1 vccd1 _16899_/X sky130_fd_sc_hd__mux2_1
XFILLER_224_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_204_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17421__A0 _15768_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_209_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09440_ _09440_/A _09440_/B _09440_/C _09440_/D vssd1 vssd1 vccd1 vccd1 _09464_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_80_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18638_ _19810_/CLK _18638_/D repeater226/X vssd1 vssd1 vccd1 vccd1 _18638_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_65_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_224_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09371_ _20006_/Q vssd1 vssd1 vccd1 vccd1 _09467_/A sky130_fd_sc_hd__inv_2
X_18569_ _19846_/CLK _18569_/D repeater272/X vssd1 vssd1 vccd1 vccd1 _18569_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_220_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_240_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_220_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_177_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_178_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12228__A _12228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_192_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14710__B2 _14701_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_248_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_181_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17886__S1 _18759_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16463__B2 _16394_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09707_ _09794_/A _19411_/Q _09750_/A _19423_/Q _09706_/X vssd1 vssd1 vccd1 vccd1
+ _09713_/B sky130_fd_sc_hd__o221a_1
XFILLER_244_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17412__A0 _15963_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09638_ _19977_/Q vssd1 vssd1 vccd1 vccd1 _09789_/A sky130_fd_sc_hd__inv_2
XANTENNA__20055__RESET_B repeater204/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09569_ _09607_/A vssd1 vssd1 vccd1 vccd1 _09604_/B sky130_fd_sc_hd__clkbuf_4
XPHY_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11600_ _11600_/A vssd1 vssd1 vccd1 vccd1 _11600_/Y sky130_fd_sc_hd__inv_2
XPHY_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_212_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12580_ _19044_/Q _12576_/X _12406_/X _12577_/X vssd1 vssd1 vccd1 vccd1 _19044_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_184_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11531_ _11467_/A _11531_/A2 _11523_/X _11529_/Y vssd1 vssd1 vccd1 vccd1 _19586_/D
+ sky130_fd_sc_hd__a211oi_4
XPHY_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17810__S1 _18750_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14250_ _14251_/A vssd1 vssd1 vccd1 vccd1 _14250_/X sky130_fd_sc_hd__clkbuf_2
X_11462_ _11462_/A _11538_/A vssd1 vssd1 vccd1 vccd1 _11463_/B sky130_fd_sc_hd__or2_2
XPHY_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_52_HCLK clkbuf_opt_1_HCLK/A vssd1 vssd1 vccd1 vccd1 _19794_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13201_ _13069_/B _13200_/A _18896_/Q _13200_/Y _13162_/X vssd1 vssd1 vccd1 vccd1
+ _18896_/D sky130_fd_sc_hd__o221a_1
XANTENNA__11977__A _11977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10413_ _10147_/X _10408_/X _10413_/S vssd1 vssd1 vccd1 vccd1 _19847_/D sky130_fd_sc_hd__mux2_1
X_14181_ _19101_/Q vssd1 vssd1 vccd1 vccd1 _16467_/A sky130_fd_sc_hd__inv_2
XFILLER_152_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11393_ _19135_/Q vssd1 vssd1 vccd1 vccd1 _11393_/Y sky130_fd_sc_hd__inv_2
XANTENNA__10881__A hold237/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_180_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13132_ _19170_/Q vssd1 vssd1 vccd1 vccd1 _13132_/Y sky130_fd_sc_hd__inv_2
X_10344_ _19864_/Q _10344_/B vssd1 vssd1 vccd1 vccd1 _10344_/Y sky130_fd_sc_hd__nor2_1
XFILLER_152_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16979__S _17524_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19991__RESET_B repeater192/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18511__CLK _19780_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17940_ _19842_/CLK _17940_/D vssd1 vssd1 vccd1 vccd1 _17940_/Q sky130_fd_sc_hd__dfxtp_1
X_13063_ _13063_/A _13210_/A vssd1 vssd1 vccd1 vccd1 _13064_/B sky130_fd_sc_hd__or2_1
XANTENNA__09708__B2 _19423_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10275_ _10263_/X _10268_/B _11039_/B vssd1 vssd1 vccd1 vccd1 _10275_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__19920__RESET_B repeater230/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12712__B1 hold242/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12014_ _19354_/Q _12009_/X _09037_/X _12010_/X vssd1 vssd1 vccd1 vccd1 _19354_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_105_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09184__A2 _09164_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17871_ _16156_/Y _16157_/Y _16158_/Y _16159_/Y _17913_/S0 _19632_/Q vssd1 vssd1
+ vccd1 vccd1 _17871_/X sky130_fd_sc_hd__mux4_2
Xclkbuf_4_6_0_HCLK clkbuf_4_7_0_HCLK/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_6_0_HCLK/X
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_120_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17877__S1 _18759_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_238_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19610_ _19610_/CLK _19610_/D hold343/X vssd1 vssd1 vccd1 vccd1 _19610_/Q sky130_fd_sc_hd__dfrtp_2
X_16822_ _15963_/X _09552_/Y _17534_/S vssd1 vssd1 vccd1 vccd1 _16822_/X sky130_fd_sc_hd__mux2_1
XFILLER_120_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_238_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19541_ _19541_/CLK _19541_/D repeater221/X vssd1 vssd1 vccd1 vccd1 _19541_/Q sky130_fd_sc_hd__dfrtp_1
X_16753_ _10133_/B _08986_/Y _10133_/A _08986_/A vssd1 vssd1 vccd1 vccd1 _20124_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_47_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13965_ _13802_/B _13967_/A _13802_/A vssd1 vssd1 vccd1 vccd1 _13966_/B sky130_fd_sc_hd__o21a_1
XFILLER_171_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_206_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17603__S _17605_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11217__A _19013_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15704_ _18618_/Q _15697_/A _18619_/Q vssd1 vssd1 vccd1 vccd1 _15704_/X sky130_fd_sc_hd__o21a_1
X_19472_ _19513_/CLK hold204/X repeater260/X vssd1 vssd1 vccd1 vccd1 _19472_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_47_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12916_ _12916_/A _12916_/B _12916_/C _12915_/X vssd1 vssd1 vccd1 vccd1 _12916_/X
+ sky130_fd_sc_hd__or4b_1
XFILLER_206_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16684_ _16684_/A vssd1 vssd1 vccd1 vccd1 _16684_/X sky130_fd_sc_hd__clkbuf_2
X_13896_ _19220_/Q _13830_/B _13845_/Y _18714_/Q _13895_/X vssd1 vssd1 vccd1 vccd1
+ _13897_/D sky130_fd_sc_hd__o221a_1
XFILLER_207_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_234_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18423_ _19637_/CLK _18423_/D vssd1 vssd1 vccd1 vccd1 _18423_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_234_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15635_ _18603_/Q vssd1 vssd1 vccd1 vccd1 _15635_/Y sky130_fd_sc_hd__inv_2
X_12847_ _18937_/Q vssd1 vssd1 vccd1 vccd1 _12965_/B sky130_fd_sc_hd__inv_1
XFILLER_222_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18873__RESET_B repeater208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13432__A _19260_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18354_ _18412_/CLK _18354_/D vssd1 vssd1 vccd1 vccd1 _18354_/Q sky130_fd_sc_hd__dfxtp_1
X_15566_ _15566_/A vssd1 vssd1 vccd1 vccd1 _15566_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17706__A1 _19771_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_187_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12778_ _18810_/Q vssd1 vssd1 vccd1 vccd1 _13534_/A sky130_fd_sc_hd__inv_2
XPHY_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17305_ _15768_/Y _14160_/Y _17546_/S vssd1 vssd1 vccd1 vccd1 _17305_/X sky130_fd_sc_hd__mux2_1
X_14517_ _14517_/A _14545_/B _14571_/C vssd1 vssd1 vccd1 vccd1 _14519_/A sky130_fd_sc_hd__or3_4
XFILLER_230_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_202_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18285_ _18435_/CLK _18285_/D vssd1 vssd1 vccd1 vccd1 _18285_/Q sky130_fd_sc_hd__dfxtp_1
X_11729_ _19506_/Q _11723_/X _16938_/X _11724_/X vssd1 vssd1 vccd1 vccd1 hold228/A
+ sky130_fd_sc_hd__a22o_1
X_15497_ _18569_/Q vssd1 vssd1 vccd1 vccd1 _15497_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17801__S1 _18750_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17236_ _17235_/X _13077_/A _17542_/S vssd1 vssd1 vccd1 vccd1 _17236_/X sky130_fd_sc_hd__mux2_2
X_14448_ _18371_/Q _14438_/A _14403_/X _14439_/A vssd1 vssd1 vccd1 vccd1 _18371_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_156_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17167_ _16484_/X _10206_/Y _17566_/S vssd1 vssd1 vccd1 vccd1 _17167_/X sky130_fd_sc_hd__mux2_1
X_14379_ _14490_/A _14963_/B _15058_/C vssd1 vssd1 vccd1 vccd1 _14381_/A sky130_fd_sc_hd__or3_4
XFILLER_128_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_183_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16118_ _16204_/A _18740_/Q vssd1 vssd1 vccd1 vccd1 _16118_/X sky130_fd_sc_hd__and2_1
XANTENNA__18191__CLK _18198_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17098_ _17097_/X _09855_/A _17518_/S vssd1 vssd1 vccd1 vccd1 _17098_/X sky130_fd_sc_hd__mux2_1
XANTENNA__16889__S _17546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16049_ _16303_/A vssd1 vssd1 vccd1 vccd1 _16049_/X sky130_fd_sc_hd__clkbuf_2
X_08940_ _19854_/Q vssd1 vssd1 vccd1 vccd1 _10321_/C sky130_fd_sc_hd__inv_2
XANTENNA__19661__RESET_B repeater270/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12703__B1 _12536_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17868__S1 _18759_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19808_ _19808_/CLK _19808_/D repeater224/X vssd1 vssd1 vccd1 vccd1 _19808_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_57_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09092__A hold326/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19739_ _20050_/CLK _19739_/D repeater206/X vssd1 vssd1 vccd1 vccd1 _19739_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_225_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17513__S _17513_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16748__A2 _18757_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_241_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09423_ _19917_/Q vssd1 vssd1 vccd1 vccd1 _10015_/C sky130_fd_sc_hd__inv_2
XFILLER_198_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09354_ _20023_/Q vssd1 vssd1 vccd1 vccd1 _09483_/A sky130_fd_sc_hd__inv_2
XANTENNA__18543__RESET_B repeater221/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_178_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09285_ _09293_/A vssd1 vssd1 vccd1 vccd1 _09285_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_leaf_134_HCLK_A clkbuf_4_6_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_220_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_193_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__19749__RESET_B repeater204/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14173__A _19111_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11745__B2 _11731_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16799__S _17541_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_192_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14144__C1 _14106_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10060_ _10047_/A _10059_/A _19931_/Q _10059_/Y _10053_/X vssd1 vssd1 vccd1 vccd1
+ _19931_/D sky130_fd_sc_hd__o221a_1
XANTENNA__19331__RESET_B hold371/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_248_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17859__S1 _18761_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14447__B1 _14419_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17423__S _17545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10962_ _10962_/A _10992_/A vssd1 vssd1 vccd1 vccd1 _10987_/A sky130_fd_sc_hd__or2_1
X_13750_ _13750_/A vssd1 vssd1 vccd1 vccd1 _13751_/A sky130_fd_sc_hd__inv_2
XFILLER_244_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13670__A1 _18778_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16739__A2 _16493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__20017__CLK _20091_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16547__B _16583_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_204_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12701_ _18965_/Q _12698_/X _12602_/X _12699_/X vssd1 vssd1 vccd1 vccd1 _18965_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_244_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_216_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10893_ _10894_/A vssd1 vssd1 vccd1 vccd1 _10893_/X sky130_fd_sc_hd__clkbuf_2
X_13681_ _18773_/Q _13671_/X _13680_/X _13672_/X vssd1 vssd1 vccd1 vccd1 _18773_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10876__A hold248/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_14_0_HCLK clkbuf_3_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_3_HCLK/A
+ sky130_fd_sc_hd__clkbuf_1
X_15420_ _19611_/Q vssd1 vssd1 vccd1 vccd1 _15420_/Y sky130_fd_sc_hd__inv_2
XPHY_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12632_ _19012_/Q _12629_/X _12404_/X _12630_/X vssd1 vssd1 vccd1 vccd1 _19012_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15351_ _18497_/Q _14227_/B _14228_/B vssd1 vssd1 vccd1 vccd1 _15351_/X sky130_fd_sc_hd__a21bo_1
X_12563_ _12577_/A vssd1 vssd1 vccd1 vccd1 _12563_/X sky130_fd_sc_hd__buf_1
XPHY_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16563__A _16638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17795__S0 _17923_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11514_ _11514_/A vssd1 vssd1 vccd1 vccd1 _11514_/Y sky130_fd_sc_hd__inv_2
X_14302_ _14517_/A _14450_/B _14557_/C vssd1 vssd1 vccd1 vccd1 _14304_/A sky130_fd_sc_hd__or3_4
XFILLER_157_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18070_ _18169_/CLK _18070_/D vssd1 vssd1 vccd1 vccd1 _18070_/Q sky130_fd_sc_hd__dfxtp_1
X_15282_ _15282_/A vssd1 vssd1 vccd1 vccd1 _18555_/D sky130_fd_sc_hd__inv_2
XFILLER_200_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12494_ _19091_/Q _12489_/X _12380_/X _12492_/X vssd1 vssd1 vccd1 vccd1 _19091_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17021_ _17020_/X _09490_/A _17482_/S vssd1 vssd1 vccd1 vccd1 _17021_/X sky130_fd_sc_hd__mux2_1
X_14233_ _18503_/Q _14233_/B vssd1 vssd1 vccd1 vccd1 _14236_/A sky130_fd_sc_hd__or2_4
X_11445_ _19155_/Q vssd1 vssd1 vccd1 vccd1 _11445_/Y sky130_fd_sc_hd__inv_2
XFILLER_172_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_56_HCLK_A clkbuf_4_9_0_HCLK/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14164_ _16644_/A _18694_/Q _19115_/Q _14024_/A vssd1 vssd1 vccd1 vccd1 _14164_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_109_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11376_ _11639_/C _19127_/Q _11582_/A _19149_/Q vssd1 vssd1 vccd1 vccd1 _11376_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__19419__RESET_B repeater192/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_180_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16675__A1 _17070_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10327_ _10327_/A _10357_/A vssd1 vssd1 vccd1 vccd1 _10352_/A sky130_fd_sc_hd__or2_1
X_13115_ _19184_/Q vssd1 vssd1 vccd1 vccd1 _13115_/Y sky130_fd_sc_hd__inv_2
X_18972_ _19595_/CLK _18972_/D repeater282/X vssd1 vssd1 vccd1 vccd1 _18972_/Q sky130_fd_sc_hd__dfrtp_4
X_14095_ _14116_/A vssd1 vssd1 vccd1 vccd1 _14112_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_98_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14686__B1 _14604_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17923_ _18297_/Q _18289_/Q _18281_/Q _18449_/Q _17923_/S0 _19646_/Q vssd1 vssd1
+ vccd1 vccd1 _17923_/X sky130_fd_sc_hd__mux4_2
X_13046_ _18900_/Q vssd1 vssd1 vccd1 vccd1 _13072_/A sky130_fd_sc_hd__inv_2
XFILLER_124_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10258_ _15296_/A _11027_/B vssd1 vssd1 vccd1 vccd1 _11029_/A sky130_fd_sc_hd__nand2_2
X_17854_ _17850_/X _17851_/X _17852_/X _17853_/X _19633_/Q _19634_/Q vssd1 vssd1 vccd1
+ vccd1 _17854_/X sky130_fd_sc_hd__mux4_2
XFILLER_67_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10189_ _19330_/Q vssd1 vssd1 vccd1 vccd1 _11869_/A sky130_fd_sc_hd__inv_2
XANTENNA__10172__B1 _09086_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16805_ _16804_/X _12902_/Y _17487_/S vssd1 vssd1 vccd1 vccd1 _16805_/X sky130_fd_sc_hd__mux2_1
XFILLER_208_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17785_ _18318_/Q _18438_/Q _18430_/Q _18422_/Q _17923_/S0 _19646_/Q vssd1 vssd1
+ vccd1 vccd1 _17785_/X sky130_fd_sc_hd__mux4_1
XFILLER_19_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14997_ _18056_/Q _14991_/X _14996_/X _14994_/X vssd1 vssd1 vccd1 vccd1 _18056_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_47_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19524_ _19771_/CLK _19524_/D repeater190/X vssd1 vssd1 vccd1 vccd1 _19524_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__17333__S _17546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16736_ _19092_/Q vssd1 vssd1 vccd1 vccd1 _16736_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_207_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_0_HCLK clkbuf_0_HCLK/X vssd1 vssd1 vccd1 vccd1 clkbuf_1_1_1_HCLK/A sky130_fd_sc_hd__clkbuf_1
XFILLER_47_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13948_ _13948_/A _13957_/A vssd1 vssd1 vccd1 vccd1 _13949_/B sky130_fd_sc_hd__or2_2
XFILLER_223_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_98_HCLK clkbuf_4_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19208_/CLK sky130_fd_sc_hd__clkbuf_16
X_19455_ _19462_/CLK _19455_/D repeater272/X vssd1 vssd1 vccd1 vccd1 _19455_/Q sky130_fd_sc_hd__dfrtp_1
X_16667_ _16667_/A _16668_/B vssd1 vssd1 vccd1 vccd1 _16667_/Y sky130_fd_sc_hd__nor2_1
X_13879_ _19205_/Q vssd1 vssd1 vccd1 vccd1 _13879_/Y sky130_fd_sc_hd__inv_2
XANTENNA__14258__A _14259_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18406_ _18473_/CLK _18406_/D vssd1 vssd1 vccd1 vccd1 _18406_/Q sky130_fd_sc_hd__dfxtp_1
X_15618_ _15618_/A _15618_/B vssd1 vssd1 vccd1 vccd1 _15618_/Y sky130_fd_sc_hd__nor2_1
X_19386_ _19933_/CLK _19386_/D repeater235/X vssd1 vssd1 vccd1 vccd1 _19386_/Q sky130_fd_sc_hd__dfrtp_2
X_16598_ _16598_/A vssd1 vssd1 vccd1 vccd1 _16598_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__14610__B1 _14582_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18557__CLK _19992_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18337_ _19849_/CLK _18337_/D vssd1 vssd1 vccd1 vccd1 _18337_/Q sky130_fd_sc_hd__dfxtp_1
X_15549_ _18581_/Q vssd1 vssd1 vccd1 vccd1 _15552_/A sky130_fd_sc_hd__inv_2
XFILLER_175_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_202_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17786__S0 _17923_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_175_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09070_ hold240/X vssd1 vssd1 vccd1 vccd1 hold239/A sky130_fd_sc_hd__buf_4
X_18268_ _18268_/CLK _18268_/D vssd1 vssd1 vccd1 vccd1 _18268_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_4_HCLK clkbuf_4_0_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19849_/CLK sky130_fd_sc_hd__clkbuf_16
X_17219_ _15963_/X _12816_/Y _17534_/S vssd1 vssd1 vccd1 vccd1 _17219_/X sky130_fd_sc_hd__mux2_1
XFILLER_116_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19842__RESET_B repeater270/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18199_ _18216_/CLK _18199_/D vssd1 vssd1 vccd1 vccd1 _18199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17508__S _17568_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10026__A _10026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09972_ _09972_/A vssd1 vssd1 vccd1 vccd1 _09972_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08923_ _19863_/Q vssd1 vssd1 vccd1 vccd1 _10329_/A sky130_fd_sc_hd__inv_2
X_20092_ _20120_/CLK _20092_/D repeater234/X vssd1 vssd1 vccd1 vccd1 _20092_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__12241__A _14405_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_242_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10163__B1 _09105_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17091__A1 _12913_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18795__RESET_B repeater261/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17243__S _17545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_226_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18724__RESET_B repeater253/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_241_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_226_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_241_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09406_ _19915_/Q vssd1 vssd1 vccd1 vccd1 _10087_/A sky130_fd_sc_hd__inv_2
XFILLER_198_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_201_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_187_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09337_ _20039_/Q _13766_/D _10786_/B vssd1 vssd1 vccd1 vccd1 _20039_/D sky130_fd_sc_hd__a21o_1
XFILLER_139_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11966__A1 _19380_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17777__S0 _17923_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09268_ _09340_/B _12436_/C vssd1 vssd1 vccd1 vccd1 _09270_/A sky130_fd_sc_hd__or2_4
XFILLER_138_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_194_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_hold307_A HWDATA[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_194_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_193_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09199_ _09199_/A vssd1 vssd1 vccd1 vccd1 _13283_/B sky130_fd_sc_hd__inv_2
XANTENNA__11718__A1 _19515_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11230_ _19007_/Q vssd1 vssd1 vccd1 vccd1 _11230_/Y sky130_fd_sc_hd__inv_2
XFILLER_146_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11161_ _19616_/Q _11161_/B vssd1 vssd1 vccd1 vccd1 _11162_/B sky130_fd_sc_hd__or2_1
XANTENNA__17418__S _17543_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10112_ _18558_/Q _15453_/A _18559_/Q vssd1 vssd1 vccd1 vccd1 _15457_/A sky130_fd_sc_hd__or3_1
X_11092_ _11059_/Y _11076_/X _11070_/Y _11091_/X vssd1 vssd1 vccd1 vccd1 _19640_/D
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_248_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10043_ _10043_/A _10065_/A vssd1 vssd1 vccd1 vccd1 _10044_/B sky130_fd_sc_hd__or2_2
X_14920_ _14922_/A vssd1 vssd1 vccd1 vccd1 _14920_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_49_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20070__RESET_B repeater207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14851_ _18142_/Q _14845_/X _14810_/X _14847_/X vssd1 vssd1 vccd1 vccd1 _18142_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_input25_A HADDR[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11075__A1_N _19632_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15093__B1 _09255_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17153__S _17541_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13802_ _13802_/A _13802_/B _13964_/C vssd1 vssd1 vccd1 vccd1 _13944_/C sky130_fd_sc_hd__or3_1
X_17570_ _19822_/Q _19773_/Q _18519_/Q vssd1 vssd1 vccd1 vccd1 _17570_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14782_ hold321/X vssd1 vssd1 vccd1 vccd1 _14782_/X sky130_fd_sc_hd__buf_2
XFILLER_205_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11994_ _15774_/A _11998_/A vssd1 vssd1 vccd1 vccd1 _11995_/S sky130_fd_sc_hd__or2_1
XFILLER_72_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16521_ _17292_/X _16508_/X _17279_/X _16235_/X _16520_/X vssd1 vssd1 vccd1 vccd1
+ _16521_/X sky130_fd_sc_hd__o221a_1
X_13733_ _13733_/A _14286_/B vssd1 vssd1 vccd1 vccd1 _13733_/Y sky130_fd_sc_hd__nor2_1
X_10945_ _19670_/Q _10618_/X _10601_/X vssd1 vssd1 vccd1 vccd1 _19670_/D sky130_fd_sc_hd__o21a_1
XANTENNA__16992__S _17488_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_216_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_231_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19240_ _19314_/CLK _19240_/D repeater239/X vssd1 vssd1 vccd1 vccd1 _19240_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_188_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16452_ _19772_/Q vssd1 vssd1 vccd1 vccd1 _16452_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_231_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13664_ _13671_/A vssd1 vssd1 vccd1 vccd1 _13664_/X sky130_fd_sc_hd__clkbuf_2
X_10876_ hold248/X vssd1 vssd1 vccd1 vccd1 _14273_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_188_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15403_ _18534_/Q _13221_/B _13222_/B vssd1 vssd1 vccd1 vccd1 _15403_/X sky130_fd_sc_hd__a21bo_1
XPHY_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12615_ _12651_/A vssd1 vssd1 vccd1 vccd1 _12630_/A sky130_fd_sc_hd__clkbuf_2
X_19171_ _19208_/CLK _19171_/D hold370/X vssd1 vssd1 vccd1 vccd1 _19171_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16383_ _16381_/Y _16303_/X _16382_/Y _15850_/B vssd1 vssd1 vccd1 vccd1 _16383_/X
+ sky130_fd_sc_hd__o22a_1
XPHY_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13595_ _18815_/Q _13597_/B _13591_/X _13595_/C1 vssd1 vssd1 vccd1 vccd1 _18815_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17768__S0 _17923_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18122_ _18260_/CLK _18122_/D vssd1 vssd1 vccd1 vccd1 _18122_/Q sky130_fd_sc_hd__dfxtp_1
X_15334_ _15334_/A _15334_/B _15334_/C vssd1 vssd1 vccd1 vccd1 _18481_/D sky130_fd_sc_hd__nor3_1
XPHY_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_185_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_200_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12546_ hold242/X _12556_/A _17614_/S _12249_/A _12545_/Y vssd1 vssd1 vccd1 vccd1
+ _12551_/C sky130_fd_sc_hd__a221o_1
XFILLER_118_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19975__CLK _19984_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18053_ _18142_/CLK _18053_/D vssd1 vssd1 vccd1 vccd1 _18053_/Q sky130_fd_sc_hd__dfxtp_1
X_15265_ _15259_/A _15242_/Y _15263_/Y _15250_/Y _15264_/X vssd1 vssd1 vccd1 vccd1
+ _15266_/B sky130_fd_sc_hd__o32a_1
XFILLER_177_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12477_ _19100_/Q _12471_/X _12296_/X _12472_/X vssd1 vssd1 vccd1 vccd1 _19100_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12906__B1 _12905_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17004_ _17003_/X _15657_/A _17318_/S vssd1 vssd1 vccd1 vccd1 _17004_/X sky130_fd_sc_hd__mux2_1
XFILLER_126_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14216_ _19117_/Q _14026_/A _19094_/Q _14004_/A vssd1 vssd1 vccd1 vccd1 _14216_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA_output93_A _16656_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11428_ _19151_/Q vssd1 vssd1 vccd1 vccd1 _11428_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15196_ _15196_/A vssd1 vssd1 vccd1 vccd1 _17564_/S sky130_fd_sc_hd__clkinv_8
XANTENNA__17328__S _17535_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11359_ _19609_/Q _11358_/Y _19602_/Q _11301_/Y vssd1 vssd1 vccd1 vccd1 _11359_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_4_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14147_ _14005_/A _14147_/A2 _14145_/Y _14106_/X vssd1 vssd1 vccd1 vccd1 _18674_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_193_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14659__B1 _14600_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14078_ _14077_/Y _18687_/Q _19076_/Q _14017_/A vssd1 vssd1 vccd1 vccd1 _14078_/X
+ sky130_fd_sc_hd__o22a_1
X_18955_ _18959_/CLK _18955_/D repeater257/X vssd1 vssd1 vccd1 vccd1 _18955_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_140_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17906_ _15806_/Y _15807_/Y _15808_/Y _15809_/Y _17908_/S0 _18759_/Q vssd1 vssd1
+ vccd1 vccd1 _17906_/X sky130_fd_sc_hd__mux4_2
X_13029_ _18917_/Q vssd1 vssd1 vccd1 vccd1 _13089_/A sky130_fd_sc_hd__inv_2
X_18886_ _18886_/CLK _18886_/D repeater220/X vssd1 vssd1 vccd1 vccd1 _18886_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_121_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17073__A1 _20111_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_227_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10696__A1 _10448_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17837_ _16425_/Y _16426_/Y _16427_/Y _16428_/Y _17908_/S0 _18759_/Q vssd1 vssd1
+ vccd1 vccd1 _17837_/X sky130_fd_sc_hd__mux4_1
XANTENNA__11893__B1 hold314/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17063__S _17548_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xrebuffer16 _13071_/B vssd1 vssd1 vccd1 vccd1 _13197_/C1 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer27 _13061_/B vssd1 vssd1 vccd1 vccd1 _13213_/A sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_208_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17768_ _18290_/Q _18282_/Q _18274_/Q _18442_/Q _17923_/S0 _19646_/Q vssd1 vssd1
+ vccd1 vccd1 _17768_/X sky130_fd_sc_hd__mux4_2
Xrebuffer38 _19418_/Q vssd1 vssd1 vccd1 vccd1 _09722_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_47_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xrebuffer49 _18730_/Q vssd1 vssd1 vccd1 vccd1 _13782_/A sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_212_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_207_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_223_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_208_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16719_ _16719_/A _16721_/B vssd1 vssd1 vccd1 vccd1 _16719_/Y sky130_fd_sc_hd__nor2_1
X_19507_ _19510_/CLK hold218/X repeater256/X vssd1 vssd1 vccd1 vccd1 _19507_/Q sky130_fd_sc_hd__dfrtp_1
X_17699_ _19819_/Q _19761_/Q _18548_/Q vssd1 vssd1 vccd1 vccd1 _17699_/X sky130_fd_sc_hd__mux2_1
XFILLER_212_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_223_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19438_ _19905_/CLK _19438_/D repeater210/X vssd1 vssd1 vccd1 vccd1 _19438_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_50_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_211_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_195_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19369_ _19971_/CLK _19369_/D repeater241/X vssd1 vssd1 vccd1 vccd1 _19369_/Q sky130_fd_sc_hd__dfrtp_4
X_09122_ _20082_/Q vssd1 vssd1 vccd1 vccd1 _09149_/A sky130_fd_sc_hd__inv_2
Xrebuffer106 _13536_/B vssd1 vssd1 vccd1 vccd1 _13600_/A2 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer117 _13532_/B vssd1 vssd1 vccd1 vccd1 _13606_/A2 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_176_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_175_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09053_ _09084_/A vssd1 vssd1 vccd1 vccd1 _09053_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_176_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12236__A _13678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_191_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_105_HCLK clkbuf_4_7_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19224_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_144_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16650__B _16673_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16639__A1 _16912_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13570__B1 _13560_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17238__S _17546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09955_ _19968_/Q _09954_/Y _09950_/X _09877_/B vssd1 vssd1 vccd1 vccd1 _19968_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_131_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20075_ _20076_/CLK _20075_/D repeater196/X vssd1 vssd1 vccd1 vccd1 _20075_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09886_ _19957_/Q _09883_/Y _09870_/A _19354_/Q _09885_/X vssd1 vssd1 vccd1 vccd1
+ _09895_/B sky130_fd_sc_hd__o221a_1
XFILLER_106_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18905__RESET_B repeater188/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17064__A1 _19421_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_245_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15075__B1 hold236/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_245_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_213_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10730_ _19765_/Q _10721_/A _10427_/X _10722_/A vssd1 vssd1 vccd1 vccd1 _19765_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_241_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_213_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_213_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13389__B1 _20113_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_241_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10661_ _10676_/A vssd1 vssd1 vccd1 vccd1 _10661_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_185_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12400_ _12400_/A vssd1 vssd1 vccd1 vccd1 _12400_/X sky130_fd_sc_hd__buf_1
X_13380_ _20110_/Q vssd1 vssd1 vccd1 vccd1 _13380_/Y sky130_fd_sc_hd__clkinv_1
XFILLER_167_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10592_ _19804_/Q _10592_/B _19803_/Q vssd1 vssd1 vccd1 vccd1 _10594_/B sky130_fd_sc_hd__nor3b_4
XANTENNA__16327__B1 _15859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_222_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_194_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12331_ _19182_/Q _12327_/X _12088_/X _12328_/X vssd1 vssd1 vccd1 vccd1 _19182_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_31_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15050_ _18025_/Q _15047_/X _14992_/X _15049_/X vssd1 vssd1 vccd1 vccd1 _18025_/D
+ sky130_fd_sc_hd__a22o_1
X_12262_ _12300_/A vssd1 vssd1 vccd1 vccd1 _12277_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_107_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_181_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11213_ _19597_/Q vssd1 vssd1 vccd1 vccd1 _11477_/A sky130_fd_sc_hd__inv_2
X_14001_ _18673_/Q vssd1 vssd1 vccd1 vccd1 _14004_/A sky130_fd_sc_hd__inv_2
XANTENNA__17148__S _17517_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12193_ _19258_/Q _12189_/X _12069_/X _12192_/X vssd1 vssd1 vccd1 vccd1 _19258_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_135_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17922__S0 _17923_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11144_ _11144_/A _11144_/B vssd1 vssd1 vccd1 vccd1 _11144_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__16987__S _17546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput85 _16568_/Y vssd1 vssd1 vccd1 vccd1 HRDATA[15] sky130_fd_sc_hd__clkbuf_2
XFILLER_163_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput96 _16691_/Y vssd1 vssd1 vccd1 vccd1 HRDATA[25] sky130_fd_sc_hd__clkbuf_2
X_18740_ _20066_/CLK _18740_/D repeater209/X vssd1 vssd1 vccd1 vccd1 _18740_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11075_ _19632_/Q _11074_/Y _19632_/Q _11074_/Y vssd1 vssd1 vccd1 vccd1 _11103_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_15952_ _17954_/Q vssd1 vssd1 vccd1 vccd1 _15952_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_237_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_209_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10026_ _10026_/A vssd1 vssd1 vccd1 vccd1 _10026_/X sky130_fd_sc_hd__clkbuf_2
X_14903_ _18109_/Q _14896_/X _14709_/X _14898_/X vssd1 vssd1 vccd1 vccd1 _18109_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_37_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18671_ _18686_/CLK _18671_/D repeater252/X vssd1 vssd1 vccd1 vccd1 _18671_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA_output131_A _18642_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15883_ _15883_/A vssd1 vssd1 vccd1 vccd1 _15884_/A sky130_fd_sc_hd__buf_1
XFILLER_237_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17622_ _20040_/Q _15728_/Y _17622_/S vssd1 vssd1 vccd1 vccd1 _17622_/X sky130_fd_sc_hd__mux2_1
X_14834_ _14834_/A vssd1 vssd1 vccd1 vccd1 _14834_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__13705__A _18760_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14813__B1 _14812_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17553_ _17552_/X _20036_/Q _19497_/Q vssd1 vssd1 vccd1 vccd1 _17553_/X sky130_fd_sc_hd__mux2_1
X_14765_ _18190_/Q _14759_/X _14723_/X _14761_/X vssd1 vssd1 vccd1 vccd1 _18190_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_189_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11977_ _11977_/A vssd1 vssd1 vccd1 vccd1 _11977_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_205_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17611__S _17614_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16504_ _16504_/A vssd1 vssd1 vccd1 vccd1 _16504_/X sky130_fd_sc_hd__buf_4
X_13716_ _14641_/B _13704_/B _14628_/B _18758_/Q _13715_/Y vssd1 vssd1 vccd1 vccd1
+ _13721_/B sky130_fd_sc_hd__a221o_1
X_17484_ _17483_/X _13398_/Y _17535_/S vssd1 vssd1 vccd1 vccd1 _17484_/X sky130_fd_sc_hd__mux2_1
X_10928_ _17724_/X _10923_/X _19677_/Q _10924_/X vssd1 vssd1 vccd1 vccd1 _19677_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16566__B1 _17158_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14696_ _15195_/B _14696_/B vssd1 vssd1 vccd1 vccd1 _15121_/C sky130_fd_sc_hd__or2_2
XANTENNA__16735__B _16735_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19223_ _19293_/CLK _19223_/D repeater186/X vssd1 vssd1 vccd1 vccd1 _19223_/Q sky130_fd_sc_hd__dfrtp_1
X_16435_ _17312_/X _16435_/B vssd1 vssd1 vccd1 vccd1 _16435_/Y sky130_fd_sc_hd__nand2_1
X_13647_ _16957_/X _13644_/X _18794_/Q _13646_/X vssd1 vssd1 vccd1 vccd1 _18794_/D
+ sky130_fd_sc_hd__o22a_1
X_10859_ _19707_/Q _10855_/X _10448_/X _10857_/X vssd1 vssd1 vccd1 vccd1 _19707_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_158_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19154_ _19157_/CLK _19154_/D repeater268/X vssd1 vssd1 vccd1 vccd1 _19154_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16366_ _20065_/Q _16436_/B vssd1 vssd1 vccd1 vccd1 _16366_/Y sky130_fd_sc_hd__nand2_1
X_13578_ _18825_/Q _13577_/Y _13574_/X _13578_/C1 vssd1 vssd1 vccd1 vccd1 _18825_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_157_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_128_HCLK clkbuf_4_4_0_HCLK/X vssd1 vssd1 vccd1 vccd1 _19437_/CLK sky130_fd_sc_hd__clkbuf_16
X_18105_ _20077_/CLK _18105_/D vssd1 vssd1 vccd1 vccd1 _18105_/Q sky130_fd_sc_hd__dfxtp_1
X_15317_ _15439_/A _15261_/X _15316_/X vssd1 vssd1 vccd1 vccd1 _18626_/D sky130_fd_sc_hd__a21bo_1
XFILLER_158_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19085_ _19119_/CLK _19085_/D hold355/X vssd1 vssd1 vccd1 vccd1 _19085_/Q sky130_fd_sc_hd__dfrtp_4
X_12529_ _12529_/A vssd1 vssd1 vccd1 vccd1 _12529_/X sky130_fd_sc_hd__clkbuf_2
X_16297_ _20064_/Q _16436_/B vssd1 vssd1 vccd1 vccd1 _16297_/Y sky130_fd_sc_hd__nand2_1
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18036_ _19851_/CLK _18036_/D vssd1 vssd1 vccd1 vccd1 _18036_/Q sky130_fd_sc_hd__dfxtp_1
X_15248_ _19778_/Q _19777_/Q vssd1 vssd1 vccd1 vccd1 _18517_/D sky130_fd_sc_hd__or2_1
XFILLER_126_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12355__A1 _19169_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17058__S _17318_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15179_ _17938_/Q _15171_/A _09339_/X _15172_/A vssd1 vssd1 vccd1 vccd1 _17938_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_141_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17913__S0 _17913_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16897__S _17522_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19987_ _19992_/CLK _19987_/D repeater193/X vssd1 vssd1 vccd1 vccd1 _19987_/Q sky130_fd_sc_hd__dfrtp_1
X_09740_ _09740_/A _09740_/B vssd1 vssd1 vccd1 vccd1 _09784_/A sky130_fd_sc_hd__or2_1
X_18938_ _19325_/CLK _18938_/D repeater213/X vssd1 vssd1 vccd1 vccd1 _18938_/Q sky130_fd_sc_hd__dfrtp_2
.ends

