VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO DFFRAM_4K
  CLASS BLOCK ;
  FOREIGN DFFRAM_4K ;
  ORIGIN 0.000 0.000 ;
  SIZE 1100.000 BY 1400.000 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.290 1396.000 446.570 1400.000 ;
    END
  END A[0]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.090 1396.000 460.370 1400.000 ;
    END
  END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.890 1396.000 474.170 1400.000 ;
    END
  END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.690 1396.000 487.970 1400.000 ;
    END
  END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.030 1396.000 501.310 1400.000 ;
    END
  END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.830 1396.000 515.110 1400.000 ;
    END
  END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.630 1396.000 528.910 1400.000 ;
    END
  END A[6]
  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.430 1396.000 542.710 1400.000 ;
    END
  END A[7]
  PIN A[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.230 1396.000 556.510 1400.000 ;
    END
  END A[8]
  PIN A[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.030 1396.000 570.310 1400.000 ;
    END
  END A[9]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 583.830 1396.000 584.110 1400.000 ;
    END
  END CLK
  PIN Di[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.170 1396.000 666.450 1400.000 ;
    END
  END Di[0]
  PIN Di[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 803.710 1396.000 803.990 1400.000 ;
    END
  END Di[10]
  PIN Di[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.510 1396.000 817.790 1400.000 ;
    END
  END Di[11]
  PIN Di[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 831.310 1396.000 831.590 1400.000 ;
    END
  END Di[12]
  PIN Di[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 845.110 1396.000 845.390 1400.000 ;
    END
  END Di[13]
  PIN Di[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 858.910 1396.000 859.190 1400.000 ;
    END
  END Di[14]
  PIN Di[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 872.250 1396.000 872.530 1400.000 ;
    END
  END Di[15]
  PIN Di[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 886.050 1396.000 886.330 1400.000 ;
    END
  END Di[16]
  PIN Di[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 899.850 1396.000 900.130 1400.000 ;
    END
  END Di[17]
  PIN Di[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 913.650 1396.000 913.930 1400.000 ;
    END
  END Di[18]
  PIN Di[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.450 1396.000 927.730 1400.000 ;
    END
  END Di[19]
  PIN Di[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.970 1396.000 680.250 1400.000 ;
    END
  END Di[1]
  PIN Di[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 941.250 1396.000 941.530 1400.000 ;
    END
  END Di[20]
  PIN Di[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 955.050 1396.000 955.330 1400.000 ;
    END
  END Di[21]
  PIN Di[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 968.850 1396.000 969.130 1400.000 ;
    END
  END Di[22]
  PIN Di[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 982.650 1396.000 982.930 1400.000 ;
    END
  END Di[23]
  PIN Di[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.990 1396.000 996.270 1400.000 ;
    END
  END Di[24]
  PIN Di[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1009.790 1396.000 1010.070 1400.000 ;
    END
  END Di[25]
  PIN Di[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1023.590 1396.000 1023.870 1400.000 ;
    END
  END Di[26]
  PIN Di[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1037.390 1396.000 1037.670 1400.000 ;
    END
  END Di[27]
  PIN Di[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1051.190 1396.000 1051.470 1400.000 ;
    END
  END Di[28]
  PIN Di[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1064.990 1396.000 1065.270 1400.000 ;
    END
  END Di[29]
  PIN Di[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 693.770 1396.000 694.050 1400.000 ;
    END
  END Di[2]
  PIN Di[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1078.790 1396.000 1079.070 1400.000 ;
    END
  END Di[30]
  PIN Di[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1092.590 1396.000 1092.870 1400.000 ;
    END
  END Di[31]
  PIN Di[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.570 1396.000 707.850 1400.000 ;
    END
  END Di[3]
  PIN Di[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.370 1396.000 721.650 1400.000 ;
    END
  END Di[4]
  PIN Di[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.170 1396.000 735.450 1400.000 ;
    END
  END Di[5]
  PIN Di[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.510 1396.000 748.790 1400.000 ;
    END
  END Di[6]
  PIN Di[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 762.310 1396.000 762.590 1400.000 ;
    END
  END Di[7]
  PIN Di[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.110 1396.000 776.390 1400.000 ;
    END
  END Di[8]
  PIN Di[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.910 1396.000 790.190 1400.000 ;
    END
  END Di[9]
  PIN Do[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 1396.000 6.810 1400.000 ;
    END
  END Do[0]
  PIN Do[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 1396.000 143.890 1400.000 ;
    END
  END Do[10]
  PIN Do[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.410 1396.000 157.690 1400.000 ;
    END
  END Do[11]
  PIN Do[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.210 1396.000 171.490 1400.000 ;
    END
  END Do[12]
  PIN Do[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 1396.000 185.290 1400.000 ;
    END
  END Do[13]
  PIN Do[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.810 1396.000 199.090 1400.000 ;
    END
  END Do[14]
  PIN Do[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 1396.000 212.890 1400.000 ;
    END
  END Do[15]
  PIN Do[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 1396.000 226.690 1400.000 ;
    END
  END Do[16]
  PIN Do[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.210 1396.000 240.490 1400.000 ;
    END
  END Do[17]
  PIN Do[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.550 1396.000 253.830 1400.000 ;
    END
  END Do[18]
  PIN Do[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 1396.000 267.630 1400.000 ;
    END
  END Do[19]
  PIN Do[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 1396.000 20.150 1400.000 ;
    END
  END Do[1]
  PIN Do[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.150 1396.000 281.430 1400.000 ;
    END
  END Do[20]
  PIN Do[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.950 1396.000 295.230 1400.000 ;
    END
  END Do[21]
  PIN Do[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.750 1396.000 309.030 1400.000 ;
    END
  END Do[22]
  PIN Do[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.550 1396.000 322.830 1400.000 ;
    END
  END Do[23]
  PIN Do[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.350 1396.000 336.630 1400.000 ;
    END
  END Do[24]
  PIN Do[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.150 1396.000 350.430 1400.000 ;
    END
  END Do[25]
  PIN Do[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 1396.000 364.230 1400.000 ;
    END
  END Do[26]
  PIN Do[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.290 1396.000 377.570 1400.000 ;
    END
  END Do[27]
  PIN Do[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.090 1396.000 391.370 1400.000 ;
    END
  END Do[28]
  PIN Do[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.890 1396.000 405.170 1400.000 ;
    END
  END Do[29]
  PIN Do[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 1396.000 33.950 1400.000 ;
    END
  END Do[2]
  PIN Do[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 1396.000 418.970 1400.000 ;
    END
  END Do[30]
  PIN Do[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.490 1396.000 432.770 1400.000 ;
    END
  END Do[31]
  PIN Do[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 1396.000 47.750 1400.000 ;
    END
  END Do[3]
  PIN Do[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 1396.000 61.550 1400.000 ;
    END
  END Do[4]
  PIN Do[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 1396.000 75.350 1400.000 ;
    END
  END Do[5]
  PIN Do[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 1396.000 89.150 1400.000 ;
    END
  END Do[6]
  PIN Do[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.670 1396.000 102.950 1400.000 ;
    END
  END Do[7]
  PIN Do[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.470 1396.000 116.750 1400.000 ;
    END
  END Do[8]
  PIN Do[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 1396.000 130.090 1400.000 ;
    END
  END Do[9]
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.370 1396.000 652.650 1400.000 ;
    END
  END EN
  PIN WE[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.630 1396.000 597.910 1400.000 ;
    END
  END WE[0]
  PIN WE[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.430 1396.000 611.710 1400.000 ;
    END
  END WE[1]
  PIN WE[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.770 1396.000 625.050 1400.000 ;
    END
  END WE[2]
  PIN WE[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 638.570 1396.000 638.850 1400.000 ;
    END
  END WE[3]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1387.440 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1387.440 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1387.440 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1387.440 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1387.440 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1387.440 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1387.440 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1387.440 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1387.440 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1387.440 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1387.440 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1387.440 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1387.440 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1387.440 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 1385.785 1094.530 1387.390 ;
        RECT 5.330 1380.345 1094.530 1383.175 ;
        RECT 5.330 1374.905 1094.530 1377.735 ;
        RECT 5.330 1372.245 346.455 1372.295 ;
        RECT 5.330 1369.515 1094.530 1372.245 ;
        RECT 5.330 1369.465 304.595 1369.515 ;
        RECT 5.330 1366.805 161.995 1366.855 ;
        RECT 5.330 1364.075 1094.530 1366.805 ;
        RECT 5.330 1364.025 53.040 1364.075 ;
        RECT 5.330 1361.365 30.500 1361.415 ;
        RECT 5.330 1358.635 1094.530 1361.365 ;
        RECT 5.330 1358.585 78.735 1358.635 ;
        RECT 5.330 1355.925 30.435 1355.975 ;
        RECT 5.330 1353.195 1094.530 1355.925 ;
        RECT 5.330 1353.145 142.215 1353.195 ;
        RECT 5.330 1350.485 31.420 1350.535 ;
        RECT 5.330 1347.755 1094.530 1350.485 ;
        RECT 5.330 1347.705 81.560 1347.755 ;
        RECT 5.330 1345.045 378.195 1345.095 ;
        RECT 5.330 1342.315 1094.530 1345.045 ;
        RECT 5.330 1342.265 219.560 1342.315 ;
        RECT 5.330 1339.605 28.595 1339.655 ;
        RECT 5.330 1336.875 1094.530 1339.605 ;
        RECT 5.330 1336.825 259.975 1336.875 ;
        RECT 5.330 1334.165 28.595 1334.215 ;
        RECT 5.330 1331.435 1094.530 1334.165 ;
        RECT 5.330 1331.385 87.935 1331.435 ;
        RECT 5.330 1328.725 65.855 1328.775 ;
        RECT 5.330 1325.995 1094.530 1328.725 ;
        RECT 5.330 1325.945 111.855 1325.995 ;
        RECT 5.330 1323.285 32.340 1323.335 ;
        RECT 5.330 1320.555 1094.530 1323.285 ;
        RECT 5.330 1320.505 252.615 1320.555 ;
        RECT 5.330 1317.845 297.235 1317.895 ;
        RECT 5.330 1315.115 1094.530 1317.845 ;
        RECT 5.330 1315.065 111.855 1315.115 ;
        RECT 5.330 1312.405 80.575 1312.455 ;
        RECT 5.330 1309.675 1094.530 1312.405 ;
        RECT 5.330 1309.625 23.140 1309.675 ;
        RECT 5.330 1306.965 472.955 1307.015 ;
        RECT 5.330 1304.235 1094.530 1306.965 ;
        RECT 5.330 1304.185 112.315 1304.235 ;
        RECT 5.330 1301.525 29.975 1301.575 ;
        RECT 5.330 1298.795 1094.530 1301.525 ;
        RECT 5.330 1298.745 74.200 1298.795 ;
        RECT 5.330 1296.085 177.635 1296.135 ;
        RECT 5.330 1293.355 1094.530 1296.085 ;
        RECT 5.330 1293.305 47.915 1293.355 ;
        RECT 5.330 1290.645 31.880 1290.695 ;
        RECT 5.330 1287.915 1094.530 1290.645 ;
        RECT 5.330 1287.865 99.500 1287.915 ;
        RECT 5.330 1285.205 28.200 1285.255 ;
        RECT 5.330 1282.475 1094.530 1285.205 ;
        RECT 5.330 1282.425 296.315 1282.475 ;
        RECT 5.330 1279.765 29.055 1279.815 ;
        RECT 5.330 1277.035 1094.530 1279.765 ;
        RECT 5.330 1276.985 245.780 1277.035 ;
        RECT 5.330 1274.325 221.335 1274.375 ;
        RECT 5.330 1271.595 1094.530 1274.325 ;
        RECT 5.330 1271.545 29.120 1271.595 ;
        RECT 5.330 1268.885 115.075 1268.935 ;
        RECT 5.330 1266.155 1094.530 1268.885 ;
        RECT 5.330 1266.105 29.120 1266.155 ;
        RECT 5.330 1263.445 30.435 1263.495 ;
        RECT 5.330 1260.715 1094.530 1263.445 ;
        RECT 5.330 1260.665 77.815 1260.715 ;
        RECT 5.330 1258.005 453.240 1258.055 ;
        RECT 5.330 1255.275 1094.530 1258.005 ;
        RECT 5.330 1255.225 66.840 1255.275 ;
        RECT 5.330 1252.565 140.375 1252.615 ;
        RECT 5.330 1249.835 1094.530 1252.565 ;
        RECT 5.330 1249.785 64.015 1249.835 ;
        RECT 5.330 1247.125 66.840 1247.175 ;
        RECT 5.330 1244.395 1094.530 1247.125 ;
        RECT 5.330 1244.345 182.235 1244.395 ;
        RECT 5.330 1241.685 46.535 1241.735 ;
        RECT 5.330 1238.955 1094.530 1241.685 ;
        RECT 5.330 1238.905 146.815 1238.955 ;
        RECT 5.330 1236.245 31.420 1236.295 ;
        RECT 5.330 1233.515 1094.530 1236.245 ;
        RECT 5.330 1233.465 297.695 1233.515 ;
        RECT 5.330 1230.805 49.360 1230.855 ;
        RECT 5.330 1228.075 1094.530 1230.805 ;
        RECT 5.330 1228.025 65.855 1228.075 ;
        RECT 5.330 1225.365 32.340 1225.415 ;
        RECT 5.330 1222.635 1094.530 1225.365 ;
        RECT 5.330 1222.585 66.840 1222.635 ;
        RECT 5.330 1219.925 30.435 1219.975 ;
        RECT 5.330 1217.195 1094.530 1219.925 ;
        RECT 5.330 1217.145 65.920 1217.195 ;
        RECT 5.330 1214.485 39.635 1214.535 ;
        RECT 5.330 1211.755 1094.530 1214.485 ;
        RECT 5.330 1211.705 96.675 1211.755 ;
        RECT 5.330 1209.045 135.315 1209.095 ;
        RECT 5.330 1206.315 1094.530 1209.045 ;
        RECT 5.330 1206.265 26.295 1206.315 ;
        RECT 5.330 1203.605 29.580 1203.655 ;
        RECT 5.330 1200.875 1094.530 1203.605 ;
        RECT 5.330 1200.825 231.915 1200.875 ;
        RECT 5.330 1198.165 493.195 1198.215 ;
        RECT 5.330 1195.435 1094.530 1198.165 ;
        RECT 5.330 1195.385 340.935 1195.435 ;
        RECT 5.330 1192.725 196.955 1192.775 ;
        RECT 5.330 1189.995 1094.530 1192.725 ;
        RECT 5.330 1189.945 77.420 1189.995 ;
        RECT 5.330 1187.285 81.035 1187.335 ;
        RECT 5.330 1184.555 1094.530 1187.285 ;
        RECT 5.330 1184.505 36.940 1184.555 ;
        RECT 5.330 1181.845 52.055 1181.895 ;
        RECT 5.330 1179.115 1094.530 1181.845 ;
        RECT 5.330 1179.065 227.380 1179.115 ;
        RECT 5.330 1176.405 30.500 1176.455 ;
        RECT 5.330 1173.675 1094.530 1176.405 ;
        RECT 5.330 1173.625 101.340 1173.675 ;
        RECT 5.330 1170.965 343.760 1171.015 ;
        RECT 5.330 1168.235 1094.530 1170.965 ;
        RECT 5.330 1168.185 167.120 1168.235 ;
        RECT 5.330 1165.525 164.295 1165.575 ;
        RECT 5.330 1162.795 1094.530 1165.525 ;
        RECT 5.330 1162.745 47.060 1162.795 ;
        RECT 5.330 1160.085 92.075 1160.135 ;
        RECT 5.330 1157.355 1094.530 1160.085 ;
        RECT 5.330 1157.305 709.920 1157.355 ;
        RECT 5.330 1154.645 81.955 1154.695 ;
        RECT 5.330 1151.915 1094.530 1154.645 ;
        RECT 5.330 1151.865 550.695 1151.915 ;
        RECT 5.330 1149.205 30.500 1149.255 ;
        RECT 5.330 1146.475 1094.530 1149.205 ;
        RECT 5.330 1146.425 33.195 1146.475 ;
        RECT 5.330 1143.765 293.555 1143.815 ;
        RECT 5.330 1141.035 1094.530 1143.765 ;
        RECT 5.330 1140.985 129.335 1141.035 ;
        RECT 5.330 1138.325 50.280 1138.375 ;
        RECT 5.330 1135.595 1094.530 1138.325 ;
        RECT 5.330 1135.545 69.600 1135.595 ;
        RECT 5.330 1132.885 196.035 1132.935 ;
        RECT 5.330 1130.155 1094.530 1132.885 ;
        RECT 5.330 1130.105 68.615 1130.155 ;
        RECT 5.330 1127.445 234.675 1127.495 ;
        RECT 5.330 1124.715 1094.530 1127.445 ;
        RECT 5.330 1124.665 36.940 1124.715 ;
        RECT 5.330 1122.005 54.420 1122.055 ;
        RECT 5.330 1119.275 1094.530 1122.005 ;
        RECT 5.330 1119.225 378.720 1119.275 ;
        RECT 5.330 1116.565 30.040 1116.615 ;
        RECT 5.330 1113.835 1094.530 1116.565 ;
        RECT 5.330 1113.785 174.875 1113.835 ;
        RECT 5.330 1111.125 165.675 1111.175 ;
        RECT 5.330 1108.395 1094.530 1111.125 ;
        RECT 5.330 1108.345 69.995 1108.395 ;
        RECT 5.330 1105.685 31.420 1105.735 ;
        RECT 5.330 1102.955 1094.530 1105.685 ;
        RECT 5.330 1102.905 65.000 1102.955 ;
        RECT 5.330 1100.245 492.275 1100.295 ;
        RECT 5.330 1097.515 1094.530 1100.245 ;
        RECT 5.330 1097.465 411.380 1097.515 ;
        RECT 5.330 1094.805 417.755 1094.855 ;
        RECT 5.330 1092.075 1094.530 1094.805 ;
        RECT 5.330 1092.025 460.995 1092.075 ;
        RECT 5.330 1089.365 580.595 1089.415 ;
        RECT 5.330 1086.635 1094.530 1089.365 ;
        RECT 5.330 1086.585 460.995 1086.635 ;
        RECT 5.330 1083.925 511.135 1083.975 ;
        RECT 5.330 1081.195 1094.530 1083.925 ;
        RECT 5.330 1081.145 433.855 1081.195 ;
        RECT 5.330 1078.485 7.895 1078.535 ;
        RECT 5.330 1075.755 1094.530 1078.485 ;
        RECT 5.330 1075.705 39.240 1075.755 ;
        RECT 5.330 1073.045 52.055 1073.095 ;
        RECT 5.330 1070.315 1094.530 1073.045 ;
        RECT 5.330 1070.265 26.820 1070.315 ;
        RECT 5.330 1067.605 157.855 1067.655 ;
        RECT 5.330 1064.875 1094.530 1067.605 ;
        RECT 5.330 1064.825 52.515 1064.875 ;
        RECT 5.330 1062.165 106.795 1062.215 ;
        RECT 5.330 1059.435 1094.530 1062.165 ;
        RECT 5.330 1059.385 236.055 1059.435 ;
        RECT 5.330 1056.725 39.635 1056.775 ;
        RECT 5.330 1053.995 1094.530 1056.725 ;
        RECT 5.330 1053.945 10.720 1053.995 ;
        RECT 5.330 1051.285 257.675 1051.335 ;
        RECT 5.330 1048.555 1094.530 1051.285 ;
        RECT 5.330 1048.505 25.835 1048.555 ;
        RECT 5.330 1045.845 38.255 1045.895 ;
        RECT 5.330 1043.115 1094.530 1045.845 ;
        RECT 5.330 1043.065 92.995 1043.115 ;
        RECT 5.330 1040.405 35.495 1040.455 ;
        RECT 5.330 1037.675 1094.530 1040.405 ;
        RECT 5.330 1037.625 69.535 1037.675 ;
        RECT 5.330 1034.965 24.060 1035.015 ;
        RECT 5.330 1032.235 1094.530 1034.965 ;
        RECT 5.330 1032.185 271.015 1032.235 ;
        RECT 5.330 1029.525 104.495 1029.575 ;
        RECT 5.330 1026.795 1094.530 1029.525 ;
        RECT 5.330 1026.745 93.455 1026.795 ;
        RECT 5.330 1024.085 23.075 1024.135 ;
        RECT 5.330 1021.355 1094.530 1024.085 ;
        RECT 5.330 1021.305 94.375 1021.355 ;
        RECT 5.330 1018.645 39.635 1018.695 ;
        RECT 5.330 1015.915 1094.530 1018.645 ;
        RECT 5.330 1015.865 41.015 1015.915 ;
        RECT 5.330 1013.205 20.775 1013.255 ;
        RECT 5.330 1010.475 1094.530 1013.205 ;
        RECT 5.330 1010.425 34.115 1010.475 ;
        RECT 5.330 1007.765 23.140 1007.815 ;
        RECT 5.330 1005.035 1094.530 1007.765 ;
        RECT 5.330 1004.985 169.355 1005.035 ;
        RECT 5.330 1002.325 165.740 1002.375 ;
        RECT 5.330 999.595 1094.530 1002.325 ;
        RECT 5.330 999.545 167.055 999.595 ;
        RECT 5.330 996.885 245.255 996.935 ;
        RECT 5.330 994.155 1094.530 996.885 ;
        RECT 5.330 994.105 127.955 994.155 ;
        RECT 5.330 991.445 246.240 991.495 ;
        RECT 5.330 988.715 1094.530 991.445 ;
        RECT 5.330 988.665 123.815 988.715 ;
        RECT 5.330 986.005 221.335 986.055 ;
        RECT 5.330 983.275 1094.530 986.005 ;
        RECT 5.330 983.225 125.260 983.275 ;
        RECT 5.330 980.565 345.995 980.615 ;
        RECT 5.330 977.835 1094.530 980.565 ;
        RECT 5.330 977.785 24.060 977.835 ;
        RECT 5.330 975.125 104.955 975.175 ;
        RECT 5.330 972.395 1094.530 975.125 ;
        RECT 5.330 972.345 35.495 972.395 ;
        RECT 5.330 969.685 54.355 969.735 ;
        RECT 5.330 966.955 1094.530 969.685 ;
        RECT 5.330 966.905 98.055 966.955 ;
        RECT 5.330 964.245 10.720 964.295 ;
        RECT 5.330 961.515 1094.530 964.245 ;
        RECT 5.330 961.465 73.215 961.515 ;
        RECT 5.330 958.805 39.635 958.855 ;
        RECT 5.330 956.075 1094.530 958.805 ;
        RECT 5.330 956.025 10.720 956.075 ;
        RECT 5.330 953.365 36.020 953.415 ;
        RECT 5.330 950.635 1094.530 953.365 ;
        RECT 5.330 950.585 314.715 950.635 ;
        RECT 5.330 947.925 533.280 947.975 ;
        RECT 5.330 945.195 1094.530 947.925 ;
        RECT 5.330 945.145 291.320 945.195 ;
        RECT 5.330 942.485 160.155 942.535 ;
        RECT 5.330 939.755 1094.530 942.485 ;
        RECT 5.330 939.705 20.840 939.755 ;
        RECT 5.330 937.045 51.595 937.095 ;
        RECT 5.330 934.315 1094.530 937.045 ;
        RECT 5.330 934.265 54.420 934.315 ;
        RECT 5.330 931.605 187.295 931.655 ;
        RECT 5.330 928.875 1094.530 931.605 ;
        RECT 5.330 928.825 272.460 928.875 ;
        RECT 5.330 926.165 346.915 926.215 ;
        RECT 5.330 923.435 1094.530 926.165 ;
        RECT 5.330 923.385 144.975 923.435 ;
        RECT 5.330 920.725 241.180 920.775 ;
        RECT 5.330 917.995 1094.530 920.725 ;
        RECT 5.330 917.945 379.575 917.995 ;
        RECT 5.330 915.285 109.620 915.335 ;
        RECT 5.330 912.555 1094.530 915.285 ;
        RECT 5.330 912.505 78.735 912.555 ;
        RECT 5.330 909.845 107.715 909.895 ;
        RECT 5.330 907.115 1094.530 909.845 ;
        RECT 5.330 907.065 72.820 907.115 ;
        RECT 5.330 904.405 109.160 904.455 ;
        RECT 5.330 901.675 1094.530 904.405 ;
        RECT 5.330 901.625 45.680 901.675 ;
        RECT 5.330 898.965 23.600 899.015 ;
        RECT 5.330 896.235 1094.530 898.965 ;
        RECT 5.330 896.185 23.140 896.235 ;
        RECT 5.330 893.525 49.360 893.575 ;
        RECT 5.330 890.795 1094.530 893.525 ;
        RECT 5.330 890.745 60.335 890.795 ;
        RECT 5.330 888.085 376.355 888.135 ;
        RECT 5.330 885.355 1094.530 888.085 ;
        RECT 5.330 885.305 403.035 885.355 ;
        RECT 5.330 882.645 619.300 882.695 ;
        RECT 5.330 879.915 1094.530 882.645 ;
        RECT 5.330 879.865 550.695 879.915 ;
        RECT 5.330 877.205 161.995 877.255 ;
        RECT 5.330 874.475 1094.530 877.205 ;
        RECT 5.330 874.425 23.995 874.475 ;
        RECT 5.330 871.765 25.440 871.815 ;
        RECT 5.330 869.035 1094.530 871.765 ;
        RECT 5.330 868.985 29.120 869.035 ;
        RECT 5.330 866.325 86.095 866.375 ;
        RECT 5.330 863.595 1094.530 866.325 ;
        RECT 5.330 863.545 52.515 863.595 ;
        RECT 5.330 860.885 297.300 860.935 ;
        RECT 5.330 858.155 1094.530 860.885 ;
        RECT 5.330 858.105 34.575 858.155 ;
        RECT 5.330 855.445 24.915 855.495 ;
        RECT 5.330 852.715 1094.530 855.445 ;
        RECT 5.330 852.665 29.120 852.715 ;
        RECT 5.330 850.005 144.515 850.055 ;
        RECT 5.330 847.275 1094.530 850.005 ;
        RECT 5.330 847.225 75.580 847.275 ;
        RECT 5.330 844.565 103.640 844.615 ;
        RECT 5.330 841.835 1094.530 844.565 ;
        RECT 5.330 841.785 78.735 841.835 ;
        RECT 5.330 839.125 308.735 839.175 ;
        RECT 5.330 836.395 1094.530 839.125 ;
        RECT 5.330 836.345 7.895 836.395 ;
        RECT 5.330 833.685 65.855 833.735 ;
        RECT 5.330 830.955 1094.530 833.685 ;
        RECT 5.330 830.905 160.220 830.955 ;
        RECT 5.330 828.245 267.335 828.295 ;
        RECT 5.330 825.515 1094.530 828.245 ;
        RECT 5.330 825.465 35.035 825.515 ;
        RECT 5.330 822.805 272.000 822.855 ;
        RECT 5.330 820.075 1094.530 822.805 ;
        RECT 5.330 820.025 22.155 820.075 ;
        RECT 5.330 817.365 24.520 817.415 ;
        RECT 5.330 814.635 1094.530 817.365 ;
        RECT 5.330 814.585 463.755 814.635 ;
        RECT 5.330 811.925 308.735 811.975 ;
        RECT 5.330 809.195 1094.530 811.925 ;
        RECT 5.330 809.145 352.895 809.195 ;
        RECT 5.330 806.485 107.255 806.535 ;
        RECT 5.330 803.755 1094.530 806.485 ;
        RECT 5.330 803.705 105.480 803.755 ;
        RECT 5.330 801.045 53.960 801.095 ;
        RECT 5.330 798.315 1094.530 801.045 ;
        RECT 5.330 798.265 36.940 798.315 ;
        RECT 5.330 795.605 235.135 795.655 ;
        RECT 5.330 792.875 1094.530 795.605 ;
        RECT 5.330 792.825 629.355 792.875 ;
        RECT 5.330 790.165 300.915 790.215 ;
        RECT 5.330 787.435 1094.530 790.165 ;
        RECT 5.330 787.385 111.855 787.435 ;
        RECT 5.330 784.725 107.255 784.775 ;
        RECT 5.330 781.995 1094.530 784.725 ;
        RECT 5.330 781.945 22.220 781.995 ;
        RECT 5.330 779.285 32.275 779.335 ;
        RECT 5.330 776.555 1094.530 779.285 ;
        RECT 5.330 776.505 74.595 776.555 ;
        RECT 5.330 773.845 223.175 773.895 ;
        RECT 5.330 771.115 1094.530 773.845 ;
        RECT 5.330 771.065 307.815 771.115 ;
        RECT 5.330 768.405 293.160 768.455 ;
        RECT 5.330 765.675 1094.530 768.405 ;
        RECT 5.330 765.625 410.855 765.675 ;
        RECT 5.330 762.965 256.295 763.015 ;
        RECT 5.330 760.235 1094.530 762.965 ;
        RECT 5.330 760.185 19.855 760.235 ;
        RECT 5.330 757.525 38.715 757.575 ;
        RECT 5.330 754.795 1094.530 757.525 ;
        RECT 5.330 754.745 85.635 754.795 ;
        RECT 5.330 752.085 7.895 752.135 ;
        RECT 5.330 749.355 1094.530 752.085 ;
        RECT 5.330 749.305 48.375 749.355 ;
        RECT 5.330 746.645 51.135 746.695 ;
        RECT 5.330 743.915 1094.530 746.645 ;
        RECT 5.330 743.865 39.700 743.915 ;
        RECT 5.330 741.205 10.720 741.255 ;
        RECT 5.330 738.475 1094.530 741.205 ;
        RECT 5.330 738.425 227.315 738.475 ;
        RECT 5.330 735.765 223.700 735.815 ;
        RECT 5.330 733.035 1094.530 735.765 ;
        RECT 5.330 732.985 119.215 733.035 ;
        RECT 5.330 730.325 224.160 730.375 ;
        RECT 5.330 727.595 1094.530 730.325 ;
        RECT 5.330 727.545 75.515 727.595 ;
        RECT 5.330 724.885 7.895 724.935 ;
        RECT 5.330 722.155 1094.530 724.885 ;
        RECT 5.330 722.105 103.115 722.155 ;
        RECT 5.330 719.445 154.700 719.495 ;
        RECT 5.330 716.715 1094.530 719.445 ;
        RECT 5.330 716.665 25.440 716.715 ;
        RECT 5.330 714.005 38.780 714.055 ;
        RECT 5.330 711.275 1094.530 714.005 ;
        RECT 5.330 711.225 52.055 711.275 ;
        RECT 5.330 708.565 20.775 708.615 ;
        RECT 5.330 705.835 1094.530 708.565 ;
        RECT 5.330 705.785 86.095 705.835 ;
        RECT 5.330 703.125 226.000 703.175 ;
        RECT 5.330 700.395 1094.530 703.125 ;
        RECT 5.330 700.345 69.995 700.395 ;
        RECT 5.330 697.685 428.795 697.735 ;
        RECT 5.330 694.955 1094.530 697.685 ;
        RECT 5.330 694.905 7.895 694.955 ;
        RECT 5.330 692.245 225.080 692.295 ;
        RECT 5.330 689.515 1094.530 692.245 ;
        RECT 5.330 689.465 25.440 689.515 ;
        RECT 5.330 686.805 179.015 686.855 ;
        RECT 5.330 684.075 1094.530 686.805 ;
        RECT 5.330 684.025 103.115 684.075 ;
        RECT 5.330 681.365 39.700 681.415 ;
        RECT 5.330 678.635 1094.530 681.365 ;
        RECT 5.330 678.585 51.660 678.635 ;
        RECT 5.330 675.925 49.755 675.975 ;
        RECT 5.330 673.195 1094.530 675.925 ;
        RECT 5.330 673.145 245.780 673.195 ;
        RECT 5.330 670.485 39.175 670.535 ;
        RECT 5.330 667.755 1094.530 670.485 ;
        RECT 5.330 667.705 123.815 667.755 ;
        RECT 5.330 665.045 46.535 665.095 ;
        RECT 5.330 662.315 1094.530 665.045 ;
        RECT 5.330 662.265 7.895 662.315 ;
        RECT 5.330 659.605 232.900 659.655 ;
        RECT 5.330 656.875 1094.530 659.605 ;
        RECT 5.330 656.825 387.920 656.875 ;
        RECT 5.330 654.165 390.615 654.215 ;
        RECT 5.330 651.435 1094.530 654.165 ;
        RECT 5.330 651.385 575.075 651.435 ;
        RECT 5.330 648.725 278.440 648.775 ;
        RECT 5.330 645.995 1094.530 648.725 ;
        RECT 5.330 645.945 311.955 645.995 ;
        RECT 5.330 643.285 251.760 643.335 ;
        RECT 5.330 640.555 1094.530 643.285 ;
        RECT 5.330 640.505 254.980 640.555 ;
        RECT 5.330 637.845 222.320 637.895 ;
        RECT 5.330 635.115 1094.530 637.845 ;
        RECT 5.330 635.065 363.475 635.115 ;
        RECT 5.330 632.405 577.835 632.455 ;
        RECT 5.330 629.675 1094.530 632.405 ;
        RECT 5.330 629.625 445.815 629.675 ;
        RECT 5.330 626.965 362.095 627.015 ;
        RECT 5.330 624.235 1094.530 626.965 ;
        RECT 5.330 624.185 401.195 624.235 ;
        RECT 5.330 621.525 39.700 621.575 ;
        RECT 5.330 618.795 1094.530 621.525 ;
        RECT 5.330 618.745 69.995 618.795 ;
        RECT 5.330 616.085 35.560 616.135 ;
        RECT 5.330 613.355 1094.530 616.085 ;
        RECT 5.330 613.305 47.455 613.355 ;
        RECT 5.330 610.645 28.595 610.695 ;
        RECT 5.330 607.915 1094.530 610.645 ;
        RECT 5.330 607.865 7.895 607.915 ;
        RECT 5.330 605.205 204.775 605.255 ;
        RECT 5.330 602.475 1094.530 605.205 ;
        RECT 5.330 602.425 61.715 602.475 ;
        RECT 5.330 599.765 47.455 599.815 ;
        RECT 5.330 597.035 1094.530 599.765 ;
        RECT 5.330 596.985 24.980 597.035 ;
        RECT 5.330 594.325 784.835 594.375 ;
        RECT 5.330 591.595 1094.530 594.325 ;
        RECT 5.330 591.545 77.355 591.595 ;
        RECT 5.330 588.885 291.255 588.935 ;
        RECT 5.330 586.155 1094.530 588.885 ;
        RECT 5.330 586.105 173.955 586.155 ;
        RECT 5.330 583.445 75.580 583.495 ;
        RECT 5.330 580.715 1094.530 583.445 ;
        RECT 5.330 580.665 27.280 580.715 ;
        RECT 5.330 578.005 7.895 578.055 ;
        RECT 5.330 575.275 1094.530 578.005 ;
        RECT 5.330 575.225 341.920 575.275 ;
        RECT 5.330 572.565 23.600 572.615 ;
        RECT 5.330 569.835 1094.530 572.565 ;
        RECT 5.330 569.785 35.955 569.835 ;
        RECT 5.330 567.125 83.335 567.175 ;
        RECT 5.330 564.395 1094.530 567.125 ;
        RECT 5.330 564.345 68.220 564.395 ;
        RECT 5.330 561.685 65.000 561.735 ;
        RECT 5.330 558.955 1094.530 561.685 ;
        RECT 5.330 558.905 111.855 558.955 ;
        RECT 5.330 556.245 164.755 556.295 ;
        RECT 5.330 553.515 1094.530 556.245 ;
        RECT 5.330 553.465 7.895 553.515 ;
        RECT 5.330 550.805 87.080 550.855 ;
        RECT 5.330 548.075 1094.530 550.805 ;
        RECT 5.330 548.025 97.595 548.075 ;
        RECT 5.330 545.365 192.815 545.415 ;
        RECT 5.330 542.635 1094.530 545.365 ;
        RECT 5.330 542.585 190.515 542.635 ;
        RECT 5.330 539.925 39.635 539.975 ;
        RECT 5.330 537.195 1094.530 539.925 ;
        RECT 5.330 537.145 43.380 537.195 ;
        RECT 5.330 534.485 7.895 534.535 ;
        RECT 5.330 531.755 1094.530 534.485 ;
        RECT 5.330 531.705 429.320 531.755 ;
        RECT 5.330 529.045 173.560 529.095 ;
        RECT 5.330 526.315 1094.530 529.045 ;
        RECT 5.330 526.265 169.815 526.315 ;
        RECT 5.330 523.605 7.895 523.655 ;
        RECT 5.330 520.875 1094.530 523.605 ;
        RECT 5.330 520.825 76.895 520.875 ;
        RECT 5.330 518.165 23.995 518.215 ;
        RECT 5.330 515.435 1094.530 518.165 ;
        RECT 5.330 515.385 296.315 515.435 ;
        RECT 5.330 512.725 54.880 512.775 ;
        RECT 5.330 509.995 1094.530 512.725 ;
        RECT 5.330 509.945 191.435 509.995 ;
        RECT 5.330 507.285 248.540 507.335 ;
        RECT 5.330 504.555 1094.530 507.285 ;
        RECT 5.330 504.505 103.640 504.555 ;
        RECT 5.330 501.845 432.935 501.895 ;
        RECT 5.330 499.115 1094.530 501.845 ;
        RECT 5.330 499.065 98.580 499.115 ;
        RECT 5.330 496.405 72.755 496.455 ;
        RECT 5.330 493.675 1094.530 496.405 ;
        RECT 5.330 493.625 36.415 493.675 ;
        RECT 5.330 490.965 7.895 491.015 ;
        RECT 5.330 488.235 1094.530 490.965 ;
        RECT 5.330 488.185 21.695 488.235 ;
        RECT 5.330 485.525 101.800 485.575 ;
        RECT 5.330 482.795 1094.530 485.525 ;
        RECT 5.330 482.745 70.520 482.795 ;
        RECT 5.330 480.085 230.075 480.135 ;
        RECT 5.330 477.355 1094.530 480.085 ;
        RECT 5.330 477.305 988.615 477.355 ;
        RECT 5.330 474.645 351.120 474.695 ;
        RECT 5.330 471.915 1094.530 474.645 ;
        RECT 5.330 471.865 123.815 471.915 ;
        RECT 5.330 469.205 7.895 469.255 ;
        RECT 5.330 466.475 1094.530 469.205 ;
        RECT 5.330 466.425 28.200 466.475 ;
        RECT 5.330 463.765 65.000 463.815 ;
        RECT 5.330 461.035 1094.530 463.765 ;
        RECT 5.330 460.985 343.300 461.035 ;
        RECT 5.330 458.325 30.435 458.375 ;
        RECT 5.330 455.595 1094.530 458.325 ;
        RECT 5.330 455.545 107.780 455.595 ;
        RECT 5.330 452.885 126.115 452.935 ;
        RECT 5.330 450.155 1094.530 452.885 ;
        RECT 5.330 450.105 164.295 450.155 ;
        RECT 5.330 447.445 125.195 447.495 ;
        RECT 5.330 444.715 1094.530 447.445 ;
        RECT 5.330 444.665 7.895 444.715 ;
        RECT 5.330 442.005 296.315 442.055 ;
        RECT 5.330 439.275 1094.530 442.005 ;
        RECT 5.330 439.225 64.080 439.275 ;
        RECT 5.330 436.565 50.740 436.615 ;
        RECT 5.330 433.835 1094.530 436.565 ;
        RECT 5.330 433.785 68.155 433.835 ;
        RECT 5.330 431.125 230.075 431.175 ;
        RECT 5.330 428.395 1094.530 431.125 ;
        RECT 5.330 428.345 100.880 428.395 ;
        RECT 5.330 425.685 21.235 425.735 ;
        RECT 5.330 422.955 1094.530 425.685 ;
        RECT 5.330 422.905 45.220 422.955 ;
        RECT 5.330 420.245 282.515 420.295 ;
        RECT 5.330 417.515 1094.530 420.245 ;
        RECT 5.330 417.465 43.380 417.515 ;
        RECT 5.330 414.805 73.215 414.855 ;
        RECT 5.330 412.075 1094.530 414.805 ;
        RECT 5.330 412.025 41.475 412.075 ;
        RECT 5.330 409.365 7.895 409.415 ;
        RECT 5.330 406.635 1094.530 409.365 ;
        RECT 5.330 406.585 71.440 406.635 ;
        RECT 5.330 403.925 492.275 403.975 ;
        RECT 5.330 401.195 1094.530 403.925 ;
        RECT 5.330 401.145 24.520 401.195 ;
        RECT 5.330 398.485 177.635 398.535 ;
        RECT 5.330 395.755 1094.530 398.485 ;
        RECT 5.330 395.705 122.895 395.755 ;
        RECT 5.330 393.045 125.195 393.095 ;
        RECT 5.330 390.315 1094.530 393.045 ;
        RECT 5.330 390.265 25.375 390.315 ;
        RECT 5.330 387.605 81.495 387.655 ;
        RECT 5.330 384.875 1094.530 387.605 ;
        RECT 5.330 384.825 69.600 384.875 ;
        RECT 5.330 382.165 394.755 382.215 ;
        RECT 5.330 379.435 1094.530 382.165 ;
        RECT 5.330 379.385 38.255 379.435 ;
        RECT 5.330 376.725 10.720 376.775 ;
        RECT 5.330 373.995 1094.530 376.725 ;
        RECT 5.330 373.945 53.960 373.995 ;
        RECT 5.330 371.285 261.815 371.335 ;
        RECT 5.330 368.555 1094.530 371.285 ;
        RECT 5.330 368.505 527.300 368.555 ;
        RECT 5.330 365.845 128.020 365.895 ;
        RECT 5.330 363.115 1094.530 365.845 ;
        RECT 5.330 363.065 179.015 363.115 ;
        RECT 5.330 360.405 7.895 360.455 ;
        RECT 5.330 357.675 1094.530 360.405 ;
        RECT 5.330 357.625 37.400 357.675 ;
        RECT 5.330 354.965 101.800 355.015 ;
        RECT 5.330 352.235 1094.530 354.965 ;
        RECT 5.330 352.185 574.615 352.235 ;
        RECT 5.330 349.525 528.220 349.575 ;
        RECT 5.330 346.795 1094.530 349.525 ;
        RECT 5.330 346.745 648.215 346.795 ;
        RECT 5.330 344.085 728.255 344.135 ;
        RECT 5.330 341.355 1094.530 344.085 ;
        RECT 5.330 341.305 545.175 341.355 ;
        RECT 5.330 338.645 526.775 338.695 ;
        RECT 5.330 335.915 1094.530 338.645 ;
        RECT 5.330 335.865 326.215 335.915 ;
        RECT 5.330 333.205 426.035 333.255 ;
        RECT 5.330 330.475 1094.530 333.205 ;
        RECT 5.330 330.425 403.100 330.475 ;
        RECT 5.330 327.765 448.115 327.815 ;
        RECT 5.330 325.035 1094.530 327.765 ;
        RECT 5.330 324.985 140.835 325.035 ;
        RECT 5.330 322.325 91.155 322.375 ;
        RECT 5.330 319.595 1094.530 322.325 ;
        RECT 5.330 319.545 21.760 319.595 ;
        RECT 5.330 316.885 22.155 316.935 ;
        RECT 5.330 314.155 1094.530 316.885 ;
        RECT 5.330 314.105 25.900 314.155 ;
        RECT 5.330 311.445 22.155 311.495 ;
        RECT 5.330 308.715 1094.530 311.445 ;
        RECT 5.330 308.665 112.775 308.715 ;
        RECT 5.330 306.005 65.855 306.055 ;
        RECT 5.330 303.275 1094.530 306.005 ;
        RECT 5.330 303.225 69.600 303.275 ;
        RECT 5.330 300.565 129.795 300.615 ;
        RECT 5.330 297.835 1094.530 300.565 ;
        RECT 5.330 297.785 192.355 297.835 ;
        RECT 5.330 295.125 210.755 295.175 ;
        RECT 5.330 292.395 1094.530 295.125 ;
        RECT 5.330 292.345 40.095 292.395 ;
        RECT 5.330 289.685 106.795 289.735 ;
        RECT 5.330 286.955 1094.530 289.685 ;
        RECT 5.330 286.905 262.275 286.955 ;
        RECT 5.330 284.245 24.520 284.295 ;
        RECT 5.330 281.515 1094.530 284.245 ;
        RECT 5.330 281.465 22.615 281.515 ;
        RECT 5.330 278.805 39.635 278.855 ;
        RECT 5.330 276.075 1094.530 278.805 ;
        RECT 5.330 276.025 26.360 276.075 ;
        RECT 5.330 273.365 314.780 273.415 ;
        RECT 5.330 270.635 1094.530 273.365 ;
        RECT 5.330 270.585 104.955 270.635 ;
        RECT 5.330 267.925 27.675 267.975 ;
        RECT 5.330 265.195 1094.530 267.925 ;
        RECT 5.330 265.145 78.735 265.195 ;
        RECT 5.330 262.485 203.855 262.535 ;
        RECT 5.330 259.755 1094.530 262.485 ;
        RECT 5.330 259.705 223.700 259.755 ;
        RECT 5.330 257.045 343.695 257.095 ;
        RECT 5.330 254.315 1094.530 257.045 ;
        RECT 5.330 254.265 23.995 254.315 ;
        RECT 5.330 251.605 24.980 251.655 ;
        RECT 5.330 248.875 1094.530 251.605 ;
        RECT 5.330 248.825 100.420 248.875 ;
        RECT 5.330 246.165 29.515 246.215 ;
        RECT 5.330 243.435 1094.530 246.165 ;
        RECT 5.330 243.385 151.415 243.435 ;
        RECT 5.330 237.995 1094.530 240.775 ;
        RECT 5.330 237.945 24.520 237.995 ;
        RECT 5.330 235.285 91.615 235.335 ;
        RECT 5.330 232.555 1094.530 235.285 ;
        RECT 5.330 232.505 74.200 232.555 ;
        RECT 5.330 229.845 68.680 229.895 ;
        RECT 5.330 227.115 1094.530 229.845 ;
        RECT 5.330 227.065 177.635 227.115 ;
        RECT 5.330 224.405 144.515 224.455 ;
        RECT 5.330 221.675 1094.530 224.405 ;
        RECT 5.330 221.625 198.795 221.675 ;
        RECT 5.330 218.965 247.555 219.015 ;
        RECT 5.330 216.235 1094.530 218.965 ;
        RECT 5.330 216.185 306.500 216.235 ;
        RECT 5.330 213.525 37.860 213.575 ;
        RECT 5.330 210.795 1094.530 213.525 ;
        RECT 5.330 210.745 35.955 210.795 ;
        RECT 5.330 208.085 26.820 208.135 ;
        RECT 5.330 205.355 1094.530 208.085 ;
        RECT 5.330 205.305 115.535 205.355 ;
        RECT 5.330 202.645 65.460 202.695 ;
        RECT 5.330 199.915 1094.530 202.645 ;
        RECT 5.330 199.865 78.275 199.915 ;
        RECT 5.330 197.205 113.695 197.255 ;
        RECT 5.330 194.475 1094.530 197.205 ;
        RECT 5.330 194.425 24.980 194.475 ;
        RECT 5.330 191.765 90.695 191.815 ;
        RECT 5.330 189.035 1094.530 191.765 ;
        RECT 5.330 188.985 200.175 189.035 ;
        RECT 5.330 186.325 687.775 186.375 ;
        RECT 5.330 183.595 1094.530 186.325 ;
        RECT 5.330 183.545 200.175 183.595 ;
        RECT 5.330 180.885 212.595 180.935 ;
        RECT 5.330 178.155 1094.530 180.885 ;
        RECT 5.330 178.105 18.935 178.155 ;
        RECT 5.330 175.445 92.075 175.495 ;
        RECT 5.330 172.715 1094.530 175.445 ;
        RECT 5.330 172.665 576.520 172.715 ;
        RECT 5.330 170.005 29.975 170.055 ;
        RECT 5.330 167.275 1094.530 170.005 ;
        RECT 5.330 167.225 29.120 167.275 ;
        RECT 5.330 164.565 267.795 164.615 ;
        RECT 5.330 161.835 1094.530 164.565 ;
        RECT 5.330 161.785 29.120 161.835 ;
        RECT 5.330 159.125 29.055 159.175 ;
        RECT 5.330 156.395 1094.530 159.125 ;
        RECT 5.330 156.345 317.540 156.395 ;
        RECT 5.330 153.685 138.535 153.735 ;
        RECT 5.330 150.955 1094.530 153.685 ;
        RECT 5.330 150.905 139.455 150.955 ;
        RECT 5.330 148.245 67.300 148.295 ;
        RECT 5.330 145.515 1094.530 148.245 ;
        RECT 5.330 145.465 171.655 145.515 ;
        RECT 5.330 142.805 65.855 142.855 ;
        RECT 5.330 140.075 1094.530 142.805 ;
        RECT 5.330 140.025 26.820 140.075 ;
        RECT 5.330 137.365 92.075 137.415 ;
        RECT 5.330 134.635 1094.530 137.365 ;
        RECT 5.330 134.585 26.360 134.635 ;
        RECT 5.330 131.925 262.275 131.975 ;
        RECT 5.330 129.195 1094.530 131.925 ;
        RECT 5.330 129.145 317.540 129.195 ;
        RECT 5.330 126.485 85.700 126.535 ;
        RECT 5.330 123.755 1094.530 126.485 ;
        RECT 5.330 123.705 62.240 123.755 ;
        RECT 5.330 121.045 58.955 121.095 ;
        RECT 5.330 118.315 1094.530 121.045 ;
        RECT 5.330 118.265 27.740 118.315 ;
        RECT 5.330 115.605 60.860 115.655 ;
        RECT 5.330 112.875 1094.530 115.605 ;
        RECT 5.330 112.825 193.275 112.875 ;
        RECT 5.330 110.165 27.675 110.215 ;
        RECT 5.330 107.435 1094.530 110.165 ;
        RECT 5.330 107.385 28.660 107.435 ;
        RECT 5.330 104.725 113.300 104.775 ;
        RECT 5.330 101.995 1094.530 104.725 ;
        RECT 5.330 101.945 254.455 101.995 ;
        RECT 5.330 99.285 158.775 99.335 ;
        RECT 5.330 96.555 1094.530 99.285 ;
        RECT 5.330 96.505 26.295 96.555 ;
        RECT 5.330 93.845 590.255 93.895 ;
        RECT 5.330 91.115 1094.530 93.845 ;
        RECT 5.330 91.065 99.960 91.115 ;
        RECT 5.330 88.405 141.295 88.455 ;
        RECT 5.330 85.675 1094.530 88.405 ;
        RECT 5.330 85.625 47.520 85.675 ;
        RECT 5.330 82.965 92.075 83.015 ;
        RECT 5.330 80.235 1094.530 82.965 ;
        RECT 5.330 80.185 47.520 80.235 ;
        RECT 5.330 77.525 29.120 77.575 ;
        RECT 5.330 74.795 1094.530 77.525 ;
        RECT 5.330 74.745 667.140 74.795 ;
        RECT 5.330 72.085 131.175 72.135 ;
        RECT 5.330 69.355 1094.530 72.085 ;
        RECT 5.330 69.305 175.335 69.355 ;
        RECT 5.330 66.645 128.020 66.695 ;
        RECT 5.330 63.915 1094.530 66.645 ;
        RECT 5.330 63.865 148.195 63.915 ;
        RECT 5.330 61.205 39.635 61.255 ;
        RECT 5.330 58.475 1094.530 61.205 ;
        RECT 5.330 58.425 59.415 58.475 ;
        RECT 5.330 55.765 28.200 55.815 ;
        RECT 5.330 53.035 1094.530 55.765 ;
        RECT 5.330 52.985 116.455 53.035 ;
        RECT 5.330 50.325 81.035 50.375 ;
        RECT 5.330 47.595 1094.530 50.325 ;
        RECT 5.330 47.545 203.395 47.595 ;
        RECT 5.330 44.885 77.880 44.935 ;
        RECT 5.330 42.155 1094.530 44.885 ;
        RECT 5.330 42.105 19.920 42.155 ;
        RECT 5.330 39.445 23.140 39.495 ;
        RECT 5.330 36.715 1094.530 39.445 ;
        RECT 5.330 36.665 93.455 36.715 ;
        RECT 5.330 34.005 57.115 34.055 ;
        RECT 5.330 31.275 1094.530 34.005 ;
        RECT 5.330 31.225 18.475 31.275 ;
        RECT 5.330 28.565 20.315 28.615 ;
        RECT 5.330 25.835 1094.530 28.565 ;
        RECT 5.330 25.785 307.420 25.835 ;
        RECT 5.330 20.345 1094.530 23.175 ;
        RECT 5.330 14.905 1094.530 17.735 ;
        RECT 5.330 10.690 1094.530 12.295 ;
      LAYER li1 ;
        RECT 5.520 10.795 1095.115 1387.285 ;
      LAYER met1 ;
        RECT 5.520 9.560 1095.175 1387.440 ;
      LAYER met2 ;
        RECT 7.090 1395.720 19.590 1396.000 ;
        RECT 20.430 1395.720 33.390 1396.000 ;
        RECT 34.230 1395.720 47.190 1396.000 ;
        RECT 48.030 1395.720 60.990 1396.000 ;
        RECT 61.830 1395.720 74.790 1396.000 ;
        RECT 75.630 1395.720 88.590 1396.000 ;
        RECT 89.430 1395.720 102.390 1396.000 ;
        RECT 103.230 1395.720 116.190 1396.000 ;
        RECT 117.030 1395.720 129.530 1396.000 ;
        RECT 130.370 1395.720 143.330 1396.000 ;
        RECT 144.170 1395.720 157.130 1396.000 ;
        RECT 157.970 1395.720 170.930 1396.000 ;
        RECT 171.770 1395.720 184.730 1396.000 ;
        RECT 185.570 1395.720 198.530 1396.000 ;
        RECT 199.370 1395.720 212.330 1396.000 ;
        RECT 213.170 1395.720 226.130 1396.000 ;
        RECT 226.970 1395.720 239.930 1396.000 ;
        RECT 240.770 1395.720 253.270 1396.000 ;
        RECT 254.110 1395.720 267.070 1396.000 ;
        RECT 267.910 1395.720 280.870 1396.000 ;
        RECT 281.710 1395.720 294.670 1396.000 ;
        RECT 295.510 1395.720 308.470 1396.000 ;
        RECT 309.310 1395.720 322.270 1396.000 ;
        RECT 323.110 1395.720 336.070 1396.000 ;
        RECT 336.910 1395.720 349.870 1396.000 ;
        RECT 350.710 1395.720 363.670 1396.000 ;
        RECT 364.510 1395.720 377.010 1396.000 ;
        RECT 377.850 1395.720 390.810 1396.000 ;
        RECT 391.650 1395.720 404.610 1396.000 ;
        RECT 405.450 1395.720 418.410 1396.000 ;
        RECT 419.250 1395.720 432.210 1396.000 ;
        RECT 433.050 1395.720 446.010 1396.000 ;
        RECT 446.850 1395.720 459.810 1396.000 ;
        RECT 460.650 1395.720 473.610 1396.000 ;
        RECT 474.450 1395.720 487.410 1396.000 ;
        RECT 488.250 1395.720 500.750 1396.000 ;
        RECT 501.590 1395.720 514.550 1396.000 ;
        RECT 515.390 1395.720 528.350 1396.000 ;
        RECT 529.190 1395.720 542.150 1396.000 ;
        RECT 542.990 1395.720 555.950 1396.000 ;
        RECT 556.790 1395.720 569.750 1396.000 ;
        RECT 570.590 1395.720 583.550 1396.000 ;
        RECT 584.390 1395.720 597.350 1396.000 ;
        RECT 598.190 1395.720 611.150 1396.000 ;
        RECT 611.990 1395.720 624.490 1396.000 ;
        RECT 625.330 1395.720 638.290 1396.000 ;
        RECT 639.130 1395.720 652.090 1396.000 ;
        RECT 652.930 1395.720 665.890 1396.000 ;
        RECT 666.730 1395.720 679.690 1396.000 ;
        RECT 680.530 1395.720 693.490 1396.000 ;
        RECT 694.330 1395.720 707.290 1396.000 ;
        RECT 708.130 1395.720 721.090 1396.000 ;
        RECT 721.930 1395.720 734.890 1396.000 ;
        RECT 735.730 1395.720 748.230 1396.000 ;
        RECT 749.070 1395.720 762.030 1396.000 ;
        RECT 762.870 1395.720 775.830 1396.000 ;
        RECT 776.670 1395.720 789.630 1396.000 ;
        RECT 790.470 1395.720 803.430 1396.000 ;
        RECT 804.270 1395.720 817.230 1396.000 ;
        RECT 818.070 1395.720 831.030 1396.000 ;
        RECT 831.870 1395.720 844.830 1396.000 ;
        RECT 845.670 1395.720 858.630 1396.000 ;
        RECT 859.470 1395.720 871.970 1396.000 ;
        RECT 872.810 1395.720 885.770 1396.000 ;
        RECT 886.610 1395.720 899.570 1396.000 ;
        RECT 900.410 1395.720 913.370 1396.000 ;
        RECT 914.210 1395.720 927.170 1396.000 ;
        RECT 928.010 1395.720 940.970 1396.000 ;
        RECT 941.810 1395.720 954.770 1396.000 ;
        RECT 955.610 1395.720 968.570 1396.000 ;
        RECT 969.410 1395.720 982.370 1396.000 ;
        RECT 983.210 1395.720 995.710 1396.000 ;
        RECT 996.550 1395.720 1009.510 1396.000 ;
        RECT 1010.350 1395.720 1023.310 1396.000 ;
        RECT 1024.150 1395.720 1037.110 1396.000 ;
        RECT 1037.950 1395.720 1050.910 1396.000 ;
        RECT 1051.750 1395.720 1064.710 1396.000 ;
        RECT 1065.550 1395.720 1078.510 1396.000 ;
        RECT 1079.350 1395.720 1092.310 1396.000 ;
        RECT 1093.150 1395.720 1093.320 1396.000 ;
        RECT 6.540 9.530 1093.320 1395.720 ;
      LAYER met3 ;
        RECT 6.965 10.715 1092.895 1387.365 ;
      LAYER met4 ;
        RECT 19.615 43.015 20.640 1384.985 ;
        RECT 23.040 43.015 97.440 1384.985 ;
        RECT 99.840 43.015 174.240 1384.985 ;
        RECT 176.640 43.015 251.040 1384.985 ;
        RECT 253.440 43.015 327.840 1384.985 ;
        RECT 330.240 43.015 404.640 1384.985 ;
        RECT 407.040 43.015 481.440 1384.985 ;
        RECT 483.840 43.015 558.240 1384.985 ;
        RECT 560.640 43.015 635.040 1384.985 ;
        RECT 637.440 43.015 711.840 1384.985 ;
        RECT 714.240 43.015 788.640 1384.985 ;
        RECT 791.040 43.015 865.440 1384.985 ;
        RECT 867.840 43.015 942.240 1384.985 ;
        RECT 944.640 43.015 1019.040 1384.985 ;
        RECT 1021.440 43.015 1083.465 1384.985 ;
  END
END DFFRAM_4K
END LIBRARY

