VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO DFFRAM_1Kx32
  CLASS BLOCK ;
  FOREIGN DFFRAM_1Kx32 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1100.000 BY 1400.000 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.290 1396.000 446.570 1400.000 ;
    END
  END A[0]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.090 1396.000 460.370 1400.000 ;
    END
  END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.890 1396.000 474.170 1400.000 ;
    END
  END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.690 1396.000 487.970 1400.000 ;
    END
  END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.030 1396.000 501.310 1400.000 ;
    END
  END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.830 1396.000 515.110 1400.000 ;
    END
  END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.630 1396.000 528.910 1400.000 ;
    END
  END A[6]
  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.430 1396.000 542.710 1400.000 ;
    END
  END A[7]
  PIN A[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.230 1396.000 556.510 1400.000 ;
    END
  END A[8]
  PIN A[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.030 1396.000 570.310 1400.000 ;
    END
  END A[9]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 583.830 1396.000 584.110 1400.000 ;
    END
  END CLK
  PIN Di[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.170 1396.000 666.450 1400.000 ;
    END
  END Di[0]
  PIN Di[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 803.710 1396.000 803.990 1400.000 ;
    END
  END Di[10]
  PIN Di[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.510 1396.000 817.790 1400.000 ;
    END
  END Di[11]
  PIN Di[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 831.310 1396.000 831.590 1400.000 ;
    END
  END Di[12]
  PIN Di[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 845.110 1396.000 845.390 1400.000 ;
    END
  END Di[13]
  PIN Di[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 858.910 1396.000 859.190 1400.000 ;
    END
  END Di[14]
  PIN Di[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 872.250 1396.000 872.530 1400.000 ;
    END
  END Di[15]
  PIN Di[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 886.050 1396.000 886.330 1400.000 ;
    END
  END Di[16]
  PIN Di[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 899.850 1396.000 900.130 1400.000 ;
    END
  END Di[17]
  PIN Di[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 913.650 1396.000 913.930 1400.000 ;
    END
  END Di[18]
  PIN Di[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.450 1396.000 927.730 1400.000 ;
    END
  END Di[19]
  PIN Di[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.970 1396.000 680.250 1400.000 ;
    END
  END Di[1]
  PIN Di[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 941.250 1396.000 941.530 1400.000 ;
    END
  END Di[20]
  PIN Di[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 955.050 1396.000 955.330 1400.000 ;
    END
  END Di[21]
  PIN Di[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 968.850 1396.000 969.130 1400.000 ;
    END
  END Di[22]
  PIN Di[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 982.650 1396.000 982.930 1400.000 ;
    END
  END Di[23]
  PIN Di[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.990 1396.000 996.270 1400.000 ;
    END
  END Di[24]
  PIN Di[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1009.790 1396.000 1010.070 1400.000 ;
    END
  END Di[25]
  PIN Di[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1023.590 1396.000 1023.870 1400.000 ;
    END
  END Di[26]
  PIN Di[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1037.390 1396.000 1037.670 1400.000 ;
    END
  END Di[27]
  PIN Di[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1051.190 1396.000 1051.470 1400.000 ;
    END
  END Di[28]
  PIN Di[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1064.990 1396.000 1065.270 1400.000 ;
    END
  END Di[29]
  PIN Di[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 693.770 1396.000 694.050 1400.000 ;
    END
  END Di[2]
  PIN Di[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1078.790 1396.000 1079.070 1400.000 ;
    END
  END Di[30]
  PIN Di[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1092.590 1396.000 1092.870 1400.000 ;
    END
  END Di[31]
  PIN Di[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.570 1396.000 707.850 1400.000 ;
    END
  END Di[3]
  PIN Di[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.370 1396.000 721.650 1400.000 ;
    END
  END Di[4]
  PIN Di[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.170 1396.000 735.450 1400.000 ;
    END
  END Di[5]
  PIN Di[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.510 1396.000 748.790 1400.000 ;
    END
  END Di[6]
  PIN Di[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 762.310 1396.000 762.590 1400.000 ;
    END
  END Di[7]
  PIN Di[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.110 1396.000 776.390 1400.000 ;
    END
  END Di[8]
  PIN Di[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.910 1396.000 790.190 1400.000 ;
    END
  END Di[9]
  PIN Do[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 1396.000 6.810 1400.000 ;
    END
  END Do[0]
  PIN Do[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 1396.000 143.890 1400.000 ;
    END
  END Do[10]
  PIN Do[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.410 1396.000 157.690 1400.000 ;
    END
  END Do[11]
  PIN Do[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.210 1396.000 171.490 1400.000 ;
    END
  END Do[12]
  PIN Do[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 1396.000 185.290 1400.000 ;
    END
  END Do[13]
  PIN Do[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.810 1396.000 199.090 1400.000 ;
    END
  END Do[14]
  PIN Do[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 1396.000 212.890 1400.000 ;
    END
  END Do[15]
  PIN Do[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 1396.000 226.690 1400.000 ;
    END
  END Do[16]
  PIN Do[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.210 1396.000 240.490 1400.000 ;
    END
  END Do[17]
  PIN Do[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.550 1396.000 253.830 1400.000 ;
    END
  END Do[18]
  PIN Do[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 1396.000 267.630 1400.000 ;
    END
  END Do[19]
  PIN Do[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 1396.000 20.150 1400.000 ;
    END
  END Do[1]
  PIN Do[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.150 1396.000 281.430 1400.000 ;
    END
  END Do[20]
  PIN Do[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.950 1396.000 295.230 1400.000 ;
    END
  END Do[21]
  PIN Do[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.750 1396.000 309.030 1400.000 ;
    END
  END Do[22]
  PIN Do[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.550 1396.000 322.830 1400.000 ;
    END
  END Do[23]
  PIN Do[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.350 1396.000 336.630 1400.000 ;
    END
  END Do[24]
  PIN Do[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.150 1396.000 350.430 1400.000 ;
    END
  END Do[25]
  PIN Do[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 1396.000 364.230 1400.000 ;
    END
  END Do[26]
  PIN Do[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.290 1396.000 377.570 1400.000 ;
    END
  END Do[27]
  PIN Do[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.090 1396.000 391.370 1400.000 ;
    END
  END Do[28]
  PIN Do[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.890 1396.000 405.170 1400.000 ;
    END
  END Do[29]
  PIN Do[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 1396.000 33.950 1400.000 ;
    END
  END Do[2]
  PIN Do[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 1396.000 418.970 1400.000 ;
    END
  END Do[30]
  PIN Do[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.490 1396.000 432.770 1400.000 ;
    END
  END Do[31]
  PIN Do[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 1396.000 47.750 1400.000 ;
    END
  END Do[3]
  PIN Do[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 1396.000 61.550 1400.000 ;
    END
  END Do[4]
  PIN Do[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 1396.000 75.350 1400.000 ;
    END
  END Do[5]
  PIN Do[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 1396.000 89.150 1400.000 ;
    END
  END Do[6]
  PIN Do[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.670 1396.000 102.950 1400.000 ;
    END
  END Do[7]
  PIN Do[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.470 1396.000 116.750 1400.000 ;
    END
  END Do[8]
  PIN Do[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 1396.000 130.090 1400.000 ;
    END
  END Do[9]
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.370 1396.000 652.650 1400.000 ;
    END
  END EN
  PIN WE[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.630 1396.000 597.910 1400.000 ;
    END
  END WE[0]
  PIN WE[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.430 1396.000 611.710 1400.000 ;
    END
  END WE[1]
  PIN WE[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.770 1396.000 625.050 1400.000 ;
    END
  END WE[2]
  PIN WE[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 638.570 1396.000 638.850 1400.000 ;
    END
  END WE[3]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1387.440 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1387.440 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1387.440 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1387.440 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1387.440 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1387.440 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1387.440 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1387.440 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1387.440 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1387.440 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1387.440 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1387.440 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1387.440 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1387.440 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 1385.785 1094.530 1387.390 ;
        RECT 5.330 1380.345 1094.530 1383.175 ;
        RECT 5.330 1374.905 1094.530 1377.735 ;
        RECT 5.330 1369.515 1094.530 1372.295 ;
        RECT 5.330 1369.465 454.555 1369.515 ;
        RECT 5.330 1366.805 327.660 1366.855 ;
        RECT 5.330 1364.075 1094.530 1366.805 ;
        RECT 5.330 1364.025 114.680 1364.075 ;
        RECT 5.330 1361.365 274.695 1361.415 ;
        RECT 5.330 1358.635 1094.530 1361.365 ;
        RECT 5.330 1358.585 127.035 1358.635 ;
        RECT 5.330 1355.925 106.335 1355.975 ;
        RECT 5.330 1353.195 1094.530 1355.925 ;
        RECT 5.330 1353.145 176.255 1353.195 ;
        RECT 5.330 1350.485 42.460 1350.535 ;
        RECT 5.330 1347.755 1094.530 1350.485 ;
        RECT 5.330 1347.705 36.480 1347.755 ;
        RECT 5.330 1345.045 86.095 1345.095 ;
        RECT 5.330 1342.315 1094.530 1345.045 ;
        RECT 5.330 1342.265 21.760 1342.315 ;
        RECT 5.330 1339.605 24.520 1339.655 ;
        RECT 5.330 1336.875 1094.530 1339.605 ;
        RECT 5.330 1336.825 25.900 1336.875 ;
        RECT 5.330 1334.165 115.535 1334.215 ;
        RECT 5.330 1331.435 1094.530 1334.165 ;
        RECT 5.330 1331.385 89.775 1331.435 ;
        RECT 5.330 1328.725 284.355 1328.775 ;
        RECT 5.330 1325.995 1094.530 1328.725 ;
        RECT 5.330 1325.945 69.075 1325.995 ;
        RECT 5.330 1323.285 222.715 1323.335 ;
        RECT 5.330 1320.555 1094.530 1323.285 ;
        RECT 5.330 1320.505 179.080 1320.555 ;
        RECT 5.330 1317.845 241.115 1317.895 ;
        RECT 5.330 1315.115 1094.530 1317.845 ;
        RECT 5.330 1315.065 23.600 1315.115 ;
        RECT 5.330 1312.405 84.715 1312.455 ;
        RECT 5.330 1309.675 1094.530 1312.405 ;
        RECT 5.330 1309.625 40.555 1309.675 ;
        RECT 5.330 1306.965 59.940 1307.015 ;
        RECT 5.330 1304.235 1094.530 1306.965 ;
        RECT 5.330 1304.185 41.540 1304.235 ;
        RECT 5.330 1301.525 24.980 1301.575 ;
        RECT 5.330 1298.795 1094.530 1301.525 ;
        RECT 5.330 1298.745 236.055 1298.795 ;
        RECT 5.330 1296.085 184.075 1296.135 ;
        RECT 5.330 1293.355 1094.530 1296.085 ;
        RECT 5.330 1293.305 236.055 1293.355 ;
        RECT 5.330 1290.645 25.440 1290.695 ;
        RECT 5.330 1287.915 1094.530 1290.645 ;
        RECT 5.330 1287.865 72.360 1287.915 ;
        RECT 5.330 1285.205 24.915 1285.255 ;
        RECT 5.330 1282.475 1094.530 1285.205 ;
        RECT 5.330 1282.425 185.520 1282.475 ;
        RECT 5.330 1279.765 206.680 1279.815 ;
        RECT 5.330 1277.035 1094.530 1279.765 ;
        RECT 5.330 1276.985 128.415 1277.035 ;
        RECT 5.330 1274.325 184.995 1274.375 ;
        RECT 5.330 1271.595 1094.530 1274.325 ;
        RECT 5.330 1271.545 49.820 1271.595 ;
        RECT 5.330 1268.885 85.175 1268.935 ;
        RECT 5.330 1266.155 1094.530 1268.885 ;
        RECT 5.330 1266.105 27.280 1266.155 ;
        RECT 5.330 1263.445 180.460 1263.495 ;
        RECT 5.330 1260.715 1094.530 1263.445 ;
        RECT 5.330 1260.665 114.155 1260.715 ;
        RECT 5.330 1258.005 344.155 1258.055 ;
        RECT 5.330 1255.275 1094.530 1258.005 ;
        RECT 5.330 1255.225 99.435 1255.275 ;
        RECT 5.330 1252.565 267.795 1252.615 ;
        RECT 5.330 1249.835 1094.530 1252.565 ;
        RECT 5.330 1249.785 22.615 1249.835 ;
        RECT 5.330 1247.125 24.520 1247.175 ;
        RECT 5.330 1244.395 1094.530 1247.125 ;
        RECT 5.330 1244.345 45.155 1244.395 ;
        RECT 5.330 1241.685 130.715 1241.735 ;
        RECT 5.330 1238.955 1094.530 1241.685 ;
        RECT 5.330 1238.905 49.820 1238.955 ;
        RECT 5.330 1236.245 64.015 1236.295 ;
        RECT 5.330 1233.515 1094.530 1236.245 ;
        RECT 5.330 1233.465 111.855 1233.515 ;
        RECT 5.330 1230.805 35.495 1230.855 ;
        RECT 5.330 1228.075 1094.530 1230.805 ;
        RECT 5.330 1228.025 85.635 1228.075 ;
        RECT 5.330 1225.365 23.140 1225.415 ;
        RECT 5.330 1222.635 1094.530 1225.365 ;
        RECT 5.330 1222.585 243.415 1222.635 ;
        RECT 5.330 1219.925 180.460 1219.975 ;
        RECT 5.330 1217.195 1094.530 1219.925 ;
        RECT 5.330 1217.145 21.300 1217.195 ;
        RECT 5.330 1214.485 224.620 1214.535 ;
        RECT 5.330 1211.755 1094.530 1214.485 ;
        RECT 5.330 1211.705 85.635 1211.755 ;
        RECT 5.330 1209.045 32.340 1209.095 ;
        RECT 5.330 1206.315 1094.530 1209.045 ;
        RECT 5.330 1206.265 62.240 1206.315 ;
        RECT 5.330 1203.605 118.360 1203.655 ;
        RECT 5.330 1200.875 1094.530 1203.605 ;
        RECT 5.330 1200.825 115.535 1200.875 ;
        RECT 5.330 1198.165 24.520 1198.215 ;
        RECT 5.330 1195.435 1094.530 1198.165 ;
        RECT 5.330 1195.385 45.220 1195.435 ;
        RECT 5.330 1192.725 116.455 1192.775 ;
        RECT 5.330 1189.995 1094.530 1192.725 ;
        RECT 5.330 1189.945 105.940 1189.995 ;
        RECT 5.330 1187.285 46.535 1187.335 ;
        RECT 5.330 1184.555 1094.530 1187.285 ;
        RECT 5.330 1184.505 847.855 1184.555 ;
        RECT 5.330 1181.845 28.660 1181.895 ;
        RECT 5.330 1179.115 1094.530 1181.845 ;
        RECT 5.330 1179.065 886.560 1179.115 ;
        RECT 5.330 1176.405 115.995 1176.455 ;
        RECT 5.330 1173.675 1094.530 1176.405 ;
        RECT 5.330 1173.625 48.375 1173.675 ;
        RECT 5.330 1170.965 101.735 1171.015 ;
        RECT 5.330 1168.235 1094.530 1170.965 ;
        RECT 5.330 1168.185 25.440 1168.235 ;
        RECT 5.330 1165.525 222.715 1165.575 ;
        RECT 5.330 1162.795 1094.530 1165.525 ;
        RECT 5.330 1162.745 78.735 1162.795 ;
        RECT 5.330 1160.085 974.880 1160.135 ;
        RECT 5.330 1157.355 1094.530 1160.085 ;
        RECT 5.330 1157.305 24.915 1157.355 ;
        RECT 5.330 1154.645 23.075 1154.695 ;
        RECT 5.330 1151.915 1094.530 1154.645 ;
        RECT 5.330 1151.865 21.760 1151.915 ;
        RECT 5.330 1149.205 108.635 1149.255 ;
        RECT 5.330 1146.475 1094.530 1149.205 ;
        RECT 5.330 1146.425 25.900 1146.475 ;
        RECT 5.330 1143.765 82.415 1143.815 ;
        RECT 5.330 1141.035 1094.530 1143.765 ;
        RECT 5.330 1140.985 21.760 1141.035 ;
        RECT 5.330 1138.325 125.195 1138.375 ;
        RECT 5.330 1135.595 1094.530 1138.325 ;
        RECT 5.330 1135.545 62.240 1135.595 ;
        RECT 5.330 1132.885 205.235 1132.935 ;
        RECT 5.330 1130.155 1094.530 1132.885 ;
        RECT 5.330 1130.105 426.495 1130.155 ;
        RECT 5.330 1127.445 355.720 1127.495 ;
        RECT 5.330 1124.715 1094.530 1127.445 ;
        RECT 5.330 1124.665 142.215 1124.715 ;
        RECT 5.330 1122.005 64.080 1122.055 ;
        RECT 5.330 1119.275 1094.530 1122.005 ;
        RECT 5.330 1119.225 408.555 1119.275 ;
        RECT 5.330 1116.565 49.360 1116.615 ;
        RECT 5.330 1113.835 1094.530 1116.565 ;
        RECT 5.330 1113.785 52.580 1113.835 ;
        RECT 5.330 1111.125 623.375 1111.175 ;
        RECT 5.330 1108.395 1094.530 1111.125 ;
        RECT 5.330 1108.345 186.440 1108.395 ;
        RECT 5.330 1105.685 614.635 1105.735 ;
        RECT 5.330 1102.955 1094.530 1105.685 ;
        RECT 5.330 1102.905 235.135 1102.955 ;
        RECT 5.330 1100.245 214.895 1100.295 ;
        RECT 5.330 1097.515 1094.530 1100.245 ;
        RECT 5.330 1097.465 183.615 1097.515 ;
        RECT 5.330 1094.805 354.340 1094.855 ;
        RECT 5.330 1092.075 1094.530 1094.805 ;
        RECT 5.330 1092.025 206.220 1092.075 ;
        RECT 5.330 1089.365 347.440 1089.415 ;
        RECT 5.330 1086.635 1094.530 1089.365 ;
        RECT 5.330 1086.585 176.255 1086.635 ;
        RECT 5.330 1083.925 221.860 1083.975 ;
        RECT 5.330 1081.195 1094.530 1083.925 ;
        RECT 5.330 1081.145 178.620 1081.195 ;
        RECT 5.330 1078.485 522.175 1078.535 ;
        RECT 5.330 1075.755 1094.530 1078.485 ;
        RECT 5.330 1075.705 514.420 1075.755 ;
        RECT 5.330 1073.045 957.335 1073.095 ;
        RECT 5.330 1070.315 1094.530 1073.045 ;
        RECT 5.330 1070.265 92.535 1070.315 ;
        RECT 5.330 1067.605 125.195 1067.655 ;
        RECT 5.330 1064.875 1094.530 1067.605 ;
        RECT 5.330 1064.825 54.880 1064.875 ;
        RECT 5.330 1062.165 23.140 1062.215 ;
        RECT 5.330 1059.435 1094.530 1062.165 ;
        RECT 5.330 1059.385 26.295 1059.435 ;
        RECT 5.330 1056.725 418.215 1056.775 ;
        RECT 5.330 1053.995 1094.530 1056.725 ;
        RECT 5.330 1053.945 363.475 1053.995 ;
        RECT 5.330 1051.285 330.880 1051.335 ;
        RECT 5.330 1048.555 1094.530 1051.285 ;
        RECT 5.330 1048.505 21.760 1048.555 ;
        RECT 5.330 1045.845 485.440 1045.895 ;
        RECT 5.330 1043.115 1094.530 1045.845 ;
        RECT 5.330 1043.065 24.915 1043.115 ;
        RECT 5.330 1040.405 49.360 1040.455 ;
        RECT 5.330 1037.675 1094.530 1040.405 ;
        RECT 5.330 1037.625 69.995 1037.675 ;
        RECT 5.330 1034.965 72.755 1035.015 ;
        RECT 5.330 1032.235 1094.530 1034.965 ;
        RECT 5.330 1032.185 27.740 1032.235 ;
        RECT 5.330 1029.525 267.335 1029.575 ;
        RECT 5.330 1026.795 1094.530 1029.525 ;
        RECT 5.330 1026.745 329.895 1026.795 ;
        RECT 5.330 1024.085 249.920 1024.135 ;
        RECT 5.330 1021.355 1094.530 1024.085 ;
        RECT 5.330 1021.305 68.155 1021.355 ;
        RECT 5.330 1018.645 26.820 1018.695 ;
        RECT 5.330 1015.915 1094.530 1018.645 ;
        RECT 5.330 1015.865 25.375 1015.915 ;
        RECT 5.330 1013.205 46.995 1013.255 ;
        RECT 5.330 1010.475 1094.530 1013.205 ;
        RECT 5.330 1010.425 380.955 1010.475 ;
        RECT 5.330 1007.765 686.920 1007.815 ;
        RECT 5.330 1005.035 1094.530 1007.765 ;
        RECT 5.330 1004.985 186.440 1005.035 ;
        RECT 5.330 1002.325 162.915 1002.375 ;
        RECT 5.330 999.595 1094.530 1002.325 ;
        RECT 5.330 999.545 329.895 999.595 ;
        RECT 5.330 996.885 196.955 996.935 ;
        RECT 5.330 994.155 1094.530 996.885 ;
        RECT 5.330 994.105 351.120 994.155 ;
        RECT 5.330 991.445 112.315 991.495 ;
        RECT 5.330 988.715 1094.530 991.445 ;
        RECT 5.330 988.665 53.040 988.715 ;
        RECT 5.330 986.005 58.560 986.055 ;
        RECT 5.330 983.275 1094.530 986.005 ;
        RECT 5.330 983.225 27.740 983.275 ;
        RECT 5.330 980.565 23.600 980.615 ;
        RECT 5.330 977.835 1094.530 980.565 ;
        RECT 5.330 977.785 28.660 977.835 ;
        RECT 5.330 975.125 983.555 975.175 ;
        RECT 5.330 972.395 1094.530 975.125 ;
        RECT 5.330 972.345 71.375 972.395 ;
        RECT 5.330 969.685 28.595 969.735 ;
        RECT 5.330 966.955 1094.530 969.685 ;
        RECT 5.330 966.905 202.540 966.955 ;
        RECT 5.330 964.245 108.175 964.295 ;
        RECT 5.330 961.515 1094.530 964.245 ;
        RECT 5.330 961.465 21.760 961.515 ;
        RECT 5.330 958.805 23.140 958.855 ;
        RECT 5.330 956.075 1094.530 958.805 ;
        RECT 5.330 956.025 334.100 956.075 ;
        RECT 5.330 953.365 185.455 953.415 ;
        RECT 5.330 950.635 1094.530 953.365 ;
        RECT 5.330 950.585 70.915 950.635 ;
        RECT 5.330 947.925 25.440 947.975 ;
        RECT 5.330 945.195 1094.530 947.925 ;
        RECT 5.330 945.145 204.840 945.195 ;
        RECT 5.330 942.485 52.580 942.535 ;
        RECT 5.330 939.755 1094.530 942.485 ;
        RECT 5.330 939.705 27.740 939.755 ;
        RECT 5.330 937.045 162.060 937.095 ;
        RECT 5.330 934.315 1094.530 937.045 ;
        RECT 5.330 934.265 254.060 934.315 ;
        RECT 5.330 931.605 49.360 931.655 ;
        RECT 5.330 928.875 1094.530 931.605 ;
        RECT 5.330 928.825 60.795 928.875 ;
        RECT 5.330 926.165 106.795 926.215 ;
        RECT 5.330 923.435 1094.530 926.165 ;
        RECT 5.330 923.385 419.135 923.435 ;
        RECT 5.330 920.725 59.415 920.775 ;
        RECT 5.330 917.995 1094.530 920.725 ;
        RECT 5.330 917.945 26.360 917.995 ;
        RECT 5.330 915.285 23.140 915.335 ;
        RECT 5.330 912.555 1094.530 915.285 ;
        RECT 5.330 912.505 249.855 912.555 ;
        RECT 5.330 909.845 92.075 909.895 ;
        RECT 5.330 907.115 1094.530 909.845 ;
        RECT 5.330 907.065 186.440 907.115 ;
        RECT 5.330 904.405 167.975 904.455 ;
        RECT 5.330 901.675 1094.530 904.405 ;
        RECT 5.330 901.625 22.680 901.675 ;
        RECT 5.330 898.965 64.015 899.015 ;
        RECT 5.330 896.235 1094.530 898.965 ;
        RECT 5.330 896.185 127.495 896.235 ;
        RECT 5.330 893.525 346.980 893.575 ;
        RECT 5.330 890.795 1094.530 893.525 ;
        RECT 5.330 890.745 217.655 890.795 ;
        RECT 5.330 888.085 345.075 888.135 ;
        RECT 5.330 885.355 1094.530 888.085 ;
        RECT 5.330 885.305 28.200 885.355 ;
        RECT 5.330 882.645 78.735 882.695 ;
        RECT 5.330 879.915 1094.530 882.645 ;
        RECT 5.330 879.865 28.660 879.915 ;
        RECT 5.330 877.205 29.975 877.255 ;
        RECT 5.330 874.475 1094.530 877.205 ;
        RECT 5.330 874.425 114.680 874.475 ;
        RECT 5.330 871.765 186.375 871.815 ;
        RECT 5.330 869.035 1094.530 871.765 ;
        RECT 5.330 868.985 24.915 869.035 ;
        RECT 5.330 866.325 267.335 866.375 ;
        RECT 5.330 863.595 1094.530 866.325 ;
        RECT 5.330 863.545 219.035 863.595 ;
        RECT 5.330 860.885 161.075 860.935 ;
        RECT 5.330 858.155 1094.530 860.885 ;
        RECT 5.330 858.105 586.575 858.155 ;
        RECT 5.330 855.445 233.755 855.495 ;
        RECT 5.330 852.715 1094.530 855.445 ;
        RECT 5.330 852.665 167.120 852.715 ;
        RECT 5.330 850.005 173.560 850.055 ;
        RECT 5.330 847.275 1094.530 850.005 ;
        RECT 5.330 847.225 482.680 847.275 ;
        RECT 5.330 844.565 24.520 844.615 ;
        RECT 5.330 841.835 1094.530 844.565 ;
        RECT 5.330 841.785 53.040 841.835 ;
        RECT 5.330 839.125 25.375 839.175 ;
        RECT 5.330 836.395 1094.530 839.125 ;
        RECT 5.330 836.345 28.660 836.395 ;
        RECT 5.330 833.685 265.035 833.735 ;
        RECT 5.330 830.955 1094.530 833.685 ;
        RECT 5.330 830.905 71.375 830.955 ;
        RECT 5.330 828.245 652.420 828.295 ;
        RECT 5.330 825.515 1094.530 828.245 ;
        RECT 5.330 825.465 483.140 825.515 ;
        RECT 5.330 822.805 164.360 822.855 ;
        RECT 5.330 820.075 1094.530 822.805 ;
        RECT 5.330 820.025 71.835 820.075 ;
        RECT 5.330 817.365 32.800 817.415 ;
        RECT 5.330 814.635 1094.530 817.365 ;
        RECT 5.330 814.585 238.420 814.635 ;
        RECT 5.330 811.925 104.955 811.975 ;
        RECT 5.330 809.195 1094.530 811.925 ;
        RECT 5.330 809.145 87.015 809.195 ;
        RECT 5.330 806.485 30.500 806.535 ;
        RECT 5.330 803.755 1094.530 806.485 ;
        RECT 5.330 803.705 48.900 803.755 ;
        RECT 5.330 801.045 29.055 801.095 ;
        RECT 5.330 798.315 1094.530 801.045 ;
        RECT 5.330 798.265 20.775 798.315 ;
        RECT 5.330 795.605 88.395 795.655 ;
        RECT 5.330 792.875 1094.530 795.605 ;
        RECT 5.330 792.825 166.135 792.875 ;
        RECT 5.330 790.165 23.140 790.215 ;
        RECT 5.330 787.435 1094.530 790.165 ;
        RECT 5.330 787.385 182.235 787.435 ;
        RECT 5.330 784.725 348.755 784.775 ;
        RECT 5.330 781.995 1094.530 784.725 ;
        RECT 5.330 781.945 218.115 781.995 ;
        RECT 5.330 779.285 182.300 779.335 ;
        RECT 5.330 776.555 1094.530 779.285 ;
        RECT 5.330 776.505 201.095 776.555 ;
        RECT 5.330 773.845 337.780 773.895 ;
        RECT 5.330 771.115 1094.530 773.845 ;
        RECT 5.330 771.065 350.595 771.115 ;
        RECT 5.330 768.405 188.675 768.455 ;
        RECT 5.330 765.675 1094.530 768.405 ;
        RECT 5.330 765.625 452.715 765.675 ;
        RECT 5.330 762.965 806.915 763.015 ;
        RECT 5.330 760.235 1094.530 762.965 ;
        RECT 5.330 760.185 574.155 760.235 ;
        RECT 5.330 757.525 275.615 757.575 ;
        RECT 5.330 754.795 1094.530 757.525 ;
        RECT 5.330 754.745 332.655 754.795 ;
        RECT 5.330 752.085 248.015 752.135 ;
        RECT 5.330 749.355 1094.530 752.085 ;
        RECT 5.330 749.305 49.755 749.355 ;
        RECT 5.330 746.645 24.980 746.695 ;
        RECT 5.330 743.915 1094.530 746.645 ;
        RECT 5.330 743.865 25.440 743.915 ;
        RECT 5.330 741.205 105.875 741.255 ;
        RECT 5.330 738.475 1094.530 741.205 ;
        RECT 5.330 738.425 311.560 738.475 ;
        RECT 5.330 735.765 317.935 735.815 ;
        RECT 5.330 733.035 1094.530 735.765 ;
        RECT 5.330 732.985 295.395 733.035 ;
        RECT 5.330 730.325 68.680 730.375 ;
        RECT 5.330 727.595 1094.530 730.325 ;
        RECT 5.330 727.545 26.295 727.595 ;
        RECT 5.330 724.885 89.775 724.935 ;
        RECT 5.330 722.155 1094.530 724.885 ;
        RECT 5.330 722.105 27.740 722.155 ;
        RECT 5.330 719.445 57.115 719.495 ;
        RECT 5.330 716.715 1094.530 719.445 ;
        RECT 5.330 716.665 129.795 716.715 ;
        RECT 5.330 714.005 690.995 714.055 ;
        RECT 5.330 711.275 1094.530 714.005 ;
        RECT 5.330 711.225 24.520 711.275 ;
        RECT 5.330 708.565 115.535 708.615 ;
        RECT 5.330 705.835 1094.530 708.565 ;
        RECT 5.330 705.785 25.440 705.835 ;
        RECT 5.330 703.125 90.235 703.175 ;
        RECT 5.330 700.395 1094.530 703.125 ;
        RECT 5.330 700.345 298.220 700.395 ;
        RECT 5.330 697.685 30.895 697.735 ;
        RECT 5.330 694.955 1094.530 697.685 ;
        RECT 5.330 694.905 350.135 694.955 ;
        RECT 5.330 692.245 285.340 692.295 ;
        RECT 5.330 689.515 1094.530 692.245 ;
        RECT 5.330 689.465 71.375 689.515 ;
        RECT 5.330 686.805 278.440 686.855 ;
        RECT 5.330 684.075 1094.530 686.805 ;
        RECT 5.330 684.025 21.760 684.075 ;
        RECT 5.330 681.365 75.580 681.415 ;
        RECT 5.330 678.635 1094.530 681.365 ;
        RECT 5.330 678.585 123.815 678.635 ;
        RECT 5.330 675.925 107.255 675.975 ;
        RECT 5.330 673.195 1094.530 675.925 ;
        RECT 5.330 673.145 25.375 673.195 ;
        RECT 5.330 670.485 65.460 670.535 ;
        RECT 5.330 667.755 1094.530 670.485 ;
        RECT 5.330 667.705 640.000 667.755 ;
        RECT 5.330 665.045 728.255 665.095 ;
        RECT 5.330 662.315 1094.530 665.045 ;
        RECT 5.330 662.265 353.355 662.315 ;
        RECT 5.330 659.605 161.995 659.655 ;
        RECT 5.330 656.875 1094.530 659.605 ;
        RECT 5.330 656.825 75.515 656.875 ;
        RECT 5.330 654.165 309.655 654.215 ;
        RECT 5.330 651.435 1094.530 654.165 ;
        RECT 5.330 651.385 252.615 651.435 ;
        RECT 5.330 648.725 194.720 648.775 ;
        RECT 5.330 645.995 1094.530 648.725 ;
        RECT 5.330 645.945 20.840 645.995 ;
        RECT 5.330 643.285 76.960 643.335 ;
        RECT 5.330 640.555 1094.530 643.285 ;
        RECT 5.330 640.505 23.140 640.555 ;
        RECT 5.330 637.845 26.295 637.895 ;
        RECT 5.330 635.115 1094.530 637.845 ;
        RECT 5.330 635.065 459.615 635.115 ;
        RECT 5.330 632.405 24.455 632.455 ;
        RECT 5.330 629.675 1094.530 632.405 ;
        RECT 5.330 629.625 26.360 629.675 ;
        RECT 5.330 626.965 75.580 627.015 ;
        RECT 5.330 624.235 1094.530 626.965 ;
        RECT 5.330 624.185 28.200 624.235 ;
        RECT 5.330 621.525 25.900 621.575 ;
        RECT 5.330 618.795 1094.530 621.525 ;
        RECT 5.330 618.745 430.700 618.795 ;
        RECT 5.330 616.085 189.200 616.135 ;
        RECT 5.330 613.355 1094.530 616.085 ;
        RECT 5.330 613.305 254.915 613.355 ;
        RECT 5.330 610.645 431.620 610.695 ;
        RECT 5.330 607.915 1094.530 610.645 ;
        RECT 5.330 607.865 498.255 607.915 ;
        RECT 5.330 605.205 56.655 605.255 ;
        RECT 5.330 602.475 1094.530 605.205 ;
        RECT 5.330 602.425 24.980 602.475 ;
        RECT 5.330 599.765 130.715 599.815 ;
        RECT 5.330 597.035 1094.530 599.765 ;
        RECT 5.330 596.985 87.475 597.035 ;
        RECT 5.330 594.325 24.060 594.375 ;
        RECT 5.330 591.595 1094.530 594.325 ;
        RECT 5.330 591.545 281.595 591.595 ;
        RECT 5.330 588.885 432.540 588.935 ;
        RECT 5.330 586.155 1094.530 588.885 ;
        RECT 5.330 586.105 25.440 586.155 ;
        RECT 5.330 583.445 32.275 583.495 ;
        RECT 5.330 580.715 1094.530 583.445 ;
        RECT 5.330 580.665 156.475 580.715 ;
        RECT 5.330 578.005 46.535 578.055 ;
        RECT 5.330 575.275 1094.530 578.005 ;
        RECT 5.330 575.225 143.135 575.275 ;
        RECT 5.330 572.565 75.975 572.615 ;
        RECT 5.330 569.835 1094.530 572.565 ;
        RECT 5.330 569.785 129.335 569.835 ;
        RECT 5.330 567.125 299.535 567.175 ;
        RECT 5.330 564.395 1094.530 567.125 ;
        RECT 5.330 564.345 21.300 564.395 ;
        RECT 5.330 561.685 265.495 561.735 ;
        RECT 5.330 558.955 1094.530 561.685 ;
        RECT 5.330 558.905 90.695 558.955 ;
        RECT 5.330 556.245 76.435 556.295 ;
        RECT 5.330 553.515 1094.530 556.245 ;
        RECT 5.330 553.465 45.680 553.515 ;
        RECT 5.330 550.805 136.695 550.855 ;
        RECT 5.330 548.075 1094.530 550.805 ;
        RECT 5.330 548.025 26.295 548.075 ;
        RECT 5.330 545.365 27.740 545.415 ;
        RECT 5.330 542.635 1094.530 545.365 ;
        RECT 5.330 542.585 433.920 542.635 ;
        RECT 5.330 539.925 432.540 539.975 ;
        RECT 5.330 537.195 1094.530 539.925 ;
        RECT 5.330 537.145 93.520 537.195 ;
        RECT 5.330 534.485 37.400 534.535 ;
        RECT 5.330 531.755 1094.530 534.485 ;
        RECT 5.330 531.705 19.460 531.755 ;
        RECT 5.330 529.045 117.375 529.095 ;
        RECT 5.330 526.315 1094.530 529.045 ;
        RECT 5.330 526.265 653.735 526.315 ;
        RECT 5.330 523.605 184.995 523.655 ;
        RECT 5.330 520.875 1094.530 523.605 ;
        RECT 5.330 520.825 193.340 520.875 ;
        RECT 5.330 518.165 190.055 518.215 ;
        RECT 5.330 515.435 1094.530 518.165 ;
        RECT 5.330 515.385 429.255 515.435 ;
        RECT 5.330 512.725 191.040 512.775 ;
        RECT 5.330 509.995 1094.530 512.725 ;
        RECT 5.330 509.945 429.780 509.995 ;
        RECT 5.330 507.285 245.780 507.335 ;
        RECT 5.330 504.555 1094.530 507.285 ;
        RECT 5.330 504.505 444.435 504.555 ;
        RECT 5.330 501.845 317.935 501.895 ;
        RECT 5.330 499.115 1094.530 501.845 ;
        RECT 5.330 499.065 242.955 499.115 ;
        RECT 5.330 496.405 189.660 496.455 ;
        RECT 5.330 493.675 1094.530 496.405 ;
        RECT 5.330 493.625 183.615 493.675 ;
        RECT 5.330 490.965 431.620 491.015 ;
        RECT 5.330 488.235 1094.530 490.965 ;
        RECT 5.330 488.185 429.780 488.235 ;
        RECT 5.330 485.525 511.135 485.575 ;
        RECT 5.330 482.795 1094.530 485.525 ;
        RECT 5.330 482.745 615.095 482.795 ;
        RECT 5.330 480.085 62.635 480.135 ;
        RECT 5.330 477.355 1094.530 480.085 ;
        RECT 5.330 477.305 21.760 477.355 ;
        RECT 5.330 474.645 23.535 474.695 ;
        RECT 5.330 471.915 1094.530 474.645 ;
        RECT 5.330 471.865 69.535 471.915 ;
        RECT 5.330 469.205 23.140 469.255 ;
        RECT 5.330 466.475 1094.530 469.205 ;
        RECT 5.330 466.425 600.900 466.475 ;
        RECT 5.330 463.765 239.340 463.815 ;
        RECT 5.330 461.035 1094.530 463.765 ;
        RECT 5.330 460.985 52.055 461.035 ;
        RECT 5.330 458.325 106.795 458.375 ;
        RECT 5.330 455.595 1094.530 458.325 ;
        RECT 5.330 455.545 21.300 455.595 ;
        RECT 5.330 452.885 53.895 452.935 ;
        RECT 5.330 450.155 1094.530 452.885 ;
        RECT 5.330 450.105 73.215 450.155 ;
        RECT 5.330 447.445 56.720 447.495 ;
        RECT 5.330 444.715 1094.530 447.445 ;
        RECT 5.330 444.665 91.220 444.715 ;
        RECT 5.330 442.005 23.140 442.055 ;
        RECT 5.330 439.275 1094.530 442.005 ;
        RECT 5.330 439.225 134.000 439.275 ;
        RECT 5.330 436.565 241.180 436.615 ;
        RECT 5.330 433.835 1094.530 436.565 ;
        RECT 5.330 433.785 69.535 433.835 ;
        RECT 5.330 431.125 23.600 431.175 ;
        RECT 5.330 428.395 1094.530 431.125 ;
        RECT 5.330 428.345 53.500 428.395 ;
        RECT 5.330 425.685 141.295 425.735 ;
        RECT 5.330 422.955 1094.530 425.685 ;
        RECT 5.330 422.905 36.020 422.955 ;
        RECT 5.330 420.245 52.975 420.295 ;
        RECT 5.330 417.515 1094.530 420.245 ;
        RECT 5.330 417.465 376.880 417.515 ;
        RECT 5.330 414.805 469.735 414.855 ;
        RECT 5.330 412.075 1094.530 414.805 ;
        RECT 5.330 412.025 28.200 412.075 ;
        RECT 5.330 409.365 84.715 409.415 ;
        RECT 5.330 406.635 1094.530 409.365 ;
        RECT 5.330 406.585 26.295 406.635 ;
        RECT 5.330 403.925 144.515 403.975 ;
        RECT 5.330 401.195 1094.530 403.925 ;
        RECT 5.330 401.145 53.500 401.195 ;
        RECT 5.330 398.485 55.340 398.535 ;
        RECT 5.330 395.755 1094.530 398.485 ;
        RECT 5.330 395.705 23.140 395.755 ;
        RECT 5.330 393.045 117.835 393.095 ;
        RECT 5.330 390.315 1094.530 393.045 ;
        RECT 5.330 390.265 489.975 390.315 ;
        RECT 5.330 387.605 401.260 387.655 ;
        RECT 5.330 384.875 1094.530 387.605 ;
        RECT 5.330 384.825 134.000 384.875 ;
        RECT 5.330 382.165 54.355 382.215 ;
        RECT 5.330 379.435 1094.530 382.165 ;
        RECT 5.330 379.385 92.535 379.435 ;
        RECT 5.330 376.725 98.975 376.775 ;
        RECT 5.330 373.995 1094.530 376.725 ;
        RECT 5.330 373.945 21.300 373.995 ;
        RECT 5.330 371.285 72.755 371.335 ;
        RECT 5.330 368.555 1094.530 371.285 ;
        RECT 5.330 368.505 24.980 368.555 ;
        RECT 5.330 365.845 25.440 365.895 ;
        RECT 5.330 363.115 1094.530 365.845 ;
        RECT 5.330 363.065 55.340 363.115 ;
        RECT 5.330 360.405 102.655 360.455 ;
        RECT 5.330 357.675 1094.530 360.405 ;
        RECT 5.330 357.625 20.840 357.675 ;
        RECT 5.330 354.965 84.715 355.015 ;
        RECT 5.330 352.235 1094.530 354.965 ;
        RECT 5.330 352.185 115.075 352.235 ;
        RECT 5.330 349.525 249.395 349.575 ;
        RECT 5.330 346.795 1094.530 349.525 ;
        RECT 5.330 346.745 201.620 346.795 ;
        RECT 5.330 344.085 56.720 344.135 ;
        RECT 5.330 341.355 1094.530 344.085 ;
        RECT 5.330 341.305 20.380 341.355 ;
        RECT 5.330 338.645 53.500 338.695 ;
        RECT 5.330 335.915 1094.530 338.645 ;
        RECT 5.330 335.865 953.720 335.915 ;
        RECT 5.330 333.205 371.820 333.255 ;
        RECT 5.330 330.475 1094.530 333.205 ;
        RECT 5.330 330.425 142.215 330.475 ;
        RECT 5.330 327.765 20.315 327.815 ;
        RECT 5.330 325.035 1094.530 327.765 ;
        RECT 5.330 324.985 21.300 325.035 ;
        RECT 5.330 322.325 143.595 322.375 ;
        RECT 5.330 319.595 1094.530 322.325 ;
        RECT 5.330 319.545 64.015 319.595 ;
        RECT 5.330 316.885 66.380 316.935 ;
        RECT 5.330 314.155 1094.530 316.885 ;
        RECT 5.330 314.105 21.235 314.155 ;
        RECT 5.330 311.445 199.780 311.495 ;
        RECT 5.330 308.715 1094.530 311.445 ;
        RECT 5.330 308.665 249.460 308.715 ;
        RECT 5.330 306.005 68.680 306.055 ;
        RECT 5.330 303.275 1094.530 306.005 ;
        RECT 5.330 303.225 21.760 303.275 ;
        RECT 5.330 300.565 65.460 300.615 ;
        RECT 5.330 297.835 1094.530 300.565 ;
        RECT 5.330 297.785 54.420 297.835 ;
        RECT 5.330 295.125 270.095 295.175 ;
        RECT 5.330 292.395 1094.530 295.125 ;
        RECT 5.330 292.345 201.160 292.395 ;
        RECT 5.330 289.685 63.620 289.735 ;
        RECT 5.330 286.955 1094.530 289.685 ;
        RECT 5.330 286.905 26.295 286.955 ;
        RECT 5.330 284.245 24.980 284.295 ;
        RECT 5.330 281.515 1094.530 284.245 ;
        RECT 5.330 281.465 66.775 281.515 ;
        RECT 5.330 278.805 244.795 278.855 ;
        RECT 5.330 276.075 1094.530 278.805 ;
        RECT 5.330 276.025 131.175 276.075 ;
        RECT 5.330 273.365 145.500 273.415 ;
        RECT 5.330 270.635 1094.530 273.365 ;
        RECT 5.330 270.585 29.120 270.635 ;
        RECT 5.330 267.925 232.900 267.975 ;
        RECT 5.330 265.195 1094.530 267.925 ;
        RECT 5.330 265.145 34.575 265.195 ;
        RECT 5.330 262.485 92.075 262.535 ;
        RECT 5.330 259.755 1094.530 262.485 ;
        RECT 5.330 259.705 18.935 259.755 ;
        RECT 5.330 254.315 1094.530 257.095 ;
        RECT 5.330 254.265 19.920 254.315 ;
        RECT 5.330 251.605 39.635 251.655 ;
        RECT 5.330 248.875 1094.530 251.605 ;
        RECT 5.330 248.825 286.195 248.875 ;
        RECT 5.330 246.165 252.220 246.215 ;
        RECT 5.330 243.435 1094.530 246.165 ;
        RECT 5.330 243.385 202.015 243.435 ;
        RECT 5.330 240.725 206.680 240.775 ;
        RECT 5.330 237.995 1094.530 240.725 ;
        RECT 5.330 237.945 269.635 237.995 ;
        RECT 5.330 235.285 534.660 235.335 ;
        RECT 5.330 232.555 1094.530 235.285 ;
        RECT 5.330 232.505 954.180 232.555 ;
        RECT 5.330 229.845 199.780 229.895 ;
        RECT 5.330 227.115 1094.530 229.845 ;
        RECT 5.330 227.065 258.660 227.115 ;
        RECT 5.330 224.405 197.940 224.455 ;
        RECT 5.330 221.675 1094.530 224.405 ;
        RECT 5.330 221.625 234.215 221.675 ;
        RECT 5.330 218.965 335.875 219.015 ;
        RECT 5.330 216.235 1094.530 218.965 ;
        RECT 5.330 216.185 40.160 216.235 ;
        RECT 5.330 213.525 68.680 213.575 ;
        RECT 5.330 210.795 1094.530 213.525 ;
        RECT 5.330 210.745 38.255 210.795 ;
        RECT 5.330 208.085 41.080 208.135 ;
        RECT 5.330 205.355 1094.530 208.085 ;
        RECT 5.330 205.305 116.455 205.355 ;
        RECT 5.330 202.645 41.080 202.695 ;
        RECT 5.330 199.915 1094.530 202.645 ;
        RECT 5.330 199.865 210.360 199.915 ;
        RECT 5.330 197.205 65.855 197.255 ;
        RECT 5.330 194.475 1094.530 197.205 ;
        RECT 5.330 194.425 40.160 194.475 ;
        RECT 5.330 191.765 39.175 191.815 ;
        RECT 5.330 189.035 1094.530 191.765 ;
        RECT 5.330 188.985 37.860 189.035 ;
        RECT 5.330 186.325 39.635 186.375 ;
        RECT 5.330 183.595 1094.530 186.325 ;
        RECT 5.330 183.545 405.860 183.595 ;
        RECT 5.330 180.885 40.620 180.935 ;
        RECT 5.330 178.155 1094.530 180.885 ;
        RECT 5.330 178.105 138.075 178.155 ;
        RECT 5.330 175.445 207.600 175.495 ;
        RECT 5.330 172.715 1094.530 175.445 ;
        RECT 5.330 172.665 261.880 172.715 ;
        RECT 5.330 170.005 249.395 170.055 ;
        RECT 5.330 167.275 1094.530 170.005 ;
        RECT 5.330 167.225 388.840 167.275 ;
        RECT 5.330 164.565 964.235 164.615 ;
        RECT 5.330 161.835 1094.530 164.565 ;
        RECT 5.330 161.785 304.595 161.835 ;
        RECT 5.330 159.125 215.880 159.175 ;
        RECT 5.330 156.395 1094.530 159.125 ;
        RECT 5.330 156.345 206.155 156.395 ;
        RECT 5.330 153.685 285.735 153.735 ;
        RECT 5.330 150.955 1094.530 153.685 ;
        RECT 5.330 150.905 41.540 150.955 ;
        RECT 5.330 148.245 39.240 148.295 ;
        RECT 5.330 145.515 1094.530 148.245 ;
        RECT 5.330 145.465 104.955 145.515 ;
        RECT 5.330 142.805 37.335 142.855 ;
        RECT 5.330 140.075 1094.530 142.805 ;
        RECT 5.330 140.025 36.875 140.075 ;
        RECT 5.330 137.365 63.555 137.415 ;
        RECT 5.330 134.635 1094.530 137.365 ;
        RECT 5.330 134.585 37.860 134.635 ;
        RECT 5.330 131.925 38.780 131.975 ;
        RECT 5.330 129.195 1094.530 131.925 ;
        RECT 5.330 129.145 37.860 129.195 ;
        RECT 5.330 126.485 125.195 126.535 ;
        RECT 5.330 123.755 1094.530 126.485 ;
        RECT 5.330 123.705 37.860 123.755 ;
        RECT 5.330 121.045 39.175 121.095 ;
        RECT 5.330 118.315 1094.530 121.045 ;
        RECT 5.330 118.265 37.860 118.315 ;
        RECT 5.330 115.605 41.540 115.655 ;
        RECT 5.330 112.875 1094.530 115.605 ;
        RECT 5.330 112.825 60.795 112.875 ;
        RECT 5.330 110.165 324.375 110.215 ;
        RECT 5.330 107.435 1094.530 110.165 ;
        RECT 5.330 107.385 517.180 107.435 ;
        RECT 5.330 104.725 585.655 104.775 ;
        RECT 5.330 101.995 1094.530 104.725 ;
        RECT 5.330 101.945 275.680 101.995 ;
        RECT 5.330 99.285 423.735 99.335 ;
        RECT 5.330 96.555 1094.530 99.285 ;
        RECT 5.330 96.505 120.135 96.555 ;
        RECT 5.330 93.845 143.660 93.895 ;
        RECT 5.330 91.115 1094.530 93.845 ;
        RECT 5.330 91.065 308.800 91.115 ;
        RECT 5.330 88.405 74.135 88.455 ;
        RECT 5.330 85.675 1094.530 88.405 ;
        RECT 5.330 85.625 36.415 85.675 ;
        RECT 5.330 82.965 39.700 83.015 ;
        RECT 5.330 80.235 1094.530 82.965 ;
        RECT 5.330 80.185 52.515 80.235 ;
        RECT 5.330 77.525 40.160 77.575 ;
        RECT 5.330 74.795 1094.530 77.525 ;
        RECT 5.330 74.745 71.375 74.795 ;
        RECT 5.330 72.085 37.795 72.135 ;
        RECT 5.330 69.355 1094.530 72.085 ;
        RECT 5.330 69.305 39.240 69.355 ;
        RECT 5.330 66.645 54.355 66.695 ;
        RECT 5.330 63.915 1094.530 66.645 ;
        RECT 5.330 63.865 74.135 63.915 ;
        RECT 5.330 61.205 40.160 61.255 ;
        RECT 5.330 58.475 1094.530 61.205 ;
        RECT 5.330 58.425 52.515 58.475 ;
        RECT 5.330 55.765 39.240 55.815 ;
        RECT 5.330 53.035 1094.530 55.765 ;
        RECT 5.330 52.985 199.715 53.035 ;
        RECT 5.330 50.325 36.875 50.375 ;
        RECT 5.330 47.595 1094.530 50.325 ;
        RECT 5.330 47.545 103.575 47.595 ;
        RECT 5.330 44.885 112.380 44.935 ;
        RECT 5.330 42.155 1094.530 44.885 ;
        RECT 5.330 42.105 38.320 42.155 ;
        RECT 5.330 39.445 36.940 39.495 ;
        RECT 5.330 36.715 1094.530 39.445 ;
        RECT 5.330 36.665 39.175 36.715 ;
        RECT 5.330 34.005 40.160 34.055 ;
        RECT 5.330 31.275 1094.530 34.005 ;
        RECT 5.330 31.225 79.720 31.275 ;
        RECT 5.330 28.565 828.600 28.615 ;
        RECT 5.330 25.835 1094.530 28.565 ;
        RECT 5.330 25.785 903.055 25.835 ;
        RECT 5.330 20.345 1094.530 23.175 ;
        RECT 5.330 14.905 1094.530 17.735 ;
        RECT 5.330 10.690 1094.530 12.295 ;
      LAYER li1 ;
        RECT 5.520 10.795 1095.115 1387.285 ;
      LAYER met1 ;
        RECT 5.520 8.540 1095.175 1387.840 ;
      LAYER met2 ;
        RECT 7.090 1395.720 19.590 1396.000 ;
        RECT 20.430 1395.720 33.390 1396.000 ;
        RECT 34.230 1395.720 47.190 1396.000 ;
        RECT 48.030 1395.720 60.990 1396.000 ;
        RECT 61.830 1395.720 74.790 1396.000 ;
        RECT 75.630 1395.720 88.590 1396.000 ;
        RECT 89.430 1395.720 102.390 1396.000 ;
        RECT 103.230 1395.720 116.190 1396.000 ;
        RECT 117.030 1395.720 129.530 1396.000 ;
        RECT 130.370 1395.720 143.330 1396.000 ;
        RECT 144.170 1395.720 157.130 1396.000 ;
        RECT 157.970 1395.720 170.930 1396.000 ;
        RECT 171.770 1395.720 184.730 1396.000 ;
        RECT 185.570 1395.720 198.530 1396.000 ;
        RECT 199.370 1395.720 212.330 1396.000 ;
        RECT 213.170 1395.720 226.130 1396.000 ;
        RECT 226.970 1395.720 239.930 1396.000 ;
        RECT 240.770 1395.720 253.270 1396.000 ;
        RECT 254.110 1395.720 267.070 1396.000 ;
        RECT 267.910 1395.720 280.870 1396.000 ;
        RECT 281.710 1395.720 294.670 1396.000 ;
        RECT 295.510 1395.720 308.470 1396.000 ;
        RECT 309.310 1395.720 322.270 1396.000 ;
        RECT 323.110 1395.720 336.070 1396.000 ;
        RECT 336.910 1395.720 349.870 1396.000 ;
        RECT 350.710 1395.720 363.670 1396.000 ;
        RECT 364.510 1395.720 377.010 1396.000 ;
        RECT 377.850 1395.720 390.810 1396.000 ;
        RECT 391.650 1395.720 404.610 1396.000 ;
        RECT 405.450 1395.720 418.410 1396.000 ;
        RECT 419.250 1395.720 432.210 1396.000 ;
        RECT 433.050 1395.720 446.010 1396.000 ;
        RECT 446.850 1395.720 459.810 1396.000 ;
        RECT 460.650 1395.720 473.610 1396.000 ;
        RECT 474.450 1395.720 487.410 1396.000 ;
        RECT 488.250 1395.720 500.750 1396.000 ;
        RECT 501.590 1395.720 514.550 1396.000 ;
        RECT 515.390 1395.720 528.350 1396.000 ;
        RECT 529.190 1395.720 542.150 1396.000 ;
        RECT 542.990 1395.720 555.950 1396.000 ;
        RECT 556.790 1395.720 569.750 1396.000 ;
        RECT 570.590 1395.720 583.550 1396.000 ;
        RECT 584.390 1395.720 597.350 1396.000 ;
        RECT 598.190 1395.720 611.150 1396.000 ;
        RECT 611.990 1395.720 624.490 1396.000 ;
        RECT 625.330 1395.720 638.290 1396.000 ;
        RECT 639.130 1395.720 652.090 1396.000 ;
        RECT 652.930 1395.720 665.890 1396.000 ;
        RECT 666.730 1395.720 679.690 1396.000 ;
        RECT 680.530 1395.720 693.490 1396.000 ;
        RECT 694.330 1395.720 707.290 1396.000 ;
        RECT 708.130 1395.720 721.090 1396.000 ;
        RECT 721.930 1395.720 734.890 1396.000 ;
        RECT 735.730 1395.720 748.230 1396.000 ;
        RECT 749.070 1395.720 762.030 1396.000 ;
        RECT 762.870 1395.720 775.830 1396.000 ;
        RECT 776.670 1395.720 789.630 1396.000 ;
        RECT 790.470 1395.720 803.430 1396.000 ;
        RECT 804.270 1395.720 817.230 1396.000 ;
        RECT 818.070 1395.720 831.030 1396.000 ;
        RECT 831.870 1395.720 844.830 1396.000 ;
        RECT 845.670 1395.720 858.630 1396.000 ;
        RECT 859.470 1395.720 871.970 1396.000 ;
        RECT 872.810 1395.720 885.770 1396.000 ;
        RECT 886.610 1395.720 899.570 1396.000 ;
        RECT 900.410 1395.720 913.370 1396.000 ;
        RECT 914.210 1395.720 927.170 1396.000 ;
        RECT 928.010 1395.720 940.970 1396.000 ;
        RECT 941.810 1395.720 954.770 1396.000 ;
        RECT 955.610 1395.720 968.570 1396.000 ;
        RECT 969.410 1395.720 982.370 1396.000 ;
        RECT 983.210 1395.720 995.710 1396.000 ;
        RECT 996.550 1395.720 1009.510 1396.000 ;
        RECT 1010.350 1395.720 1023.310 1396.000 ;
        RECT 1024.150 1395.720 1037.110 1396.000 ;
        RECT 1037.950 1395.720 1050.910 1396.000 ;
        RECT 1051.750 1395.720 1064.710 1396.000 ;
        RECT 1065.550 1395.720 1078.510 1396.000 ;
        RECT 1079.350 1395.720 1092.310 1396.000 ;
        RECT 1093.150 1395.720 1094.240 1396.000 ;
        RECT 6.540 8.510 1094.240 1395.720 ;
      LAYER met3 ;
        RECT 8.805 10.715 1093.815 1387.365 ;
      LAYER met4 ;
        RECT 47.215 19.895 97.440 1385.665 ;
        RECT 99.840 19.895 174.240 1385.665 ;
        RECT 176.640 19.895 251.040 1385.665 ;
        RECT 253.440 19.895 327.840 1385.665 ;
        RECT 330.240 19.895 404.640 1385.665 ;
        RECT 407.040 19.895 481.440 1385.665 ;
        RECT 483.840 19.895 558.240 1385.665 ;
        RECT 560.640 19.895 635.040 1385.665 ;
        RECT 637.440 19.895 711.840 1385.665 ;
        RECT 714.240 19.895 788.640 1385.665 ;
        RECT 791.040 19.895 865.440 1385.665 ;
        RECT 867.840 19.895 942.240 1385.665 ;
        RECT 944.640 19.895 1019.040 1385.665 ;
        RECT 1021.440 19.895 1089.905 1385.665 ;
  END
END DFFRAM_1Kx32
END LIBRARY

