magic
tech sky130A
magscale 1 2
timestamp 1621698203
<< nwell >>
rect 1066 277157 218906 277478
rect 1066 276069 218906 276635
rect 1066 274981 218906 275547
rect 1066 273903 218906 274459
rect 1066 273893 86048 273903
rect 1066 273361 22371 273371
rect 1066 272815 218906 273361
rect 1066 272805 13552 272815
rect 1066 272273 16759 272283
rect 1066 271727 218906 272273
rect 1066 271717 14564 271727
rect 1066 271185 25407 271195
rect 1066 270639 218906 271185
rect 1066 270629 40587 270639
rect 1066 270097 123111 270107
rect 1066 269551 218906 270097
rect 1066 269541 22371 269551
rect 1066 269009 60840 269019
rect 1066 268463 218906 269009
rect 1066 268453 52087 268463
rect 1066 267921 7848 267931
rect 1066 267375 218906 267921
rect 1066 267365 14196 267375
rect 1066 266833 6652 266843
rect 1066 266287 218906 266833
rect 1066 266277 8571 266287
rect 1066 265745 6376 265755
rect 1066 265199 218906 265745
rect 1066 265189 15747 265199
rect 1066 264657 5811 264667
rect 1066 264111 218906 264657
rect 1066 264101 25591 264111
rect 1066 263569 6192 263579
rect 1066 263023 218906 263569
rect 1066 263013 52192 263023
rect 1066 262481 30375 262491
rect 1066 261935 218906 262481
rect 1066 261925 36723 261935
rect 1066 261393 5903 261403
rect 1066 260847 218906 261393
rect 1066 260837 14275 260847
rect 1066 260305 15103 260315
rect 1066 259759 218906 260305
rect 1066 259749 25315 259759
rect 1066 259217 109876 259227
rect 1066 258671 218906 259217
rect 1066 258661 56687 258671
rect 1066 258129 53375 258139
rect 1066 257583 218906 258129
rect 1066 257573 40127 257583
rect 1066 257041 6560 257051
rect 1066 256495 218906 257041
rect 1066 256485 7204 256495
rect 1066 255953 79227 255963
rect 1066 255407 218906 255953
rect 1066 255397 10411 255407
rect 1066 254865 6363 254875
rect 1066 254319 218906 254865
rect 1066 254309 36539 254319
rect 1066 253777 6836 253787
rect 1066 253231 218906 253777
rect 1066 253221 6731 253231
rect 1066 252689 31571 252699
rect 1066 252143 218906 252689
rect 1066 252133 7204 252143
rect 1066 251601 6455 251611
rect 1066 251055 218906 251601
rect 1066 251045 40035 251055
rect 1066 250513 6284 250523
rect 1066 249967 218906 250513
rect 1066 249957 11883 249967
rect 1066 249425 10135 249435
rect 1066 248879 218906 249425
rect 1066 248869 10056 248879
rect 1066 248337 5719 248347
rect 1066 247791 218906 248337
rect 1066 247781 5259 247791
rect 1066 247249 18336 247259
rect 1066 246703 218906 247249
rect 1066 246693 205004 246703
rect 1066 246161 13736 246171
rect 1066 245615 218906 246161
rect 1066 245605 31479 245615
rect 1066 245073 16207 245083
rect 1066 244527 218906 245073
rect 1066 244517 14288 244527
rect 1066 243985 25223 243995
rect 1066 243439 218906 243985
rect 1066 243429 13920 243439
rect 1066 242897 15116 242907
rect 1066 242351 218906 242897
rect 1066 242341 13815 242351
rect 1066 241809 63495 241819
rect 1066 241263 218906 241809
rect 1066 241253 14012 241263
rect 1066 240721 20360 240731
rect 1066 240175 218906 240721
rect 1066 240165 14380 240175
rect 1066 239633 63495 239643
rect 1066 239087 218906 239633
rect 1066 239077 29823 239087
rect 1066 238545 109692 238555
rect 1066 237999 218906 238545
rect 1066 237989 176484 237999
rect 1066 236911 218906 237467
rect 1066 236901 169768 236911
rect 1066 236369 56687 236379
rect 1066 235823 218906 236369
rect 1066 235813 170596 235823
rect 1066 235281 51824 235291
rect 1066 234735 218906 235281
rect 1066 234725 59999 234735
rect 1066 234193 51916 234203
rect 1066 233647 218906 234193
rect 1066 233637 86508 233647
rect 1066 233105 5640 233115
rect 1066 232559 218906 233105
rect 1066 232549 5456 232559
rect 1066 232017 8492 232027
rect 1066 231471 218906 232017
rect 1066 231461 11975 231471
rect 1066 230929 4628 230939
rect 1066 230383 218906 230929
rect 1066 230373 5088 230383
rect 1066 229841 11239 229851
rect 1066 229295 218906 229841
rect 1066 229285 31479 229295
rect 1066 228753 51824 228763
rect 1066 228207 218906 228753
rect 1066 228197 51995 228207
rect 1066 227665 100295 227675
rect 1066 227119 218906 227665
rect 1066 227109 118327 227119
rect 1066 226577 154115 226587
rect 1066 226031 218906 226577
rect 1066 226021 3511 226031
rect 1066 225489 33227 225499
rect 1066 224943 218906 225489
rect 1066 224933 59815 224943
rect 1066 224401 186223 224411
rect 1066 223855 218906 224401
rect 1066 223845 51548 223855
rect 1066 223313 48236 223323
rect 1066 222767 218906 223313
rect 1066 222757 67175 222767
rect 1066 222225 177115 222235
rect 1066 221679 218906 222225
rect 1066 221669 18875 221679
rect 1066 221137 6284 221147
rect 1066 220591 218906 221137
rect 1066 220581 11883 220591
rect 1066 220049 6468 220059
rect 1066 219503 218906 220049
rect 1066 219493 14564 219503
rect 1066 218961 5627 218971
rect 1066 218415 218906 218961
rect 1066 218405 31203 218415
rect 1066 217873 5811 217883
rect 1066 217327 218906 217873
rect 1066 217317 5824 217327
rect 1066 216785 30651 216795
rect 1066 216239 218906 216785
rect 1066 216229 50155 216239
rect 1066 215697 15300 215707
rect 1066 215151 218906 215697
rect 1066 215141 36723 215151
rect 1066 214609 4904 214619
rect 1066 214063 218906 214609
rect 1066 214053 22371 214063
rect 1066 213521 48959 213531
rect 1066 212975 218906 213521
rect 1066 212965 90543 212975
rect 1066 212433 30283 212443
rect 1066 211887 218906 212433
rect 1066 211877 29087 211887
rect 1066 211345 6100 211355
rect 1066 210799 218906 211345
rect 1066 210789 14196 210799
rect 1066 210257 7927 210267
rect 1066 209711 218906 210257
rect 1066 209701 8676 209711
rect 1066 209169 52008 209179
rect 1066 208623 218906 209169
rect 1066 208613 34515 208623
rect 1066 208081 37275 208091
rect 1066 207535 218906 208081
rect 1066 207525 64691 207535
rect 1066 206993 118616 207003
rect 1066 206447 218906 206993
rect 1066 206437 5088 206447
rect 1066 205905 6100 205915
rect 1066 205359 218906 205905
rect 1066 205349 5732 205359
rect 1066 204817 6376 204827
rect 1066 204271 218906 204817
rect 1066 204261 6915 204271
rect 1066 203729 9307 203739
rect 1066 203183 218906 203729
rect 1066 203173 14091 203183
rect 1066 202641 37183 202651
rect 1066 202095 218906 202641
rect 1066 202085 90543 202095
rect 1066 201553 89623 201563
rect 1066 201007 218906 201553
rect 1066 200997 4260 201007
rect 1066 200465 31939 200475
rect 1066 199919 218906 200465
rect 1066 199909 35527 199919
rect 1066 199377 16943 199387
rect 1066 198831 218906 199377
rect 1066 198821 5824 198831
rect 1066 198289 20163 198299
rect 1066 197743 218906 198289
rect 1066 197733 5088 197743
rect 1066 197201 17495 197211
rect 1066 196655 218906 197201
rect 1066 196645 14551 196655
rect 1066 196113 23672 196123
rect 1066 195567 218906 196113
rect 1066 195557 25867 195567
rect 1066 195025 4996 195035
rect 1066 194479 218906 195025
rect 1066 194469 9031 194479
rect 1066 193937 5627 193947
rect 1066 193391 218906 193937
rect 1066 193381 12159 193391
rect 1066 192849 31676 192859
rect 1066 192303 218906 192849
rect 1066 192293 32044 192303
rect 1066 191761 58619 191771
rect 1066 191215 218906 191761
rect 1066 191205 34896 191215
rect 1066 190673 63219 190683
rect 1066 190127 218906 190673
rect 1066 190117 31584 190127
rect 1066 189585 48788 189595
rect 1066 189039 218906 189585
rect 1066 189029 36723 189039
rect 1066 188497 32136 188507
rect 1066 187951 218906 188497
rect 1066 187941 55399 187951
rect 1066 187409 34252 187419
rect 1066 186863 218906 187409
rect 1066 186853 6639 186863
rect 1066 186321 4063 186331
rect 1066 185775 218906 186321
rect 1066 185765 8755 185775
rect 1066 185233 33503 185243
rect 1066 184687 218906 185233
rect 1066 184677 2144 184687
rect 1066 184145 7927 184155
rect 1066 183599 218906 184145
rect 1066 183589 8387 183599
rect 1066 183057 7927 183067
rect 1066 182511 218906 183057
rect 1066 182501 4352 182511
rect 1066 181969 1579 181979
rect 1066 181423 218906 181969
rect 1066 181413 8111 181423
rect 1066 180881 4523 180891
rect 1066 180335 218906 180881
rect 1066 180325 15747 180335
rect 1066 179793 7927 179803
rect 1066 179247 218906 179793
rect 1066 179237 15944 179247
rect 1066 178705 19887 178715
rect 1066 178159 218906 178705
rect 1066 178149 19887 178159
rect 1066 177617 7835 177627
rect 1066 177071 218906 177617
rect 1066 177061 41967 177071
rect 1066 176529 38300 176539
rect 1066 175983 218906 176529
rect 1066 175973 4260 175983
rect 1066 175441 48880 175451
rect 1066 174895 218906 175441
rect 1066 174885 7204 174895
rect 1066 174353 7927 174363
rect 1066 173807 218906 174353
rect 1066 173797 18047 173807
rect 1066 173265 11331 173275
rect 1066 172719 218906 173265
rect 1066 172709 18047 172719
rect 1066 172177 15011 172187
rect 1066 171631 218906 172177
rect 1066 171621 31952 171631
rect 1066 171089 5272 171099
rect 1066 170543 218906 171089
rect 1066 170533 8755 170543
rect 1066 170001 9872 170011
rect 1066 169455 218906 170001
rect 1066 169445 33595 169455
rect 1066 168913 62207 168923
rect 1066 168367 218906 168913
rect 1066 168357 17495 168367
rect 1066 167825 25880 167835
rect 1066 167279 218906 167825
rect 1066 167269 17127 167279
rect 1066 166737 39207 166747
rect 1066 166191 218906 166737
rect 1066 166181 8860 166191
rect 1066 165649 5364 165659
rect 1066 165103 218906 165649
rect 1066 165093 5824 165103
rect 1066 164561 6836 164571
rect 1066 164015 218906 164561
rect 1066 164005 7559 164015
rect 1066 163473 85864 163483
rect 1066 162927 218906 163473
rect 1066 162917 5259 162927
rect 1066 162385 103699 162395
rect 1066 161839 218906 162385
rect 1066 161829 2144 161839
rect 1066 161297 104527 161307
rect 1066 160751 218906 161297
rect 1066 160741 8387 160751
rect 1066 160209 30283 160219
rect 1066 159663 218906 160209
rect 1066 159653 3616 159663
rect 1066 159121 6455 159131
rect 1066 158575 218906 159121
rect 1066 158565 22371 158575
rect 1066 158033 18323 158043
rect 1066 157487 218906 158033
rect 1066 157477 1671 157487
rect 1066 156945 26787 156955
rect 1066 156399 218906 156945
rect 1066 156389 72603 156399
rect 1066 155857 155140 155867
rect 1066 155311 218906 155857
rect 1066 155301 14919 155311
rect 1066 154769 28903 154779
rect 1066 154223 218906 154769
rect 1066 154213 15300 154223
rect 1066 153681 9307 153691
rect 1066 153135 218906 153681
rect 1066 153125 2144 153135
rect 1066 152593 6271 152603
rect 1066 152047 218906 152593
rect 1066 152037 17692 152047
rect 1066 151505 2144 151515
rect 1066 150959 218906 151505
rect 1066 150949 94039 150959
rect 1066 150417 25775 150427
rect 1066 149871 218906 150417
rect 1066 149861 5259 149871
rect 1066 149329 60367 149339
rect 1066 148783 218906 149329
rect 1066 148773 21556 148783
rect 1066 148241 6100 148251
rect 1066 147695 218906 148241
rect 1066 147685 25696 147695
rect 1066 147153 26235 147163
rect 1066 146607 218906 147153
rect 1066 146597 26524 146607
rect 1066 146065 2144 146075
rect 1066 145519 218906 146065
rect 1066 145509 3787 145519
rect 1066 144977 15484 144987
rect 1066 144431 218906 144977
rect 1066 144421 1579 144431
rect 1066 143889 16772 143899
rect 1066 143343 218906 143889
rect 1066 143333 4628 143343
rect 1066 142801 2144 142811
rect 1066 142255 218906 142801
rect 1066 142245 60551 142255
rect 1066 141713 92304 141723
rect 1066 141167 218906 141713
rect 1066 141157 97903 141167
rect 1066 140625 6376 140635
rect 1066 140079 218906 140625
rect 1066 140069 49156 140079
rect 1066 139537 68187 139547
rect 1066 138991 218906 139537
rect 1066 138981 3616 138991
rect 1066 138449 48407 138459
rect 1066 137903 218906 138449
rect 1066 137893 54663 137903
rect 1066 137361 58908 137371
rect 1066 136815 218906 137361
rect 1066 136805 10503 136815
rect 1066 136273 50444 136283
rect 1066 135727 218906 136273
rect 1066 135717 54400 135727
rect 1066 135185 28903 135195
rect 1066 134639 218906 135185
rect 1066 134629 8847 134639
rect 1066 134097 5364 134107
rect 1066 133551 218906 134097
rect 1066 133541 4891 133551
rect 1066 133009 107563 133019
rect 1066 132463 218906 133009
rect 1066 132453 57988 132463
rect 1066 131921 114463 131931
rect 1066 131375 218906 131921
rect 1066 131365 24316 131375
rect 1066 130833 27155 130843
rect 1066 130287 218906 130833
rect 1066 130277 23488 130287
rect 1066 129745 37275 129755
rect 1066 129199 218906 129745
rect 1066 129189 24119 129199
rect 1066 128657 33963 128667
rect 1066 128111 218906 128657
rect 1066 128101 20084 128111
rect 1066 127569 25315 127579
rect 1066 127023 218906 127569
rect 1066 127013 20820 127023
rect 1066 126481 24040 126491
rect 1066 125935 218906 126481
rect 1066 125925 20636 125935
rect 1066 125393 52560 125403
rect 1066 124847 218906 125393
rect 1066 124837 28548 124847
rect 1066 124305 28167 124315
rect 1066 123759 218906 124305
rect 1066 123749 18967 123759
rect 1066 123217 20360 123227
rect 1066 122671 218906 123217
rect 1066 122661 76743 122671
rect 1066 122129 13171 122139
rect 1066 121583 218906 122129
rect 1066 121573 10135 121583
rect 1066 121041 9872 121051
rect 1066 120495 218906 121041
rect 1066 120485 10148 120495
rect 1066 119953 10332 119963
rect 1066 119407 218906 119953
rect 1066 119397 10227 119407
rect 1066 118865 10056 118875
rect 1066 118319 218906 118865
rect 1066 118309 13907 118319
rect 1066 117777 10056 117787
rect 1066 117231 218906 117777
rect 1066 117221 10240 117231
rect 1066 116689 10240 116699
rect 1066 116143 218906 116689
rect 1066 116133 10319 116143
rect 1066 115601 10148 115611
rect 1066 115055 218906 115601
rect 1066 115045 10411 115055
rect 1066 114513 26143 114523
rect 1066 113967 218906 114513
rect 1066 113957 32859 113967
rect 1066 113425 123295 113435
rect 1066 112879 218906 113425
rect 1066 112869 117328 112879
rect 1066 112337 119996 112347
rect 1066 111791 218906 112337
rect 1066 111781 19519 111791
rect 1066 111249 16404 111259
rect 1066 110703 218906 111249
rect 1066 110693 15576 110703
rect 1066 110161 15116 110171
rect 1066 109615 218906 110161
rect 1066 109605 27615 109615
rect 1066 109073 15208 109083
rect 1066 108527 218906 109073
rect 1066 108517 15747 108527
rect 1066 107985 48959 107995
rect 1066 107439 218906 107985
rect 1066 107429 28167 107439
rect 1066 106897 18415 106907
rect 1066 106351 218906 106897
rect 1066 106341 16036 106351
rect 1066 105809 23659 105819
rect 1066 105263 218906 105809
rect 1066 105253 16128 105263
rect 1066 104721 30927 104731
rect 1066 104175 218906 104721
rect 1066 104165 17692 104175
rect 1066 103633 15484 103643
rect 1066 103087 218906 103633
rect 1066 103077 25499 103087
rect 1066 102545 15392 102555
rect 1066 101999 218906 102545
rect 1066 101989 18599 101999
rect 1066 101457 49603 101467
rect 1066 100911 218906 101457
rect 1066 100901 91292 100911
rect 1066 100369 7480 100379
rect 1066 99823 218906 100369
rect 1066 99813 5272 99823
rect 1066 99281 31203 99291
rect 1066 98735 218906 99281
rect 1066 98725 73247 98735
rect 1066 98193 5548 98203
rect 1066 97647 218906 98193
rect 1066 97637 9780 97647
rect 1066 97105 16115 97115
rect 1066 96559 218906 97105
rect 1066 96549 7664 96559
rect 1066 96017 31111 96027
rect 1066 95471 218906 96017
rect 1066 95461 32859 95471
rect 1066 94929 31571 94939
rect 1066 94383 218906 94929
rect 1066 94373 18599 94383
rect 1066 93841 15116 93851
rect 1066 93295 218906 93841
rect 1066 93285 57804 93295
rect 1066 92753 32031 92763
rect 1066 92207 218906 92753
rect 1066 92197 29179 92207
rect 1066 91665 46856 91675
rect 1066 91119 218906 91665
rect 1066 91109 119707 91119
rect 1066 90577 23659 90587
rect 1066 90031 218906 90577
rect 1066 90021 49156 90031
rect 1066 89489 58632 89499
rect 1066 88943 218906 89489
rect 1066 88933 4431 88943
rect 1066 88401 9872 88411
rect 1066 87855 218906 88401
rect 1066 87845 4260 87855
rect 1066 87313 4904 87323
rect 1066 86767 218906 87313
rect 1066 86757 70027 86767
rect 1066 86225 84760 86235
rect 1066 85679 218906 86225
rect 1066 85669 4996 85679
rect 1066 85137 4339 85147
rect 1066 84591 218906 85137
rect 1066 84581 101491 84591
rect 1066 84049 45200 84059
rect 1066 83503 218906 84049
rect 1066 83493 54400 83503
rect 1066 82961 7756 82971
rect 1066 82415 218906 82961
rect 1066 82405 5364 82415
rect 1066 81873 44635 81883
rect 1066 81327 218906 81873
rect 1066 81317 53835 81327
rect 1066 80785 6744 80795
rect 1066 80239 218906 80785
rect 1066 80229 45844 80239
rect 1066 79697 24040 79707
rect 1066 79151 218906 79697
rect 1066 79141 28811 79151
rect 1066 78609 14827 78619
rect 1066 78063 218906 78609
rect 1066 78053 9951 78063
rect 1066 77521 31755 77531
rect 1066 76975 218906 77521
rect 1066 76965 4812 76975
rect 1066 76433 49892 76443
rect 1066 75887 218906 76433
rect 1066 75877 5732 75887
rect 1066 75345 22003 75355
rect 1066 74799 218906 75345
rect 1066 74789 5364 74799
rect 1066 74257 7927 74267
rect 1066 73711 218906 74257
rect 1066 73701 34515 73711
rect 1066 73169 56503 73179
rect 1066 72623 218906 73169
rect 1066 72613 30835 72623
rect 1066 72081 7664 72091
rect 1066 71535 218906 72081
rect 1066 71525 31479 71535
rect 1066 70993 15379 71003
rect 1066 70447 218906 70993
rect 1066 70437 7848 70447
rect 1066 69905 7927 69915
rect 1066 69359 218906 69905
rect 1066 69349 24947 69359
rect 1066 68817 24224 68827
rect 1066 68271 218906 68817
rect 1066 68261 17495 68271
rect 1066 67729 17127 67739
rect 1066 67183 218906 67729
rect 1066 67173 2144 67183
rect 1066 66641 10227 66651
rect 1066 66095 218906 66641
rect 1066 66085 31479 66095
rect 1066 65553 97075 65563
rect 1066 65007 218906 65553
rect 1066 64997 10135 65007
rect 1066 64465 65519 64475
rect 1066 63919 218906 64465
rect 1066 63909 83380 63919
rect 1066 63377 10043 63387
rect 1066 62831 218906 63377
rect 1066 62821 2144 62831
rect 1066 62289 4812 62299
rect 1066 61743 218906 62289
rect 1066 61733 15747 61743
rect 1066 61201 16023 61211
rect 1066 60655 218906 61201
rect 1066 60645 6915 60655
rect 1066 60113 10043 60123
rect 1066 59557 218906 60113
rect 1066 59025 83472 59035
rect 1066 58479 218906 59025
rect 1066 58469 5272 58479
rect 1066 57937 9859 57947
rect 1066 57391 218906 57937
rect 1066 57381 1579 57391
rect 1066 56849 98455 56859
rect 1066 56303 218906 56849
rect 1066 56293 6731 56303
rect 1066 55761 55123 55771
rect 1066 55215 218906 55761
rect 1066 55205 53835 55215
rect 1066 54673 49327 54683
rect 1066 54127 218906 54673
rect 1066 54117 4247 54127
rect 1066 53585 23015 53595
rect 1066 53039 218906 53585
rect 1066 53029 15287 53039
rect 1066 52497 25039 52507
rect 1066 51951 218906 52497
rect 1066 51941 3800 51951
rect 1066 51409 11331 51419
rect 1066 50863 218906 51409
rect 1066 50853 4076 50863
rect 1066 50321 7467 50331
rect 1066 49775 218906 50321
rect 1066 49765 3695 49775
rect 1066 49233 14643 49243
rect 1066 48687 218906 49233
rect 1066 48677 8479 48687
rect 1066 48145 29468 48155
rect 1066 47599 218906 48145
rect 1066 47589 13999 47599
rect 1066 47057 58067 47067
rect 1066 46511 218906 47057
rect 1066 46501 54492 46511
rect 1066 45969 29284 45979
rect 1066 45423 218906 45969
rect 1066 45413 38103 45423
rect 1066 44881 83288 44891
rect 1066 44335 218906 44881
rect 1066 44325 8847 44335
rect 1066 43793 49064 43803
rect 1066 43247 218906 43793
rect 1066 43237 29284 43247
rect 1066 42705 68647 42715
rect 1066 42159 218906 42705
rect 1066 42149 47592 42159
rect 1066 41617 29376 41627
rect 1066 41071 218906 41617
rect 1066 41061 2144 41071
rect 1066 40529 68463 40539
rect 1066 39983 218906 40529
rect 1066 39973 5548 39983
rect 1066 39441 11515 39451
rect 1066 38895 218906 39441
rect 1066 38885 4628 38895
rect 1066 38353 4628 38363
rect 1066 37807 218906 38353
rect 1066 37797 7480 37807
rect 1066 37265 23120 37275
rect 1066 36719 218906 37265
rect 1066 36709 59539 36719
rect 1066 36177 35711 36187
rect 1066 35631 218906 36177
rect 1066 35621 125884 35631
rect 1066 35089 9307 35099
rect 1066 34543 218906 35089
rect 1066 34533 14643 34543
rect 1066 34001 27155 34011
rect 1066 33455 218906 34001
rect 1066 33445 23212 33455
rect 1066 32913 23488 32923
rect 1066 32367 218906 32913
rect 1066 32357 35711 32367
rect 1066 31825 55031 31835
rect 1066 31279 218906 31825
rect 1066 31269 48591 31279
rect 1066 30737 48236 30747
rect 1066 30191 218906 30737
rect 1066 30181 3984 30191
rect 1066 29649 9872 29659
rect 1066 29103 218906 29649
rect 1066 29093 76940 29103
rect 1066 28561 163683 28571
rect 1066 28015 218906 28561
rect 1066 28005 3892 28015
rect 1066 27473 7572 27483
rect 1066 26927 218906 27473
rect 1066 26917 10043 26927
rect 1066 26385 16391 26395
rect 1066 25839 218906 26385
rect 1066 25829 26064 25839
rect 1066 25297 27444 25307
rect 1066 24751 218906 25297
rect 1066 24741 14091 24751
rect 1066 24209 27155 24219
rect 1066 23663 218906 24209
rect 1066 23653 7204 23663
rect 1066 23121 45200 23131
rect 1066 22575 218906 23121
rect 1066 22565 4352 22575
rect 1066 22033 52652 22043
rect 1066 21487 218906 22033
rect 1066 21477 9504 21487
rect 1066 20945 7296 20955
rect 1066 20399 218906 20945
rect 1066 20389 14919 20399
rect 1066 19857 1579 19867
rect 1066 19311 218906 19857
rect 1066 19301 24040 19311
rect 1066 18769 4720 18779
rect 1066 18223 218906 18769
rect 1066 18213 4996 18223
rect 1066 17681 31295 17691
rect 1066 17135 218906 17681
rect 1066 17125 25052 17135
rect 1066 16593 23948 16603
rect 1066 16047 218906 16593
rect 1066 16037 88164 16047
rect 1066 15505 52363 15515
rect 1066 14959 218906 15505
rect 1066 14949 45936 14959
rect 1066 14417 13184 14427
rect 1066 13871 218906 14417
rect 1066 13861 4983 13871
rect 1066 13329 27812 13339
rect 1066 12783 218906 13329
rect 1066 12773 15471 12783
rect 1066 12241 4628 12251
rect 1066 11695 218906 12241
rect 1066 11685 7191 11695
rect 1066 11153 12895 11163
rect 1066 10607 218906 11153
rect 1066 10597 30007 10607
rect 1066 10065 24132 10075
rect 1066 9519 218906 10065
rect 1066 9509 27615 9519
rect 1066 8977 7467 8987
rect 1066 8431 218906 8977
rect 1066 8421 2144 8431
rect 1066 7889 9583 7899
rect 1066 7343 218906 7889
rect 1066 7333 7204 7343
rect 1066 6801 68831 6811
rect 1066 6255 218906 6801
rect 1066 6245 76651 6255
rect 1066 5713 92396 5723
rect 1066 5167 218906 5713
rect 1066 5157 129735 5167
rect 1066 4069 218906 4635
rect 1066 2981 218906 3547
rect 1066 2138 218906 2459
<< obsli1 >>
rect 1104 2159 219023 277457
<< obsm1 >>
rect 1104 1980 219035 277488
<< metal2 >>
rect 1306 279200 1362 280000
rect 3974 279200 4030 280000
rect 6734 279200 6790 280000
rect 9494 279200 9550 280000
rect 12254 279200 12310 280000
rect 15014 279200 15070 280000
rect 17774 279200 17830 280000
rect 20534 279200 20590 280000
rect 23294 279200 23350 280000
rect 25962 279200 26018 280000
rect 28722 279200 28778 280000
rect 31482 279200 31538 280000
rect 34242 279200 34298 280000
rect 37002 279200 37058 280000
rect 39762 279200 39818 280000
rect 42522 279200 42578 280000
rect 45282 279200 45338 280000
rect 48042 279200 48098 280000
rect 50710 279200 50766 280000
rect 53470 279200 53526 280000
rect 56230 279200 56286 280000
rect 58990 279200 59046 280000
rect 61750 279200 61806 280000
rect 64510 279200 64566 280000
rect 67270 279200 67326 280000
rect 70030 279200 70086 280000
rect 72790 279200 72846 280000
rect 75458 279200 75514 280000
rect 78218 279200 78274 280000
rect 80978 279200 81034 280000
rect 83738 279200 83794 280000
rect 86498 279200 86554 280000
rect 89258 279200 89314 280000
rect 92018 279200 92074 280000
rect 94778 279200 94834 280000
rect 97538 279200 97594 280000
rect 100206 279200 100262 280000
rect 102966 279200 103022 280000
rect 105726 279200 105782 280000
rect 108486 279200 108542 280000
rect 111246 279200 111302 280000
rect 114006 279200 114062 280000
rect 116766 279200 116822 280000
rect 119526 279200 119582 280000
rect 122286 279200 122342 280000
rect 124954 279200 125010 280000
rect 127714 279200 127770 280000
rect 130474 279200 130530 280000
rect 133234 279200 133290 280000
rect 135994 279200 136050 280000
rect 138754 279200 138810 280000
rect 141514 279200 141570 280000
rect 144274 279200 144330 280000
rect 147034 279200 147090 280000
rect 149702 279200 149758 280000
rect 152462 279200 152518 280000
rect 155222 279200 155278 280000
rect 157982 279200 158038 280000
rect 160742 279200 160798 280000
rect 163502 279200 163558 280000
rect 166262 279200 166318 280000
rect 169022 279200 169078 280000
rect 171782 279200 171838 280000
rect 174450 279200 174506 280000
rect 177210 279200 177266 280000
rect 179970 279200 180026 280000
rect 182730 279200 182786 280000
rect 185490 279200 185546 280000
rect 188250 279200 188306 280000
rect 191010 279200 191066 280000
rect 193770 279200 193826 280000
rect 196530 279200 196586 280000
rect 199198 279200 199254 280000
rect 201958 279200 202014 280000
rect 204718 279200 204774 280000
rect 207478 279200 207534 280000
rect 210238 279200 210294 280000
rect 212998 279200 213054 280000
rect 215758 279200 215814 280000
rect 218518 279200 218574 280000
<< obsm2 >>
rect 1418 279144 3918 279200
rect 4086 279144 6678 279200
rect 6846 279144 9438 279200
rect 9606 279144 12198 279200
rect 12366 279144 14958 279200
rect 15126 279144 17718 279200
rect 17886 279144 20478 279200
rect 20646 279144 23238 279200
rect 23406 279144 25906 279200
rect 26074 279144 28666 279200
rect 28834 279144 31426 279200
rect 31594 279144 34186 279200
rect 34354 279144 36946 279200
rect 37114 279144 39706 279200
rect 39874 279144 42466 279200
rect 42634 279144 45226 279200
rect 45394 279144 47986 279200
rect 48154 279144 50654 279200
rect 50822 279144 53414 279200
rect 53582 279144 56174 279200
rect 56342 279144 58934 279200
rect 59102 279144 61694 279200
rect 61862 279144 64454 279200
rect 64622 279144 67214 279200
rect 67382 279144 69974 279200
rect 70142 279144 72734 279200
rect 72902 279144 75402 279200
rect 75570 279144 78162 279200
rect 78330 279144 80922 279200
rect 81090 279144 83682 279200
rect 83850 279144 86442 279200
rect 86610 279144 89202 279200
rect 89370 279144 91962 279200
rect 92130 279144 94722 279200
rect 94890 279144 97482 279200
rect 97650 279144 100150 279200
rect 100318 279144 102910 279200
rect 103078 279144 105670 279200
rect 105838 279144 108430 279200
rect 108598 279144 111190 279200
rect 111358 279144 113950 279200
rect 114118 279144 116710 279200
rect 116878 279144 119470 279200
rect 119638 279144 122230 279200
rect 122398 279144 124898 279200
rect 125066 279144 127658 279200
rect 127826 279144 130418 279200
rect 130586 279144 133178 279200
rect 133346 279144 135938 279200
rect 136106 279144 138698 279200
rect 138866 279144 141458 279200
rect 141626 279144 144218 279200
rect 144386 279144 146978 279200
rect 147146 279144 149646 279200
rect 149814 279144 152406 279200
rect 152574 279144 155166 279200
rect 155334 279144 157926 279200
rect 158094 279144 160686 279200
rect 160854 279144 163446 279200
rect 163614 279144 166206 279200
rect 166374 279144 168966 279200
rect 169134 279144 171726 279200
rect 171894 279144 174394 279200
rect 174562 279144 177154 279200
rect 177322 279144 179914 279200
rect 180082 279144 182674 279200
rect 182842 279144 185434 279200
rect 185602 279144 188194 279200
rect 188362 279144 190954 279200
rect 191122 279144 193714 279200
rect 193882 279144 196474 279200
rect 196642 279144 199142 279200
rect 199310 279144 201902 279200
rect 202070 279144 204662 279200
rect 204830 279144 207422 279200
rect 207590 279144 210182 279200
rect 210350 279144 212942 279200
rect 213110 279144 215702 279200
rect 215870 279144 218462 279200
rect 218630 279144 218666 279200
rect 1306 1974 218666 279144
<< obsm3 >>
rect 1301 2143 218671 277473
<< metal4 >>
rect 4208 2128 4528 277488
rect 19568 2128 19888 277488
rect 34928 2128 35248 277488
rect 50288 2128 50608 277488
rect 65648 2128 65968 277488
rect 81008 2128 81328 277488
rect 96368 2128 96688 277488
rect 111728 2128 112048 277488
rect 127088 2128 127408 277488
rect 142448 2128 142768 277488
rect 157808 2128 158128 277488
rect 173168 2128 173488 277488
rect 188528 2128 188848 277488
rect 203888 2128 204208 277488
<< obsm4 >>
rect 2819 5339 4128 276181
rect 4608 5339 19488 276181
rect 19968 5339 34848 276181
rect 35328 5339 50208 276181
rect 50688 5339 65568 276181
rect 66048 5339 80928 276181
rect 81408 5339 96288 276181
rect 96768 5339 111648 276181
rect 112128 5339 127008 276181
rect 127488 5339 142368 276181
rect 142848 5339 157728 276181
rect 158208 5339 173088 276181
rect 173568 5339 188448 276181
rect 188928 5339 203808 276181
rect 204288 5339 212829 276181
<< labels >>
rlabel metal2 s 89258 279200 89314 280000 6 A[0]
port 1 nsew signal input
rlabel metal2 s 92018 279200 92074 280000 6 A[1]
port 2 nsew signal input
rlabel metal2 s 94778 279200 94834 280000 6 A[2]
port 3 nsew signal input
rlabel metal2 s 97538 279200 97594 280000 6 A[3]
port 4 nsew signal input
rlabel metal2 s 100206 279200 100262 280000 6 A[4]
port 5 nsew signal input
rlabel metal2 s 102966 279200 103022 280000 6 A[5]
port 6 nsew signal input
rlabel metal2 s 105726 279200 105782 280000 6 A[6]
port 7 nsew signal input
rlabel metal2 s 108486 279200 108542 280000 6 A[7]
port 8 nsew signal input
rlabel metal2 s 111246 279200 111302 280000 6 A[8]
port 9 nsew signal input
rlabel metal2 s 114006 279200 114062 280000 6 A[9]
port 10 nsew signal input
rlabel metal2 s 116766 279200 116822 280000 6 CLK
port 11 nsew signal input
rlabel metal2 s 133234 279200 133290 280000 6 Di[0]
port 12 nsew signal input
rlabel metal2 s 160742 279200 160798 280000 6 Di[10]
port 13 nsew signal input
rlabel metal2 s 163502 279200 163558 280000 6 Di[11]
port 14 nsew signal input
rlabel metal2 s 166262 279200 166318 280000 6 Di[12]
port 15 nsew signal input
rlabel metal2 s 169022 279200 169078 280000 6 Di[13]
port 16 nsew signal input
rlabel metal2 s 171782 279200 171838 280000 6 Di[14]
port 17 nsew signal input
rlabel metal2 s 174450 279200 174506 280000 6 Di[15]
port 18 nsew signal input
rlabel metal2 s 177210 279200 177266 280000 6 Di[16]
port 19 nsew signal input
rlabel metal2 s 179970 279200 180026 280000 6 Di[17]
port 20 nsew signal input
rlabel metal2 s 182730 279200 182786 280000 6 Di[18]
port 21 nsew signal input
rlabel metal2 s 185490 279200 185546 280000 6 Di[19]
port 22 nsew signal input
rlabel metal2 s 135994 279200 136050 280000 6 Di[1]
port 23 nsew signal input
rlabel metal2 s 188250 279200 188306 280000 6 Di[20]
port 24 nsew signal input
rlabel metal2 s 191010 279200 191066 280000 6 Di[21]
port 25 nsew signal input
rlabel metal2 s 193770 279200 193826 280000 6 Di[22]
port 26 nsew signal input
rlabel metal2 s 196530 279200 196586 280000 6 Di[23]
port 27 nsew signal input
rlabel metal2 s 199198 279200 199254 280000 6 Di[24]
port 28 nsew signal input
rlabel metal2 s 201958 279200 202014 280000 6 Di[25]
port 29 nsew signal input
rlabel metal2 s 204718 279200 204774 280000 6 Di[26]
port 30 nsew signal input
rlabel metal2 s 207478 279200 207534 280000 6 Di[27]
port 31 nsew signal input
rlabel metal2 s 210238 279200 210294 280000 6 Di[28]
port 32 nsew signal input
rlabel metal2 s 212998 279200 213054 280000 6 Di[29]
port 33 nsew signal input
rlabel metal2 s 138754 279200 138810 280000 6 Di[2]
port 34 nsew signal input
rlabel metal2 s 215758 279200 215814 280000 6 Di[30]
port 35 nsew signal input
rlabel metal2 s 218518 279200 218574 280000 6 Di[31]
port 36 nsew signal input
rlabel metal2 s 141514 279200 141570 280000 6 Di[3]
port 37 nsew signal input
rlabel metal2 s 144274 279200 144330 280000 6 Di[4]
port 38 nsew signal input
rlabel metal2 s 147034 279200 147090 280000 6 Di[5]
port 39 nsew signal input
rlabel metal2 s 149702 279200 149758 280000 6 Di[6]
port 40 nsew signal input
rlabel metal2 s 152462 279200 152518 280000 6 Di[7]
port 41 nsew signal input
rlabel metal2 s 155222 279200 155278 280000 6 Di[8]
port 42 nsew signal input
rlabel metal2 s 157982 279200 158038 280000 6 Di[9]
port 43 nsew signal input
rlabel metal2 s 1306 279200 1362 280000 6 Do[0]
port 44 nsew signal output
rlabel metal2 s 28722 279200 28778 280000 6 Do[10]
port 45 nsew signal output
rlabel metal2 s 31482 279200 31538 280000 6 Do[11]
port 46 nsew signal output
rlabel metal2 s 34242 279200 34298 280000 6 Do[12]
port 47 nsew signal output
rlabel metal2 s 37002 279200 37058 280000 6 Do[13]
port 48 nsew signal output
rlabel metal2 s 39762 279200 39818 280000 6 Do[14]
port 49 nsew signal output
rlabel metal2 s 42522 279200 42578 280000 6 Do[15]
port 50 nsew signal output
rlabel metal2 s 45282 279200 45338 280000 6 Do[16]
port 51 nsew signal output
rlabel metal2 s 48042 279200 48098 280000 6 Do[17]
port 52 nsew signal output
rlabel metal2 s 50710 279200 50766 280000 6 Do[18]
port 53 nsew signal output
rlabel metal2 s 53470 279200 53526 280000 6 Do[19]
port 54 nsew signal output
rlabel metal2 s 3974 279200 4030 280000 6 Do[1]
port 55 nsew signal output
rlabel metal2 s 56230 279200 56286 280000 6 Do[20]
port 56 nsew signal output
rlabel metal2 s 58990 279200 59046 280000 6 Do[21]
port 57 nsew signal output
rlabel metal2 s 61750 279200 61806 280000 6 Do[22]
port 58 nsew signal output
rlabel metal2 s 64510 279200 64566 280000 6 Do[23]
port 59 nsew signal output
rlabel metal2 s 67270 279200 67326 280000 6 Do[24]
port 60 nsew signal output
rlabel metal2 s 70030 279200 70086 280000 6 Do[25]
port 61 nsew signal output
rlabel metal2 s 72790 279200 72846 280000 6 Do[26]
port 62 nsew signal output
rlabel metal2 s 75458 279200 75514 280000 6 Do[27]
port 63 nsew signal output
rlabel metal2 s 78218 279200 78274 280000 6 Do[28]
port 64 nsew signal output
rlabel metal2 s 80978 279200 81034 280000 6 Do[29]
port 65 nsew signal output
rlabel metal2 s 6734 279200 6790 280000 6 Do[2]
port 66 nsew signal output
rlabel metal2 s 83738 279200 83794 280000 6 Do[30]
port 67 nsew signal output
rlabel metal2 s 86498 279200 86554 280000 6 Do[31]
port 68 nsew signal output
rlabel metal2 s 9494 279200 9550 280000 6 Do[3]
port 69 nsew signal output
rlabel metal2 s 12254 279200 12310 280000 6 Do[4]
port 70 nsew signal output
rlabel metal2 s 15014 279200 15070 280000 6 Do[5]
port 71 nsew signal output
rlabel metal2 s 17774 279200 17830 280000 6 Do[6]
port 72 nsew signal output
rlabel metal2 s 20534 279200 20590 280000 6 Do[7]
port 73 nsew signal output
rlabel metal2 s 23294 279200 23350 280000 6 Do[8]
port 74 nsew signal output
rlabel metal2 s 25962 279200 26018 280000 6 Do[9]
port 75 nsew signal output
rlabel metal2 s 130474 279200 130530 280000 6 EN
port 76 nsew signal input
rlabel metal2 s 119526 279200 119582 280000 6 WE[0]
port 77 nsew signal input
rlabel metal2 s 122286 279200 122342 280000 6 WE[1]
port 78 nsew signal input
rlabel metal2 s 124954 279200 125010 280000 6 WE[2]
port 79 nsew signal input
rlabel metal2 s 127714 279200 127770 280000 6 WE[3]
port 80 nsew signal input
rlabel metal4 s 188528 2128 188848 277488 6 vccd1
port 81 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 277488 6 vccd1
port 82 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 277488 6 vccd1
port 83 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 277488 6 vccd1
port 84 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 277488 6 vccd1
port 85 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 277488 6 vccd1
port 86 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 277488 6 vccd1
port 87 nsew power bidirectional
rlabel metal4 s 203888 2128 204208 277488 6 vssd1
port 88 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 277488 6 vssd1
port 89 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 277488 6 vssd1
port 90 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 277488 6 vssd1
port 91 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 277488 6 vssd1
port 92 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 277488 6 vssd1
port 93 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 277488 6 vssd1
port 94 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 220000 280000
string LEFview TRUE
string GDS_FILE /project/openlane/DFFRAM_1Kx32/runs/DFFRAM_1Kx32/results/magic/DFFRAM_1Kx32.gds
string GDS_END 237891996
string GDS_START 181870
<< end >>

