VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO DMC_32x16HC
  CLASS BLOCK ;
  FOREIGN DMC_32x16HC ;
  ORIGIN 0.000 0.000 ;
  SIZE 400.000 BY 600.000 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 596.000 2.670 600.000 ;
    END
  END A[0]
  PIN A[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 596.000 56.490 600.000 ;
    END
  END A[10]
  PIN A[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 596.000 62.010 600.000 ;
    END
  END A[11]
  PIN A[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.250 596.000 67.530 600.000 ;
    END
  END A[12]
  PIN A[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 596.000 72.590 600.000 ;
    END
  END A[13]
  PIN A[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 596.000 78.110 600.000 ;
    END
  END A[14]
  PIN A[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 596.000 83.630 600.000 ;
    END
  END A[15]
  PIN A[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 596.000 89.150 600.000 ;
    END
  END A[16]
  PIN A[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 596.000 94.210 600.000 ;
    END
  END A[17]
  PIN A[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.450 596.000 99.730 600.000 ;
    END
  END A[18]
  PIN A[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.970 596.000 105.250 600.000 ;
    END
  END A[19]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 596.000 7.730 600.000 ;
    END
  END A[1]
  PIN A[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.490 596.000 110.770 600.000 ;
    END
  END A[20]
  PIN A[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.550 596.000 115.830 600.000 ;
    END
  END A[21]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 596.000 13.250 600.000 ;
    END
  END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 596.000 18.770 600.000 ;
    END
  END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 596.000 24.290 600.000 ;
    END
  END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 596.000 29.350 600.000 ;
    END
  END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 596.000 34.870 600.000 ;
    END
  END A[6]
  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 596.000 40.390 600.000 ;
    END
  END A[7]
  PIN A[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 596.000 45.910 600.000 ;
    END
  END A[8]
  PIN A[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 596.000 50.970 600.000 ;
    END
  END A[9]
  PIN A_h[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.070 596.000 121.350 600.000 ;
    END
  END A_h[0]
  PIN A_h[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.350 596.000 175.630 600.000 ;
    END
  END A_h[10]
  PIN A_h[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 596.000 180.690 600.000 ;
    END
  END A_h[11]
  PIN A_h[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.930 596.000 186.210 600.000 ;
    END
  END A_h[12]
  PIN A_h[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.450 596.000 191.730 600.000 ;
    END
  END A_h[13]
  PIN A_h[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.970 596.000 197.250 600.000 ;
    END
  END A_h[14]
  PIN A_h[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.490 596.000 202.770 600.000 ;
    END
  END A_h[15]
  PIN A_h[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.550 596.000 207.830 600.000 ;
    END
  END A_h[16]
  PIN A_h[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.070 596.000 213.350 600.000 ;
    END
  END A_h[17]
  PIN A_h[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.590 596.000 218.870 600.000 ;
    END
  END A_h[18]
  PIN A_h[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.110 596.000 224.390 600.000 ;
    END
  END A_h[19]
  PIN A_h[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.590 596.000 126.870 600.000 ;
    END
  END A_h[1]
  PIN A_h[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 596.000 132.390 600.000 ;
    END
  END A_h[2]
  PIN A_h[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.170 596.000 137.450 600.000 ;
    END
  END A_h[3]
  PIN A_h[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 596.000 142.970 600.000 ;
    END
  END A_h[4]
  PIN A_h[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 596.000 148.490 600.000 ;
    END
  END A_h[5]
  PIN A_h[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.730 596.000 154.010 600.000 ;
    END
  END A_h[6]
  PIN A_h[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.790 596.000 159.070 600.000 ;
    END
  END A_h[7]
  PIN A_h[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 596.000 164.590 600.000 ;
    END
  END A_h[8]
  PIN A_h[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.830 596.000 170.110 600.000 ;
    END
  END A_h[9]
  PIN Do[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.170 596.000 229.450 600.000 ;
    END
  END Do[0]
  PIN Do[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 596.000 283.730 600.000 ;
    END
  END Do[10]
  PIN Do[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.970 596.000 289.250 600.000 ;
    END
  END Do[11]
  PIN Do[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.030 596.000 294.310 600.000 ;
    END
  END Do[12]
  PIN Do[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 596.000 299.830 600.000 ;
    END
  END Do[13]
  PIN Do[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.070 596.000 305.350 600.000 ;
    END
  END Do[14]
  PIN Do[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.590 596.000 310.870 600.000 ;
    END
  END Do[15]
  PIN Do[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 596.000 315.930 600.000 ;
    END
  END Do[16]
  PIN Do[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.170 596.000 321.450 600.000 ;
    END
  END Do[17]
  PIN Do[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.690 596.000 326.970 600.000 ;
    END
  END Do[18]
  PIN Do[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.210 596.000 332.490 600.000 ;
    END
  END Do[19]
  PIN Do[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 596.000 234.970 600.000 ;
    END
  END Do[1]
  PIN Do[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.270 596.000 337.550 600.000 ;
    END
  END Do[20]
  PIN Do[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.790 596.000 343.070 600.000 ;
    END
  END Do[21]
  PIN Do[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.310 596.000 348.590 600.000 ;
    END
  END Do[22]
  PIN Do[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.830 596.000 354.110 600.000 ;
    END
  END Do[23]
  PIN Do[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.890 596.000 359.170 600.000 ;
    END
  END Do[24]
  PIN Do[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.410 596.000 364.690 600.000 ;
    END
  END Do[25]
  PIN Do[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.930 596.000 370.210 600.000 ;
    END
  END Do[26]
  PIN Do[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.450 596.000 375.730 600.000 ;
    END
  END Do[27]
  PIN Do[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.510 596.000 380.790 600.000 ;
    END
  END Do[28]
  PIN Do[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.030 596.000 386.310 600.000 ;
    END
  END Do[29]
  PIN Do[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.210 596.000 240.490 600.000 ;
    END
  END Do[2]
  PIN Do[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.550 596.000 391.830 600.000 ;
    END
  END Do[30]
  PIN Do[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.070 596.000 397.350 600.000 ;
    END
  END Do[31]
  PIN Do[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.730 596.000 246.010 600.000 ;
    END
  END Do[3]
  PIN Do[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.790 596.000 251.070 600.000 ;
    END
  END Do[4]
  PIN Do[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.310 596.000 256.590 600.000 ;
    END
  END Do[5]
  PIN Do[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.830 596.000 262.110 600.000 ;
    END
  END Do[6]
  PIN Do[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 596.000 267.630 600.000 ;
    END
  END Do[7]
  PIN Do[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.410 596.000 272.690 600.000 ;
    END
  END Do[8]
  PIN Do[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.930 596.000 278.210 600.000 ;
    END
  END Do[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 4.000 ;
    END
  END clk
  PIN hit
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.690 0.000 349.970 4.000 ;
    END
  END hit
  PIN line[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 2.080 400.000 2.680 ;
    END
  END line[0]
  PIN line[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 470.600 400.000 471.200 ;
    END
  END line[100]
  PIN line[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 474.680 400.000 475.280 ;
    END
  END line[101]
  PIN line[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 479.440 400.000 480.040 ;
    END
  END line[102]
  PIN line[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 484.200 400.000 484.800 ;
    END
  END line[103]
  PIN line[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 488.960 400.000 489.560 ;
    END
  END line[104]
  PIN line[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 493.720 400.000 494.320 ;
    END
  END line[105]
  PIN line[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 498.480 400.000 499.080 ;
    END
  END line[106]
  PIN line[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 503.240 400.000 503.840 ;
    END
  END line[107]
  PIN line[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 508.000 400.000 508.600 ;
    END
  END line[108]
  PIN line[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 512.760 400.000 513.360 ;
    END
  END line[109]
  PIN line[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 48.320 400.000 48.920 ;
    END
  END line[10]
  PIN line[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 516.840 400.000 517.440 ;
    END
  END line[110]
  PIN line[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 521.600 400.000 522.200 ;
    END
  END line[111]
  PIN line[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 526.360 400.000 526.960 ;
    END
  END line[112]
  PIN line[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 531.120 400.000 531.720 ;
    END
  END line[113]
  PIN line[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 535.880 400.000 536.480 ;
    END
  END line[114]
  PIN line[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 540.640 400.000 541.240 ;
    END
  END line[115]
  PIN line[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 545.400 400.000 546.000 ;
    END
  END line[116]
  PIN line[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 550.160 400.000 550.760 ;
    END
  END line[117]
  PIN line[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 554.920 400.000 555.520 ;
    END
  END line[118]
  PIN line[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 559.000 400.000 559.600 ;
    END
  END line[119]
  PIN line[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 53.080 400.000 53.680 ;
    END
  END line[11]
  PIN line[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 563.760 400.000 564.360 ;
    END
  END line[120]
  PIN line[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 568.520 400.000 569.120 ;
    END
  END line[121]
  PIN line[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 573.280 400.000 573.880 ;
    END
  END line[122]
  PIN line[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 578.040 400.000 578.640 ;
    END
  END line[123]
  PIN line[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 582.800 400.000 583.400 ;
    END
  END line[124]
  PIN line[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 587.560 400.000 588.160 ;
    END
  END line[125]
  PIN line[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 592.320 400.000 592.920 ;
    END
  END line[126]
  PIN line[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 597.080 400.000 597.680 ;
    END
  END line[127]
  PIN line[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 57.840 400.000 58.440 ;
    END
  END line[12]
  PIN line[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 62.600 400.000 63.200 ;
    END
  END line[13]
  PIN line[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 67.360 400.000 67.960 ;
    END
  END line[14]
  PIN line[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 72.120 400.000 72.720 ;
    END
  END line[15]
  PIN line[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 76.880 400.000 77.480 ;
    END
  END line[16]
  PIN line[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 81.640 400.000 82.240 ;
    END
  END line[17]
  PIN line[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 86.400 400.000 87.000 ;
    END
  END line[18]
  PIN line[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 90.480 400.000 91.080 ;
    END
  END line[19]
  PIN line[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 6.160 400.000 6.760 ;
    END
  END line[1]
  PIN line[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 95.240 400.000 95.840 ;
    END
  END line[20]
  PIN line[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 100.000 400.000 100.600 ;
    END
  END line[21]
  PIN line[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 104.760 400.000 105.360 ;
    END
  END line[22]
  PIN line[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 109.520 400.000 110.120 ;
    END
  END line[23]
  PIN line[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 114.280 400.000 114.880 ;
    END
  END line[24]
  PIN line[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 119.040 400.000 119.640 ;
    END
  END line[25]
  PIN line[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 123.800 400.000 124.400 ;
    END
  END line[26]
  PIN line[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 128.560 400.000 129.160 ;
    END
  END line[27]
  PIN line[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 132.640 400.000 133.240 ;
    END
  END line[28]
  PIN line[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 137.400 400.000 138.000 ;
    END
  END line[29]
  PIN line[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 10.920 400.000 11.520 ;
    END
  END line[2]
  PIN line[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 142.160 400.000 142.760 ;
    END
  END line[30]
  PIN line[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 146.920 400.000 147.520 ;
    END
  END line[31]
  PIN line[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 151.680 400.000 152.280 ;
    END
  END line[32]
  PIN line[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 156.440 400.000 157.040 ;
    END
  END line[33]
  PIN line[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 161.200 400.000 161.800 ;
    END
  END line[34]
  PIN line[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 165.960 400.000 166.560 ;
    END
  END line[35]
  PIN line[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 170.720 400.000 171.320 ;
    END
  END line[36]
  PIN line[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 174.800 400.000 175.400 ;
    END
  END line[37]
  PIN line[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 179.560 400.000 180.160 ;
    END
  END line[38]
  PIN line[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 184.320 400.000 184.920 ;
    END
  END line[39]
  PIN line[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 15.680 400.000 16.280 ;
    END
  END line[3]
  PIN line[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 189.080 400.000 189.680 ;
    END
  END line[40]
  PIN line[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 193.840 400.000 194.440 ;
    END
  END line[41]
  PIN line[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 198.600 400.000 199.200 ;
    END
  END line[42]
  PIN line[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 203.360 400.000 203.960 ;
    END
  END line[43]
  PIN line[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 208.120 400.000 208.720 ;
    END
  END line[44]
  PIN line[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 212.880 400.000 213.480 ;
    END
  END line[45]
  PIN line[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 216.960 400.000 217.560 ;
    END
  END line[46]
  PIN line[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 221.720 400.000 222.320 ;
    END
  END line[47]
  PIN line[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 226.480 400.000 227.080 ;
    END
  END line[48]
  PIN line[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 231.240 400.000 231.840 ;
    END
  END line[49]
  PIN line[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 20.440 400.000 21.040 ;
    END
  END line[4]
  PIN line[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 236.000 400.000 236.600 ;
    END
  END line[50]
  PIN line[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 240.760 400.000 241.360 ;
    END
  END line[51]
  PIN line[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 245.520 400.000 246.120 ;
    END
  END line[52]
  PIN line[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 250.280 400.000 250.880 ;
    END
  END line[53]
  PIN line[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 255.040 400.000 255.640 ;
    END
  END line[54]
  PIN line[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 259.120 400.000 259.720 ;
    END
  END line[55]
  PIN line[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 263.880 400.000 264.480 ;
    END
  END line[56]
  PIN line[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 268.640 400.000 269.240 ;
    END
  END line[57]
  PIN line[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 273.400 400.000 274.000 ;
    END
  END line[58]
  PIN line[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 278.160 400.000 278.760 ;
    END
  END line[59]
  PIN line[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 25.200 400.000 25.800 ;
    END
  END line[5]
  PIN line[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 282.920 400.000 283.520 ;
    END
  END line[60]
  PIN line[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 287.680 400.000 288.280 ;
    END
  END line[61]
  PIN line[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 292.440 400.000 293.040 ;
    END
  END line[62]
  PIN line[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 297.200 400.000 297.800 ;
    END
  END line[63]
  PIN line[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 301.960 400.000 302.560 ;
    END
  END line[64]
  PIN line[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 306.040 400.000 306.640 ;
    END
  END line[65]
  PIN line[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 310.800 400.000 311.400 ;
    END
  END line[66]
  PIN line[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 315.560 400.000 316.160 ;
    END
  END line[67]
  PIN line[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 320.320 400.000 320.920 ;
    END
  END line[68]
  PIN line[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 325.080 400.000 325.680 ;
    END
  END line[69]
  PIN line[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 29.960 400.000 30.560 ;
    END
  END line[6]
  PIN line[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 329.840 400.000 330.440 ;
    END
  END line[70]
  PIN line[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 334.600 400.000 335.200 ;
    END
  END line[71]
  PIN line[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 339.360 400.000 339.960 ;
    END
  END line[72]
  PIN line[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 344.120 400.000 344.720 ;
    END
  END line[73]
  PIN line[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 348.200 400.000 348.800 ;
    END
  END line[74]
  PIN line[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 352.960 400.000 353.560 ;
    END
  END line[75]
  PIN line[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 357.720 400.000 358.320 ;
    END
  END line[76]
  PIN line[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 362.480 400.000 363.080 ;
    END
  END line[77]
  PIN line[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 367.240 400.000 367.840 ;
    END
  END line[78]
  PIN line[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 372.000 400.000 372.600 ;
    END
  END line[79]
  PIN line[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 34.720 400.000 35.320 ;
    END
  END line[7]
  PIN line[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 376.760 400.000 377.360 ;
    END
  END line[80]
  PIN line[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 381.520 400.000 382.120 ;
    END
  END line[81]
  PIN line[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 386.280 400.000 386.880 ;
    END
  END line[82]
  PIN line[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 390.360 400.000 390.960 ;
    END
  END line[83]
  PIN line[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 395.120 400.000 395.720 ;
    END
  END line[84]
  PIN line[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 399.880 400.000 400.480 ;
    END
  END line[85]
  PIN line[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 404.640 400.000 405.240 ;
    END
  END line[86]
  PIN line[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 409.400 400.000 410.000 ;
    END
  END line[87]
  PIN line[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 414.160 400.000 414.760 ;
    END
  END line[88]
  PIN line[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 418.920 400.000 419.520 ;
    END
  END line[89]
  PIN line[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 39.480 400.000 40.080 ;
    END
  END line[8]
  PIN line[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 423.680 400.000 424.280 ;
    END
  END line[90]
  PIN line[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 428.440 400.000 429.040 ;
    END
  END line[91]
  PIN line[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 432.520 400.000 433.120 ;
    END
  END line[92]
  PIN line[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 437.280 400.000 437.880 ;
    END
  END line[93]
  PIN line[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 442.040 400.000 442.640 ;
    END
  END line[94]
  PIN line[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 446.800 400.000 447.400 ;
    END
  END line[95]
  PIN line[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 451.560 400.000 452.160 ;
    END
  END line[96]
  PIN line[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 456.320 400.000 456.920 ;
    END
  END line[97]
  PIN line[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 461.080 400.000 461.680 ;
    END
  END line[98]
  PIN line[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 465.840 400.000 466.440 ;
    END
  END line[99]
  PIN line[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 44.240 400.000 44.840 ;
    END
  END line[9]
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 0.000 149.870 4.000 ;
    END
  END rst_n
  PIN wr
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.870 0.000 250.150 4.000 ;
    END
  END wr
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 587.760 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 587.760 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 587.760 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 587.760 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 587.760 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 395.455 587.605 ;
      LAYER met1 ;
        RECT 5.520 6.160 397.370 587.760 ;
      LAYER met2 ;
        RECT 0.090 595.720 2.110 597.565 ;
        RECT 2.950 595.720 7.170 597.565 ;
        RECT 8.010 595.720 12.690 597.565 ;
        RECT 13.530 595.720 18.210 597.565 ;
        RECT 19.050 595.720 23.730 597.565 ;
        RECT 24.570 595.720 28.790 597.565 ;
        RECT 29.630 595.720 34.310 597.565 ;
        RECT 35.150 595.720 39.830 597.565 ;
        RECT 40.670 595.720 45.350 597.565 ;
        RECT 46.190 595.720 50.410 597.565 ;
        RECT 51.250 595.720 55.930 597.565 ;
        RECT 56.770 595.720 61.450 597.565 ;
        RECT 62.290 595.720 66.970 597.565 ;
        RECT 67.810 595.720 72.030 597.565 ;
        RECT 72.870 595.720 77.550 597.565 ;
        RECT 78.390 595.720 83.070 597.565 ;
        RECT 83.910 595.720 88.590 597.565 ;
        RECT 89.430 595.720 93.650 597.565 ;
        RECT 94.490 595.720 99.170 597.565 ;
        RECT 100.010 595.720 104.690 597.565 ;
        RECT 105.530 595.720 110.210 597.565 ;
        RECT 111.050 595.720 115.270 597.565 ;
        RECT 116.110 595.720 120.790 597.565 ;
        RECT 121.630 595.720 126.310 597.565 ;
        RECT 127.150 595.720 131.830 597.565 ;
        RECT 132.670 595.720 136.890 597.565 ;
        RECT 137.730 595.720 142.410 597.565 ;
        RECT 143.250 595.720 147.930 597.565 ;
        RECT 148.770 595.720 153.450 597.565 ;
        RECT 154.290 595.720 158.510 597.565 ;
        RECT 159.350 595.720 164.030 597.565 ;
        RECT 164.870 595.720 169.550 597.565 ;
        RECT 170.390 595.720 175.070 597.565 ;
        RECT 175.910 595.720 180.130 597.565 ;
        RECT 180.970 595.720 185.650 597.565 ;
        RECT 186.490 595.720 191.170 597.565 ;
        RECT 192.010 595.720 196.690 597.565 ;
        RECT 197.530 595.720 202.210 597.565 ;
        RECT 203.050 595.720 207.270 597.565 ;
        RECT 208.110 595.720 212.790 597.565 ;
        RECT 213.630 595.720 218.310 597.565 ;
        RECT 219.150 595.720 223.830 597.565 ;
        RECT 224.670 595.720 228.890 597.565 ;
        RECT 229.730 595.720 234.410 597.565 ;
        RECT 235.250 595.720 239.930 597.565 ;
        RECT 240.770 595.720 245.450 597.565 ;
        RECT 246.290 595.720 250.510 597.565 ;
        RECT 251.350 595.720 256.030 597.565 ;
        RECT 256.870 595.720 261.550 597.565 ;
        RECT 262.390 595.720 267.070 597.565 ;
        RECT 267.910 595.720 272.130 597.565 ;
        RECT 272.970 595.720 277.650 597.565 ;
        RECT 278.490 595.720 283.170 597.565 ;
        RECT 284.010 595.720 288.690 597.565 ;
        RECT 289.530 595.720 293.750 597.565 ;
        RECT 294.590 595.720 299.270 597.565 ;
        RECT 300.110 595.720 304.790 597.565 ;
        RECT 305.630 595.720 310.310 597.565 ;
        RECT 311.150 595.720 315.370 597.565 ;
        RECT 316.210 595.720 320.890 597.565 ;
        RECT 321.730 595.720 326.410 597.565 ;
        RECT 327.250 595.720 331.930 597.565 ;
        RECT 332.770 595.720 336.990 597.565 ;
        RECT 337.830 595.720 342.510 597.565 ;
        RECT 343.350 595.720 348.030 597.565 ;
        RECT 348.870 595.720 353.550 597.565 ;
        RECT 354.390 595.720 358.610 597.565 ;
        RECT 359.450 595.720 364.130 597.565 ;
        RECT 364.970 595.720 369.650 597.565 ;
        RECT 370.490 595.720 375.170 597.565 ;
        RECT 376.010 595.720 380.230 597.565 ;
        RECT 381.070 595.720 385.750 597.565 ;
        RECT 386.590 595.720 391.270 597.565 ;
        RECT 392.110 595.720 396.790 597.565 ;
        RECT 0.090 4.280 397.340 595.720 ;
        RECT 0.090 2.195 49.490 4.280 ;
        RECT 50.330 2.195 149.310 4.280 ;
        RECT 150.150 2.195 249.590 4.280 ;
        RECT 250.430 2.195 349.410 4.280 ;
        RECT 350.250 2.195 397.340 4.280 ;
      LAYER met3 ;
        RECT 0.065 596.680 395.600 597.545 ;
        RECT 0.065 593.320 396.000 596.680 ;
        RECT 0.065 591.920 395.600 593.320 ;
        RECT 0.065 588.560 396.000 591.920 ;
        RECT 0.065 587.160 395.600 588.560 ;
        RECT 0.065 583.800 396.000 587.160 ;
        RECT 0.065 582.400 395.600 583.800 ;
        RECT 0.065 579.040 396.000 582.400 ;
        RECT 0.065 577.640 395.600 579.040 ;
        RECT 0.065 574.280 396.000 577.640 ;
        RECT 0.065 572.880 395.600 574.280 ;
        RECT 0.065 569.520 396.000 572.880 ;
        RECT 0.065 568.120 395.600 569.520 ;
        RECT 0.065 564.760 396.000 568.120 ;
        RECT 0.065 563.360 395.600 564.760 ;
        RECT 0.065 560.000 396.000 563.360 ;
        RECT 0.065 558.600 395.600 560.000 ;
        RECT 0.065 555.920 396.000 558.600 ;
        RECT 0.065 554.520 395.600 555.920 ;
        RECT 0.065 551.160 396.000 554.520 ;
        RECT 0.065 549.760 395.600 551.160 ;
        RECT 0.065 546.400 396.000 549.760 ;
        RECT 0.065 545.000 395.600 546.400 ;
        RECT 0.065 541.640 396.000 545.000 ;
        RECT 0.065 540.240 395.600 541.640 ;
        RECT 0.065 536.880 396.000 540.240 ;
        RECT 0.065 535.480 395.600 536.880 ;
        RECT 0.065 532.120 396.000 535.480 ;
        RECT 0.065 530.720 395.600 532.120 ;
        RECT 0.065 527.360 396.000 530.720 ;
        RECT 0.065 525.960 395.600 527.360 ;
        RECT 0.065 522.600 396.000 525.960 ;
        RECT 0.065 521.200 395.600 522.600 ;
        RECT 0.065 517.840 396.000 521.200 ;
        RECT 0.065 516.440 395.600 517.840 ;
        RECT 0.065 513.760 396.000 516.440 ;
        RECT 0.065 512.360 395.600 513.760 ;
        RECT 0.065 509.000 396.000 512.360 ;
        RECT 0.065 507.600 395.600 509.000 ;
        RECT 0.065 504.240 396.000 507.600 ;
        RECT 0.065 502.840 395.600 504.240 ;
        RECT 0.065 499.480 396.000 502.840 ;
        RECT 0.065 498.080 395.600 499.480 ;
        RECT 0.065 494.720 396.000 498.080 ;
        RECT 0.065 493.320 395.600 494.720 ;
        RECT 0.065 489.960 396.000 493.320 ;
        RECT 0.065 488.560 395.600 489.960 ;
        RECT 0.065 485.200 396.000 488.560 ;
        RECT 0.065 483.800 395.600 485.200 ;
        RECT 0.065 480.440 396.000 483.800 ;
        RECT 0.065 479.040 395.600 480.440 ;
        RECT 0.065 475.680 396.000 479.040 ;
        RECT 0.065 474.280 395.600 475.680 ;
        RECT 0.065 471.600 396.000 474.280 ;
        RECT 0.065 470.200 395.600 471.600 ;
        RECT 0.065 466.840 396.000 470.200 ;
        RECT 0.065 465.440 395.600 466.840 ;
        RECT 0.065 462.080 396.000 465.440 ;
        RECT 0.065 460.680 395.600 462.080 ;
        RECT 0.065 457.320 396.000 460.680 ;
        RECT 0.065 455.920 395.600 457.320 ;
        RECT 0.065 452.560 396.000 455.920 ;
        RECT 0.065 451.160 395.600 452.560 ;
        RECT 0.065 447.800 396.000 451.160 ;
        RECT 0.065 446.400 395.600 447.800 ;
        RECT 0.065 443.040 396.000 446.400 ;
        RECT 0.065 441.640 395.600 443.040 ;
        RECT 0.065 438.280 396.000 441.640 ;
        RECT 0.065 436.880 395.600 438.280 ;
        RECT 0.065 433.520 396.000 436.880 ;
        RECT 0.065 432.120 395.600 433.520 ;
        RECT 0.065 429.440 396.000 432.120 ;
        RECT 0.065 428.040 395.600 429.440 ;
        RECT 0.065 424.680 396.000 428.040 ;
        RECT 0.065 423.280 395.600 424.680 ;
        RECT 0.065 419.920 396.000 423.280 ;
        RECT 0.065 418.520 395.600 419.920 ;
        RECT 0.065 415.160 396.000 418.520 ;
        RECT 0.065 413.760 395.600 415.160 ;
        RECT 0.065 410.400 396.000 413.760 ;
        RECT 0.065 409.000 395.600 410.400 ;
        RECT 0.065 405.640 396.000 409.000 ;
        RECT 0.065 404.240 395.600 405.640 ;
        RECT 0.065 400.880 396.000 404.240 ;
        RECT 0.065 399.480 395.600 400.880 ;
        RECT 0.065 396.120 396.000 399.480 ;
        RECT 0.065 394.720 395.600 396.120 ;
        RECT 0.065 391.360 396.000 394.720 ;
        RECT 0.065 389.960 395.600 391.360 ;
        RECT 0.065 387.280 396.000 389.960 ;
        RECT 0.065 385.880 395.600 387.280 ;
        RECT 0.065 382.520 396.000 385.880 ;
        RECT 0.065 381.120 395.600 382.520 ;
        RECT 0.065 377.760 396.000 381.120 ;
        RECT 0.065 376.360 395.600 377.760 ;
        RECT 0.065 373.000 396.000 376.360 ;
        RECT 0.065 371.600 395.600 373.000 ;
        RECT 0.065 368.240 396.000 371.600 ;
        RECT 0.065 366.840 395.600 368.240 ;
        RECT 0.065 363.480 396.000 366.840 ;
        RECT 0.065 362.080 395.600 363.480 ;
        RECT 0.065 358.720 396.000 362.080 ;
        RECT 0.065 357.320 395.600 358.720 ;
        RECT 0.065 353.960 396.000 357.320 ;
        RECT 0.065 352.560 395.600 353.960 ;
        RECT 0.065 349.200 396.000 352.560 ;
        RECT 0.065 347.800 395.600 349.200 ;
        RECT 0.065 345.120 396.000 347.800 ;
        RECT 0.065 343.720 395.600 345.120 ;
        RECT 0.065 340.360 396.000 343.720 ;
        RECT 0.065 338.960 395.600 340.360 ;
        RECT 0.065 335.600 396.000 338.960 ;
        RECT 0.065 334.200 395.600 335.600 ;
        RECT 0.065 330.840 396.000 334.200 ;
        RECT 0.065 329.440 395.600 330.840 ;
        RECT 0.065 326.080 396.000 329.440 ;
        RECT 0.065 324.680 395.600 326.080 ;
        RECT 0.065 321.320 396.000 324.680 ;
        RECT 0.065 319.920 395.600 321.320 ;
        RECT 0.065 316.560 396.000 319.920 ;
        RECT 0.065 315.160 395.600 316.560 ;
        RECT 0.065 311.800 396.000 315.160 ;
        RECT 0.065 310.400 395.600 311.800 ;
        RECT 0.065 307.040 396.000 310.400 ;
        RECT 0.065 305.640 395.600 307.040 ;
        RECT 0.065 302.960 396.000 305.640 ;
        RECT 0.065 301.560 395.600 302.960 ;
        RECT 0.065 298.200 396.000 301.560 ;
        RECT 0.065 296.800 395.600 298.200 ;
        RECT 0.065 293.440 396.000 296.800 ;
        RECT 0.065 292.040 395.600 293.440 ;
        RECT 0.065 288.680 396.000 292.040 ;
        RECT 0.065 287.280 395.600 288.680 ;
        RECT 0.065 283.920 396.000 287.280 ;
        RECT 0.065 282.520 395.600 283.920 ;
        RECT 0.065 279.160 396.000 282.520 ;
        RECT 0.065 277.760 395.600 279.160 ;
        RECT 0.065 274.400 396.000 277.760 ;
        RECT 0.065 273.000 395.600 274.400 ;
        RECT 0.065 269.640 396.000 273.000 ;
        RECT 0.065 268.240 395.600 269.640 ;
        RECT 0.065 264.880 396.000 268.240 ;
        RECT 0.065 263.480 395.600 264.880 ;
        RECT 0.065 260.120 396.000 263.480 ;
        RECT 0.065 258.720 395.600 260.120 ;
        RECT 0.065 256.040 396.000 258.720 ;
        RECT 0.065 254.640 395.600 256.040 ;
        RECT 0.065 251.280 396.000 254.640 ;
        RECT 0.065 249.880 395.600 251.280 ;
        RECT 0.065 246.520 396.000 249.880 ;
        RECT 0.065 245.120 395.600 246.520 ;
        RECT 0.065 241.760 396.000 245.120 ;
        RECT 0.065 240.360 395.600 241.760 ;
        RECT 0.065 237.000 396.000 240.360 ;
        RECT 0.065 235.600 395.600 237.000 ;
        RECT 0.065 232.240 396.000 235.600 ;
        RECT 0.065 230.840 395.600 232.240 ;
        RECT 0.065 227.480 396.000 230.840 ;
        RECT 0.065 226.080 395.600 227.480 ;
        RECT 0.065 222.720 396.000 226.080 ;
        RECT 0.065 221.320 395.600 222.720 ;
        RECT 0.065 217.960 396.000 221.320 ;
        RECT 0.065 216.560 395.600 217.960 ;
        RECT 0.065 213.880 396.000 216.560 ;
        RECT 0.065 212.480 395.600 213.880 ;
        RECT 0.065 209.120 396.000 212.480 ;
        RECT 0.065 207.720 395.600 209.120 ;
        RECT 0.065 204.360 396.000 207.720 ;
        RECT 0.065 202.960 395.600 204.360 ;
        RECT 0.065 199.600 396.000 202.960 ;
        RECT 0.065 198.200 395.600 199.600 ;
        RECT 0.065 194.840 396.000 198.200 ;
        RECT 0.065 193.440 395.600 194.840 ;
        RECT 0.065 190.080 396.000 193.440 ;
        RECT 0.065 188.680 395.600 190.080 ;
        RECT 0.065 185.320 396.000 188.680 ;
        RECT 0.065 183.920 395.600 185.320 ;
        RECT 0.065 180.560 396.000 183.920 ;
        RECT 0.065 179.160 395.600 180.560 ;
        RECT 0.065 175.800 396.000 179.160 ;
        RECT 0.065 174.400 395.600 175.800 ;
        RECT 0.065 171.720 396.000 174.400 ;
        RECT 0.065 170.320 395.600 171.720 ;
        RECT 0.065 166.960 396.000 170.320 ;
        RECT 0.065 165.560 395.600 166.960 ;
        RECT 0.065 162.200 396.000 165.560 ;
        RECT 0.065 160.800 395.600 162.200 ;
        RECT 0.065 157.440 396.000 160.800 ;
        RECT 0.065 156.040 395.600 157.440 ;
        RECT 0.065 152.680 396.000 156.040 ;
        RECT 0.065 151.280 395.600 152.680 ;
        RECT 0.065 147.920 396.000 151.280 ;
        RECT 0.065 146.520 395.600 147.920 ;
        RECT 0.065 143.160 396.000 146.520 ;
        RECT 0.065 141.760 395.600 143.160 ;
        RECT 0.065 138.400 396.000 141.760 ;
        RECT 0.065 137.000 395.600 138.400 ;
        RECT 0.065 133.640 396.000 137.000 ;
        RECT 0.065 132.240 395.600 133.640 ;
        RECT 0.065 129.560 396.000 132.240 ;
        RECT 0.065 128.160 395.600 129.560 ;
        RECT 0.065 124.800 396.000 128.160 ;
        RECT 0.065 123.400 395.600 124.800 ;
        RECT 0.065 120.040 396.000 123.400 ;
        RECT 0.065 118.640 395.600 120.040 ;
        RECT 0.065 115.280 396.000 118.640 ;
        RECT 0.065 113.880 395.600 115.280 ;
        RECT 0.065 110.520 396.000 113.880 ;
        RECT 0.065 109.120 395.600 110.520 ;
        RECT 0.065 105.760 396.000 109.120 ;
        RECT 0.065 104.360 395.600 105.760 ;
        RECT 0.065 101.000 396.000 104.360 ;
        RECT 0.065 99.600 395.600 101.000 ;
        RECT 0.065 96.240 396.000 99.600 ;
        RECT 0.065 94.840 395.600 96.240 ;
        RECT 0.065 91.480 396.000 94.840 ;
        RECT 0.065 90.080 395.600 91.480 ;
        RECT 0.065 87.400 396.000 90.080 ;
        RECT 0.065 86.000 395.600 87.400 ;
        RECT 0.065 82.640 396.000 86.000 ;
        RECT 0.065 81.240 395.600 82.640 ;
        RECT 0.065 77.880 396.000 81.240 ;
        RECT 0.065 76.480 395.600 77.880 ;
        RECT 0.065 73.120 396.000 76.480 ;
        RECT 0.065 71.720 395.600 73.120 ;
        RECT 0.065 68.360 396.000 71.720 ;
        RECT 0.065 66.960 395.600 68.360 ;
        RECT 0.065 63.600 396.000 66.960 ;
        RECT 0.065 62.200 395.600 63.600 ;
        RECT 0.065 58.840 396.000 62.200 ;
        RECT 0.065 57.440 395.600 58.840 ;
        RECT 0.065 54.080 396.000 57.440 ;
        RECT 0.065 52.680 395.600 54.080 ;
        RECT 0.065 49.320 396.000 52.680 ;
        RECT 0.065 47.920 395.600 49.320 ;
        RECT 0.065 45.240 396.000 47.920 ;
        RECT 0.065 43.840 395.600 45.240 ;
        RECT 0.065 40.480 396.000 43.840 ;
        RECT 0.065 39.080 395.600 40.480 ;
        RECT 0.065 35.720 396.000 39.080 ;
        RECT 0.065 34.320 395.600 35.720 ;
        RECT 0.065 30.960 396.000 34.320 ;
        RECT 0.065 29.560 395.600 30.960 ;
        RECT 0.065 26.200 396.000 29.560 ;
        RECT 0.065 24.800 395.600 26.200 ;
        RECT 0.065 21.440 396.000 24.800 ;
        RECT 0.065 20.040 395.600 21.440 ;
        RECT 0.065 16.680 396.000 20.040 ;
        RECT 0.065 15.280 395.600 16.680 ;
        RECT 0.065 11.920 396.000 15.280 ;
        RECT 0.065 10.520 395.600 11.920 ;
        RECT 0.065 7.160 396.000 10.520 ;
        RECT 0.065 5.760 395.600 7.160 ;
        RECT 0.065 3.080 396.000 5.760 ;
        RECT 0.065 2.215 395.600 3.080 ;
      LAYER met4 ;
        RECT 71.135 26.015 97.440 573.065 ;
        RECT 99.840 26.015 174.240 573.065 ;
        RECT 176.640 26.015 251.040 573.065 ;
        RECT 253.440 26.015 327.840 573.065 ;
        RECT 330.240 26.015 373.225 573.065 ;
  END
END DMC_32x16HC
END LIBRARY

