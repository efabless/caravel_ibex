magic
tech sky130A
magscale 1 2
timestamp 1621723670
<< obsli1 >>
rect 1104 1445 118864 157777
<< obsm1 >>
rect 474 1232 119494 157808
<< metal2 >>
rect 478 0 534 800
rect 1398 0 1454 800
rect 2410 0 2466 800
rect 3422 0 3478 800
rect 4434 0 4490 800
rect 5446 0 5502 800
rect 6458 0 6514 800
rect 7470 0 7526 800
rect 8390 0 8446 800
rect 9402 0 9458 800
rect 10414 0 10470 800
rect 11426 0 11482 800
rect 12438 0 12494 800
rect 13450 0 13506 800
rect 14462 0 14518 800
rect 15474 0 15530 800
rect 16394 0 16450 800
rect 17406 0 17462 800
rect 18418 0 18474 800
rect 19430 0 19486 800
rect 20442 0 20498 800
rect 21454 0 21510 800
rect 22466 0 22522 800
rect 23386 0 23442 800
rect 24398 0 24454 800
rect 25410 0 25466 800
rect 26422 0 26478 800
rect 27434 0 27490 800
rect 28446 0 28502 800
rect 29458 0 29514 800
rect 30470 0 30526 800
rect 31390 0 31446 800
rect 32402 0 32458 800
rect 33414 0 33470 800
rect 34426 0 34482 800
rect 35438 0 35494 800
rect 36450 0 36506 800
rect 37462 0 37518 800
rect 38382 0 38438 800
rect 39394 0 39450 800
rect 40406 0 40462 800
rect 41418 0 41474 800
rect 42430 0 42486 800
rect 43442 0 43498 800
rect 44454 0 44510 800
rect 45466 0 45522 800
rect 46386 0 46442 800
rect 47398 0 47454 800
rect 48410 0 48466 800
rect 49422 0 49478 800
rect 50434 0 50490 800
rect 51446 0 51502 800
rect 52458 0 52514 800
rect 53378 0 53434 800
rect 54390 0 54446 800
rect 55402 0 55458 800
rect 56414 0 56470 800
rect 57426 0 57482 800
rect 58438 0 58494 800
rect 59450 0 59506 800
rect 60462 0 60518 800
rect 61382 0 61438 800
rect 62394 0 62450 800
rect 63406 0 63462 800
rect 64418 0 64474 800
rect 65430 0 65486 800
rect 66442 0 66498 800
rect 67454 0 67510 800
rect 68374 0 68430 800
rect 69386 0 69442 800
rect 70398 0 70454 800
rect 71410 0 71466 800
rect 72422 0 72478 800
rect 73434 0 73490 800
rect 74446 0 74502 800
rect 75458 0 75514 800
rect 76378 0 76434 800
rect 77390 0 77446 800
rect 78402 0 78458 800
rect 79414 0 79470 800
rect 80426 0 80482 800
rect 81438 0 81494 800
rect 82450 0 82506 800
rect 83370 0 83426 800
rect 84382 0 84438 800
rect 85394 0 85450 800
rect 86406 0 86462 800
rect 87418 0 87474 800
rect 88430 0 88486 800
rect 89442 0 89498 800
rect 90454 0 90510 800
rect 91374 0 91430 800
rect 92386 0 92442 800
rect 93398 0 93454 800
rect 94410 0 94466 800
rect 95422 0 95478 800
rect 96434 0 96490 800
rect 97446 0 97502 800
rect 98366 0 98422 800
rect 99378 0 99434 800
rect 100390 0 100446 800
rect 101402 0 101458 800
rect 102414 0 102470 800
rect 103426 0 103482 800
rect 104438 0 104494 800
rect 105450 0 105506 800
rect 106370 0 106426 800
rect 107382 0 107438 800
rect 108394 0 108450 800
rect 109406 0 109462 800
rect 110418 0 110474 800
rect 111430 0 111486 800
rect 112442 0 112498 800
rect 113362 0 113418 800
rect 114374 0 114430 800
rect 115386 0 115442 800
rect 116398 0 116454 800
rect 117410 0 117466 800
rect 118422 0 118478 800
rect 119434 0 119490 800
<< obsm2 >>
rect 480 856 119488 157808
rect 590 800 1342 856
rect 1510 800 2354 856
rect 2522 800 3366 856
rect 3534 800 4378 856
rect 4546 800 5390 856
rect 5558 800 6402 856
rect 6570 800 7414 856
rect 7582 800 8334 856
rect 8502 800 9346 856
rect 9514 800 10358 856
rect 10526 800 11370 856
rect 11538 800 12382 856
rect 12550 800 13394 856
rect 13562 800 14406 856
rect 14574 800 15418 856
rect 15586 800 16338 856
rect 16506 800 17350 856
rect 17518 800 18362 856
rect 18530 800 19374 856
rect 19542 800 20386 856
rect 20554 800 21398 856
rect 21566 800 22410 856
rect 22578 800 23330 856
rect 23498 800 24342 856
rect 24510 800 25354 856
rect 25522 800 26366 856
rect 26534 800 27378 856
rect 27546 800 28390 856
rect 28558 800 29402 856
rect 29570 800 30414 856
rect 30582 800 31334 856
rect 31502 800 32346 856
rect 32514 800 33358 856
rect 33526 800 34370 856
rect 34538 800 35382 856
rect 35550 800 36394 856
rect 36562 800 37406 856
rect 37574 800 38326 856
rect 38494 800 39338 856
rect 39506 800 40350 856
rect 40518 800 41362 856
rect 41530 800 42374 856
rect 42542 800 43386 856
rect 43554 800 44398 856
rect 44566 800 45410 856
rect 45578 800 46330 856
rect 46498 800 47342 856
rect 47510 800 48354 856
rect 48522 800 49366 856
rect 49534 800 50378 856
rect 50546 800 51390 856
rect 51558 800 52402 856
rect 52570 800 53322 856
rect 53490 800 54334 856
rect 54502 800 55346 856
rect 55514 800 56358 856
rect 56526 800 57370 856
rect 57538 800 58382 856
rect 58550 800 59394 856
rect 59562 800 60406 856
rect 60574 800 61326 856
rect 61494 800 62338 856
rect 62506 800 63350 856
rect 63518 800 64362 856
rect 64530 800 65374 856
rect 65542 800 66386 856
rect 66554 800 67398 856
rect 67566 800 68318 856
rect 68486 800 69330 856
rect 69498 800 70342 856
rect 70510 800 71354 856
rect 71522 800 72366 856
rect 72534 800 73378 856
rect 73546 800 74390 856
rect 74558 800 75402 856
rect 75570 800 76322 856
rect 76490 800 77334 856
rect 77502 800 78346 856
rect 78514 800 79358 856
rect 79526 800 80370 856
rect 80538 800 81382 856
rect 81550 800 82394 856
rect 82562 800 83314 856
rect 83482 800 84326 856
rect 84494 800 85338 856
rect 85506 800 86350 856
rect 86518 800 87362 856
rect 87530 800 88374 856
rect 88542 800 89386 856
rect 89554 800 90398 856
rect 90566 800 91318 856
rect 91486 800 92330 856
rect 92498 800 93342 856
rect 93510 800 94354 856
rect 94522 800 95366 856
rect 95534 800 96378 856
rect 96546 800 97390 856
rect 97558 800 98310 856
rect 98478 800 99322 856
rect 99490 800 100334 856
rect 100502 800 101346 856
rect 101514 800 102358 856
rect 102526 800 103370 856
rect 103538 800 104382 856
rect 104550 800 105394 856
rect 105562 800 106314 856
rect 106482 800 107326 856
rect 107494 800 108338 856
rect 108506 800 109350 856
rect 109518 800 110362 856
rect 110530 800 111374 856
rect 111542 800 112386 856
rect 112554 800 113306 856
rect 113474 800 114318 856
rect 114486 800 115330 856
rect 115498 800 116342 856
rect 116510 800 117354 856
rect 117522 800 118366 856
rect 118534 800 119378 856
<< metal3 >>
rect 0 156680 800 156800
rect 0 150560 800 150680
rect 0 144440 800 144560
rect 0 138320 800 138440
rect 0 132064 800 132184
rect 0 125944 800 126064
rect 0 119824 800 119944
rect 0 113704 800 113824
rect 0 107448 800 107568
rect 0 101328 800 101448
rect 0 95208 800 95328
rect 0 89088 800 89208
rect 0 82968 800 83088
rect 0 76712 800 76832
rect 0 70592 800 70712
rect 0 64472 800 64592
rect 0 58352 800 58472
rect 0 52096 800 52216
rect 0 45976 800 46096
rect 0 39856 800 39976
rect 0 33736 800 33856
rect 0 27480 800 27600
rect 0 21360 800 21480
rect 0 15240 800 15360
rect 0 9120 800 9240
rect 0 3000 800 3120
<< obsm3 >>
rect 800 156880 112503 157793
rect 880 156600 112503 156880
rect 800 150760 112503 156600
rect 880 150480 112503 150760
rect 800 144640 112503 150480
rect 880 144360 112503 144640
rect 800 138520 112503 144360
rect 880 138240 112503 138520
rect 800 132264 112503 138240
rect 880 131984 112503 132264
rect 800 126144 112503 131984
rect 880 125864 112503 126144
rect 800 120024 112503 125864
rect 880 119744 112503 120024
rect 800 113904 112503 119744
rect 880 113624 112503 113904
rect 800 107648 112503 113624
rect 880 107368 112503 107648
rect 800 101528 112503 107368
rect 880 101248 112503 101528
rect 800 95408 112503 101248
rect 880 95128 112503 95408
rect 800 89288 112503 95128
rect 880 89008 112503 89288
rect 800 83168 112503 89008
rect 880 82888 112503 83168
rect 800 76912 112503 82888
rect 880 76632 112503 76912
rect 800 70792 112503 76632
rect 880 70512 112503 70792
rect 800 64672 112503 70512
rect 880 64392 112503 64672
rect 800 58552 112503 64392
rect 880 58272 112503 58552
rect 800 52296 112503 58272
rect 880 52016 112503 52296
rect 800 46176 112503 52016
rect 880 45896 112503 46176
rect 800 40056 112503 45896
rect 880 39776 112503 40056
rect 800 33936 112503 39776
rect 880 33656 112503 33936
rect 800 27680 112503 33656
rect 880 27400 112503 27680
rect 800 21560 112503 27400
rect 880 21280 112503 21560
rect 800 15440 112503 21280
rect 880 15160 112503 15440
rect 800 9320 112503 15160
rect 880 9040 112503 9320
rect 800 3200 112503 9040
rect 880 2920 112503 3200
rect 800 1939 112503 2920
<< metal4 >>
rect 4208 2128 4528 157808
rect 19568 2128 19888 157808
rect 34928 2128 35248 157808
rect 50288 2128 50608 157808
rect 65648 2128 65968 157808
rect 81008 2128 81328 157808
rect 96368 2128 96688 157808
rect 111728 2128 112048 157808
<< obsm4 >>
rect 2451 2048 4128 156093
rect 4608 2048 19488 156093
rect 19968 2048 34848 156093
rect 35328 2048 50208 156093
rect 50688 2048 65568 156093
rect 66048 2048 80928 156093
rect 81408 2048 93781 156093
rect 2451 1939 93781 2048
<< labels >>
rlabel metal3 s 0 156680 800 156800 6 EXT_IRQ
port 1 nsew signal input
rlabel metal2 s 478 0 534 800 6 HADDR[0]
port 2 nsew signal output
rlabel metal2 s 10414 0 10470 800 6 HADDR[10]
port 3 nsew signal output
rlabel metal2 s 11426 0 11482 800 6 HADDR[11]
port 4 nsew signal output
rlabel metal2 s 12438 0 12494 800 6 HADDR[12]
port 5 nsew signal output
rlabel metal2 s 13450 0 13506 800 6 HADDR[13]
port 6 nsew signal output
rlabel metal2 s 14462 0 14518 800 6 HADDR[14]
port 7 nsew signal output
rlabel metal2 s 15474 0 15530 800 6 HADDR[15]
port 8 nsew signal output
rlabel metal2 s 16394 0 16450 800 6 HADDR[16]
port 9 nsew signal output
rlabel metal2 s 17406 0 17462 800 6 HADDR[17]
port 10 nsew signal output
rlabel metal2 s 18418 0 18474 800 6 HADDR[18]
port 11 nsew signal output
rlabel metal2 s 19430 0 19486 800 6 HADDR[19]
port 12 nsew signal output
rlabel metal2 s 1398 0 1454 800 6 HADDR[1]
port 13 nsew signal output
rlabel metal2 s 20442 0 20498 800 6 HADDR[20]
port 14 nsew signal output
rlabel metal2 s 21454 0 21510 800 6 HADDR[21]
port 15 nsew signal output
rlabel metal2 s 22466 0 22522 800 6 HADDR[22]
port 16 nsew signal output
rlabel metal2 s 23386 0 23442 800 6 HADDR[23]
port 17 nsew signal output
rlabel metal2 s 24398 0 24454 800 6 HADDR[24]
port 18 nsew signal output
rlabel metal2 s 25410 0 25466 800 6 HADDR[25]
port 19 nsew signal output
rlabel metal2 s 26422 0 26478 800 6 HADDR[26]
port 20 nsew signal output
rlabel metal2 s 27434 0 27490 800 6 HADDR[27]
port 21 nsew signal output
rlabel metal2 s 28446 0 28502 800 6 HADDR[28]
port 22 nsew signal output
rlabel metal2 s 29458 0 29514 800 6 HADDR[29]
port 23 nsew signal output
rlabel metal2 s 2410 0 2466 800 6 HADDR[2]
port 24 nsew signal output
rlabel metal2 s 30470 0 30526 800 6 HADDR[30]
port 25 nsew signal output
rlabel metal2 s 31390 0 31446 800 6 HADDR[31]
port 26 nsew signal output
rlabel metal2 s 3422 0 3478 800 6 HADDR[3]
port 27 nsew signal output
rlabel metal2 s 4434 0 4490 800 6 HADDR[4]
port 28 nsew signal output
rlabel metal2 s 5446 0 5502 800 6 HADDR[5]
port 29 nsew signal output
rlabel metal2 s 6458 0 6514 800 6 HADDR[6]
port 30 nsew signal output
rlabel metal2 s 7470 0 7526 800 6 HADDR[7]
port 31 nsew signal output
rlabel metal2 s 8390 0 8446 800 6 HADDR[8]
port 32 nsew signal output
rlabel metal2 s 9402 0 9458 800 6 HADDR[9]
port 33 nsew signal output
rlabel metal3 s 0 3000 800 3120 6 HCLK
port 34 nsew signal input
rlabel metal2 s 32402 0 32458 800 6 HRDATA[0]
port 35 nsew signal input
rlabel metal2 s 42430 0 42486 800 6 HRDATA[10]
port 36 nsew signal input
rlabel metal2 s 43442 0 43498 800 6 HRDATA[11]
port 37 nsew signal input
rlabel metal2 s 44454 0 44510 800 6 HRDATA[12]
port 38 nsew signal input
rlabel metal2 s 45466 0 45522 800 6 HRDATA[13]
port 39 nsew signal input
rlabel metal2 s 46386 0 46442 800 6 HRDATA[14]
port 40 nsew signal input
rlabel metal2 s 47398 0 47454 800 6 HRDATA[15]
port 41 nsew signal input
rlabel metal2 s 48410 0 48466 800 6 HRDATA[16]
port 42 nsew signal input
rlabel metal2 s 49422 0 49478 800 6 HRDATA[17]
port 43 nsew signal input
rlabel metal2 s 50434 0 50490 800 6 HRDATA[18]
port 44 nsew signal input
rlabel metal2 s 51446 0 51502 800 6 HRDATA[19]
port 45 nsew signal input
rlabel metal2 s 33414 0 33470 800 6 HRDATA[1]
port 46 nsew signal input
rlabel metal2 s 52458 0 52514 800 6 HRDATA[20]
port 47 nsew signal input
rlabel metal2 s 53378 0 53434 800 6 HRDATA[21]
port 48 nsew signal input
rlabel metal2 s 54390 0 54446 800 6 HRDATA[22]
port 49 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 HRDATA[23]
port 50 nsew signal input
rlabel metal2 s 56414 0 56470 800 6 HRDATA[24]
port 51 nsew signal input
rlabel metal2 s 57426 0 57482 800 6 HRDATA[25]
port 52 nsew signal input
rlabel metal2 s 58438 0 58494 800 6 HRDATA[26]
port 53 nsew signal input
rlabel metal2 s 59450 0 59506 800 6 HRDATA[27]
port 54 nsew signal input
rlabel metal2 s 60462 0 60518 800 6 HRDATA[28]
port 55 nsew signal input
rlabel metal2 s 61382 0 61438 800 6 HRDATA[29]
port 56 nsew signal input
rlabel metal2 s 34426 0 34482 800 6 HRDATA[2]
port 57 nsew signal input
rlabel metal2 s 62394 0 62450 800 6 HRDATA[30]
port 58 nsew signal input
rlabel metal2 s 63406 0 63462 800 6 HRDATA[31]
port 59 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 HRDATA[3]
port 60 nsew signal input
rlabel metal2 s 36450 0 36506 800 6 HRDATA[4]
port 61 nsew signal input
rlabel metal2 s 37462 0 37518 800 6 HRDATA[5]
port 62 nsew signal input
rlabel metal2 s 38382 0 38438 800 6 HRDATA[6]
port 63 nsew signal input
rlabel metal2 s 39394 0 39450 800 6 HRDATA[7]
port 64 nsew signal input
rlabel metal2 s 40406 0 40462 800 6 HRDATA[8]
port 65 nsew signal input
rlabel metal2 s 41418 0 41474 800 6 HRDATA[9]
port 66 nsew signal input
rlabel metal3 s 0 21360 800 21480 6 HREADY
port 67 nsew signal input
rlabel metal3 s 0 9120 800 9240 6 HRESETn
port 68 nsew signal input
rlabel metal3 s 0 33736 800 33856 6 HSIZE[0]
port 69 nsew signal output
rlabel metal3 s 0 39856 800 39976 6 HSIZE[1]
port 70 nsew signal output
rlabel metal3 s 0 45976 800 46096 6 HSIZE[2]
port 71 nsew signal output
rlabel metal3 s 0 52096 800 52216 6 HTRANS[0]
port 72 nsew signal output
rlabel metal3 s 0 58352 800 58472 6 HTRANS[1]
port 73 nsew signal output
rlabel metal2 s 64418 0 64474 800 6 HWDATA[0]
port 74 nsew signal output
rlabel metal2 s 74446 0 74502 800 6 HWDATA[10]
port 75 nsew signal output
rlabel metal2 s 75458 0 75514 800 6 HWDATA[11]
port 76 nsew signal output
rlabel metal2 s 76378 0 76434 800 6 HWDATA[12]
port 77 nsew signal output
rlabel metal2 s 77390 0 77446 800 6 HWDATA[13]
port 78 nsew signal output
rlabel metal2 s 78402 0 78458 800 6 HWDATA[14]
port 79 nsew signal output
rlabel metal2 s 79414 0 79470 800 6 HWDATA[15]
port 80 nsew signal output
rlabel metal2 s 80426 0 80482 800 6 HWDATA[16]
port 81 nsew signal output
rlabel metal2 s 81438 0 81494 800 6 HWDATA[17]
port 82 nsew signal output
rlabel metal2 s 82450 0 82506 800 6 HWDATA[18]
port 83 nsew signal output
rlabel metal2 s 83370 0 83426 800 6 HWDATA[19]
port 84 nsew signal output
rlabel metal2 s 65430 0 65486 800 6 HWDATA[1]
port 85 nsew signal output
rlabel metal2 s 84382 0 84438 800 6 HWDATA[20]
port 86 nsew signal output
rlabel metal2 s 85394 0 85450 800 6 HWDATA[21]
port 87 nsew signal output
rlabel metal2 s 86406 0 86462 800 6 HWDATA[22]
port 88 nsew signal output
rlabel metal2 s 87418 0 87474 800 6 HWDATA[23]
port 89 nsew signal output
rlabel metal2 s 88430 0 88486 800 6 HWDATA[24]
port 90 nsew signal output
rlabel metal2 s 89442 0 89498 800 6 HWDATA[25]
port 91 nsew signal output
rlabel metal2 s 90454 0 90510 800 6 HWDATA[26]
port 92 nsew signal output
rlabel metal2 s 91374 0 91430 800 6 HWDATA[27]
port 93 nsew signal output
rlabel metal2 s 92386 0 92442 800 6 HWDATA[28]
port 94 nsew signal output
rlabel metal2 s 93398 0 93454 800 6 HWDATA[29]
port 95 nsew signal output
rlabel metal2 s 66442 0 66498 800 6 HWDATA[2]
port 96 nsew signal output
rlabel metal2 s 94410 0 94466 800 6 HWDATA[30]
port 97 nsew signal output
rlabel metal2 s 95422 0 95478 800 6 HWDATA[31]
port 98 nsew signal output
rlabel metal2 s 67454 0 67510 800 6 HWDATA[3]
port 99 nsew signal output
rlabel metal2 s 68374 0 68430 800 6 HWDATA[4]
port 100 nsew signal output
rlabel metal2 s 69386 0 69442 800 6 HWDATA[5]
port 101 nsew signal output
rlabel metal2 s 70398 0 70454 800 6 HWDATA[6]
port 102 nsew signal output
rlabel metal2 s 71410 0 71466 800 6 HWDATA[7]
port 103 nsew signal output
rlabel metal2 s 72422 0 72478 800 6 HWDATA[8]
port 104 nsew signal output
rlabel metal2 s 73434 0 73490 800 6 HWDATA[9]
port 105 nsew signal output
rlabel metal3 s 0 15240 800 15360 6 HWRITE
port 106 nsew signal output
rlabel metal3 s 0 64472 800 64592 6 IRQ[0]
port 107 nsew signal input
rlabel metal3 s 0 125944 800 126064 6 IRQ[10]
port 108 nsew signal input
rlabel metal3 s 0 132064 800 132184 6 IRQ[11]
port 109 nsew signal input
rlabel metal3 s 0 138320 800 138440 6 IRQ[12]
port 110 nsew signal input
rlabel metal3 s 0 144440 800 144560 6 IRQ[13]
port 111 nsew signal input
rlabel metal3 s 0 150560 800 150680 6 IRQ[14]
port 112 nsew signal input
rlabel metal3 s 0 70592 800 70712 6 IRQ[1]
port 113 nsew signal input
rlabel metal3 s 0 76712 800 76832 6 IRQ[2]
port 114 nsew signal input
rlabel metal3 s 0 82968 800 83088 6 IRQ[3]
port 115 nsew signal input
rlabel metal3 s 0 89088 800 89208 6 IRQ[4]
port 116 nsew signal input
rlabel metal3 s 0 95208 800 95328 6 IRQ[5]
port 117 nsew signal input
rlabel metal3 s 0 101328 800 101448 6 IRQ[6]
port 118 nsew signal input
rlabel metal3 s 0 107448 800 107568 6 IRQ[7]
port 119 nsew signal input
rlabel metal3 s 0 113704 800 113824 6 IRQ[8]
port 120 nsew signal input
rlabel metal3 s 0 119824 800 119944 6 IRQ[9]
port 121 nsew signal input
rlabel metal3 s 0 27480 800 27600 6 NMI
port 122 nsew signal input
rlabel metal2 s 96434 0 96490 800 6 SYSTICKCLKDIV[0]
port 123 nsew signal input
rlabel metal2 s 106370 0 106426 800 6 SYSTICKCLKDIV[10]
port 124 nsew signal input
rlabel metal2 s 107382 0 107438 800 6 SYSTICKCLKDIV[11]
port 125 nsew signal input
rlabel metal2 s 108394 0 108450 800 6 SYSTICKCLKDIV[12]
port 126 nsew signal input
rlabel metal2 s 109406 0 109462 800 6 SYSTICKCLKDIV[13]
port 127 nsew signal input
rlabel metal2 s 110418 0 110474 800 6 SYSTICKCLKDIV[14]
port 128 nsew signal input
rlabel metal2 s 111430 0 111486 800 6 SYSTICKCLKDIV[15]
port 129 nsew signal input
rlabel metal2 s 112442 0 112498 800 6 SYSTICKCLKDIV[16]
port 130 nsew signal input
rlabel metal2 s 113362 0 113418 800 6 SYSTICKCLKDIV[17]
port 131 nsew signal input
rlabel metal2 s 114374 0 114430 800 6 SYSTICKCLKDIV[18]
port 132 nsew signal input
rlabel metal2 s 115386 0 115442 800 6 SYSTICKCLKDIV[19]
port 133 nsew signal input
rlabel metal2 s 97446 0 97502 800 6 SYSTICKCLKDIV[1]
port 134 nsew signal input
rlabel metal2 s 116398 0 116454 800 6 SYSTICKCLKDIV[20]
port 135 nsew signal input
rlabel metal2 s 117410 0 117466 800 6 SYSTICKCLKDIV[21]
port 136 nsew signal input
rlabel metal2 s 118422 0 118478 800 6 SYSTICKCLKDIV[22]
port 137 nsew signal input
rlabel metal2 s 119434 0 119490 800 6 SYSTICKCLKDIV[23]
port 138 nsew signal input
rlabel metal2 s 98366 0 98422 800 6 SYSTICKCLKDIV[2]
port 139 nsew signal input
rlabel metal2 s 99378 0 99434 800 6 SYSTICKCLKDIV[3]
port 140 nsew signal input
rlabel metal2 s 100390 0 100446 800 6 SYSTICKCLKDIV[4]
port 141 nsew signal input
rlabel metal2 s 101402 0 101458 800 6 SYSTICKCLKDIV[5]
port 142 nsew signal input
rlabel metal2 s 102414 0 102470 800 6 SYSTICKCLKDIV[6]
port 143 nsew signal input
rlabel metal2 s 103426 0 103482 800 6 SYSTICKCLKDIV[7]
port 144 nsew signal input
rlabel metal2 s 104438 0 104494 800 6 SYSTICKCLKDIV[8]
port 145 nsew signal input
rlabel metal2 s 105450 0 105506 800 6 SYSTICKCLKDIV[9]
port 146 nsew signal input
rlabel metal4 s 96368 2128 96688 157808 6 vccd1
port 147 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 157808 6 vccd1
port 148 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 157808 6 vccd1
port 149 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 157808 6 vccd1
port 150 nsew power bidirectional
rlabel metal4 s 111728 2128 112048 157808 6 vssd1
port 151 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 157808 6 vssd1
port 152 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 157808 6 vssd1
port 153 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 157808 6 vssd1
port 154 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 120000 160000
string LEFview TRUE
string GDS_FILE ../gds/apb_sys_0.gds
string GDS_END 51979460
string GDS_START 1299454
<< end >>

