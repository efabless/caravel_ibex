magic
tech sky130A
magscale 1 2
timestamp 1617742078
<< obsli1 >>
rect 1104 2159 79183 117521
<< obsm1 >>
rect 1104 1300 79195 117552
<< metal2 >>
rect 478 119200 534 120000
rect 1398 119200 1454 120000
rect 2410 119200 2466 120000
rect 3422 119200 3478 120000
rect 4434 119200 4490 120000
rect 5446 119200 5502 120000
rect 6458 119200 6514 120000
rect 7470 119200 7526 120000
rect 8482 119200 8538 120000
rect 9402 119200 9458 120000
rect 10414 119200 10470 120000
rect 11426 119200 11482 120000
rect 12438 119200 12494 120000
rect 13450 119200 13506 120000
rect 14462 119200 14518 120000
rect 15474 119200 15530 120000
rect 16486 119200 16542 120000
rect 17406 119200 17462 120000
rect 18418 119200 18474 120000
rect 19430 119200 19486 120000
rect 20442 119200 20498 120000
rect 21454 119200 21510 120000
rect 22466 119200 22522 120000
rect 23478 119200 23534 120000
rect 24490 119200 24546 120000
rect 25410 119200 25466 120000
rect 26422 119200 26478 120000
rect 27434 119200 27490 120000
rect 28446 119200 28502 120000
rect 29458 119200 29514 120000
rect 30470 119200 30526 120000
rect 31482 119200 31538 120000
rect 32494 119200 32550 120000
rect 33414 119200 33470 120000
rect 34426 119200 34482 120000
rect 35438 119200 35494 120000
rect 36450 119200 36506 120000
rect 37462 119200 37518 120000
rect 38474 119200 38530 120000
rect 39486 119200 39542 120000
rect 40498 119200 40554 120000
rect 41418 119200 41474 120000
rect 42430 119200 42486 120000
rect 43442 119200 43498 120000
rect 44454 119200 44510 120000
rect 45466 119200 45522 120000
rect 46478 119200 46534 120000
rect 47490 119200 47546 120000
rect 48502 119200 48558 120000
rect 49422 119200 49478 120000
rect 50434 119200 50490 120000
rect 51446 119200 51502 120000
rect 52458 119200 52514 120000
rect 53470 119200 53526 120000
rect 54482 119200 54538 120000
rect 55494 119200 55550 120000
rect 56506 119200 56562 120000
rect 57426 119200 57482 120000
rect 58438 119200 58494 120000
rect 59450 119200 59506 120000
rect 60462 119200 60518 120000
rect 61474 119200 61530 120000
rect 62486 119200 62542 120000
rect 63498 119200 63554 120000
rect 64510 119200 64566 120000
rect 65430 119200 65486 120000
rect 66442 119200 66498 120000
rect 67454 119200 67510 120000
rect 68466 119200 68522 120000
rect 69478 119200 69534 120000
rect 70490 119200 70546 120000
rect 71502 119200 71558 120000
rect 72514 119200 72570 120000
rect 73434 119200 73490 120000
rect 74446 119200 74502 120000
rect 75458 119200 75514 120000
rect 76470 119200 76526 120000
rect 77482 119200 77538 120000
rect 78494 119200 78550 120000
rect 79506 119200 79562 120000
rect 9954 0 10010 800
rect 29918 0 29974 800
rect 49974 0 50030 800
rect 69938 0 69994 800
<< obsm2 >>
rect 1510 119144 2354 119513
rect 2522 119144 3366 119513
rect 3534 119144 4378 119513
rect 4546 119144 5390 119513
rect 5558 119144 6402 119513
rect 6570 119144 7414 119513
rect 7582 119144 8426 119513
rect 8594 119144 9346 119513
rect 9514 119144 10358 119513
rect 10526 119144 11370 119513
rect 11538 119144 12382 119513
rect 12550 119144 13394 119513
rect 13562 119144 14406 119513
rect 14574 119144 15418 119513
rect 15586 119144 16430 119513
rect 16598 119144 17350 119513
rect 17518 119144 18362 119513
rect 18530 119144 19374 119513
rect 19542 119144 20386 119513
rect 20554 119144 21398 119513
rect 21566 119144 22410 119513
rect 22578 119144 23422 119513
rect 23590 119144 24434 119513
rect 24602 119144 25354 119513
rect 25522 119144 26366 119513
rect 26534 119144 27378 119513
rect 27546 119144 28390 119513
rect 28558 119144 29402 119513
rect 29570 119144 30414 119513
rect 30582 119144 31426 119513
rect 31594 119144 32438 119513
rect 32606 119144 33358 119513
rect 33526 119144 34370 119513
rect 34538 119144 35382 119513
rect 35550 119144 36394 119513
rect 36562 119144 37406 119513
rect 37574 119144 38418 119513
rect 38586 119144 39430 119513
rect 39598 119144 40442 119513
rect 40610 119144 41362 119513
rect 41530 119144 42374 119513
rect 42542 119144 43386 119513
rect 43554 119144 44398 119513
rect 44566 119144 45410 119513
rect 45578 119144 46422 119513
rect 46590 119144 47434 119513
rect 47602 119144 48446 119513
rect 48614 119144 49366 119513
rect 49534 119144 50378 119513
rect 50546 119144 51390 119513
rect 51558 119144 52402 119513
rect 52570 119144 53414 119513
rect 53582 119144 54426 119513
rect 54594 119144 55438 119513
rect 55606 119144 56450 119513
rect 56618 119144 57370 119513
rect 57538 119144 58382 119513
rect 58550 119144 59394 119513
rect 59562 119144 60406 119513
rect 60574 119144 61418 119513
rect 61586 119144 62430 119513
rect 62598 119144 63442 119513
rect 63610 119144 64454 119513
rect 64622 119144 65374 119513
rect 65542 119144 66386 119513
rect 66554 119144 67398 119513
rect 67566 119144 68410 119513
rect 68578 119144 69422 119513
rect 69590 119144 70434 119513
rect 70602 119144 71446 119513
rect 71614 119144 72458 119513
rect 72626 119144 73378 119513
rect 73546 119144 74390 119513
rect 74558 119144 75402 119513
rect 75570 119144 76414 119513
rect 76582 119144 77426 119513
rect 77594 119144 78438 119513
rect 78606 119144 79450 119513
rect 1398 856 79562 119144
rect 1398 439 9898 856
rect 10066 439 29862 856
rect 30030 439 49918 856
rect 50086 439 69882 856
rect 70050 439 79562 856
<< metal3 >>
rect 79200 119416 80000 119536
rect 79200 118464 80000 118584
rect 79200 117512 80000 117632
rect 79200 116560 80000 116680
rect 79200 115608 80000 115728
rect 79200 114656 80000 114776
rect 79200 113704 80000 113824
rect 79200 112752 80000 112872
rect 79200 111800 80000 111920
rect 79200 110984 80000 111104
rect 79200 110032 80000 110152
rect 79200 109080 80000 109200
rect 79200 108128 80000 108248
rect 79200 107176 80000 107296
rect 79200 106224 80000 106344
rect 79200 105272 80000 105392
rect 79200 104320 80000 104440
rect 79200 103368 80000 103488
rect 79200 102552 80000 102672
rect 79200 101600 80000 101720
rect 79200 100648 80000 100768
rect 79200 99696 80000 99816
rect 79200 98744 80000 98864
rect 79200 97792 80000 97912
rect 79200 96840 80000 96960
rect 79200 95888 80000 96008
rect 79200 94936 80000 95056
rect 79200 94120 80000 94240
rect 79200 93168 80000 93288
rect 79200 92216 80000 92336
rect 79200 91264 80000 91384
rect 79200 90312 80000 90432
rect 79200 89360 80000 89480
rect 79200 88408 80000 88528
rect 79200 87456 80000 87576
rect 79200 86504 80000 86624
rect 79200 85688 80000 85808
rect 79200 84736 80000 84856
rect 79200 83784 80000 83904
rect 79200 82832 80000 82952
rect 79200 81880 80000 82000
rect 79200 80928 80000 81048
rect 79200 79976 80000 80096
rect 79200 79024 80000 79144
rect 79200 78072 80000 78192
rect 79200 77256 80000 77376
rect 79200 76304 80000 76424
rect 79200 75352 80000 75472
rect 79200 74400 80000 74520
rect 79200 73448 80000 73568
rect 79200 72496 80000 72616
rect 79200 71544 80000 71664
rect 79200 70592 80000 70712
rect 79200 69640 80000 69760
rect 79200 68824 80000 68944
rect 79200 67872 80000 67992
rect 79200 66920 80000 67040
rect 79200 65968 80000 66088
rect 79200 65016 80000 65136
rect 79200 64064 80000 64184
rect 79200 63112 80000 63232
rect 79200 62160 80000 62280
rect 79200 61208 80000 61328
rect 79200 60392 80000 60512
rect 79200 59440 80000 59560
rect 79200 58488 80000 58608
rect 79200 57536 80000 57656
rect 79200 56584 80000 56704
rect 79200 55632 80000 55752
rect 79200 54680 80000 54800
rect 79200 53728 80000 53848
rect 79200 52776 80000 52896
rect 79200 51824 80000 51944
rect 79200 51008 80000 51128
rect 79200 50056 80000 50176
rect 79200 49104 80000 49224
rect 79200 48152 80000 48272
rect 79200 47200 80000 47320
rect 79200 46248 80000 46368
rect 79200 45296 80000 45416
rect 79200 44344 80000 44464
rect 79200 43392 80000 43512
rect 79200 42576 80000 42696
rect 79200 41624 80000 41744
rect 79200 40672 80000 40792
rect 79200 39720 80000 39840
rect 79200 38768 80000 38888
rect 79200 37816 80000 37936
rect 79200 36864 80000 36984
rect 79200 35912 80000 36032
rect 79200 34960 80000 35080
rect 79200 34144 80000 34264
rect 79200 33192 80000 33312
rect 79200 32240 80000 32360
rect 79200 31288 80000 31408
rect 79200 30336 80000 30456
rect 79200 29384 80000 29504
rect 79200 28432 80000 28552
rect 79200 27480 80000 27600
rect 79200 26528 80000 26648
rect 79200 25712 80000 25832
rect 79200 24760 80000 24880
rect 79200 23808 80000 23928
rect 79200 22856 80000 22976
rect 79200 21904 80000 22024
rect 79200 20952 80000 21072
rect 79200 20000 80000 20120
rect 79200 19048 80000 19168
rect 79200 18096 80000 18216
rect 79200 17280 80000 17400
rect 79200 16328 80000 16448
rect 79200 15376 80000 15496
rect 79200 14424 80000 14544
rect 79200 13472 80000 13592
rect 79200 12520 80000 12640
rect 79200 11568 80000 11688
rect 79200 10616 80000 10736
rect 79200 9664 80000 9784
rect 79200 8848 80000 8968
rect 79200 7896 80000 8016
rect 79200 6944 80000 7064
rect 79200 5992 80000 6112
rect 79200 5040 80000 5160
rect 79200 4088 80000 4208
rect 79200 3136 80000 3256
rect 79200 2184 80000 2304
rect 79200 1232 80000 1352
rect 79200 416 80000 536
<< obsm3 >>
rect 1393 119336 79120 119509
rect 1393 118664 79567 119336
rect 1393 118384 79120 118664
rect 1393 117712 79567 118384
rect 1393 117432 79120 117712
rect 1393 116760 79567 117432
rect 1393 116480 79120 116760
rect 1393 115808 79567 116480
rect 1393 115528 79120 115808
rect 1393 114856 79567 115528
rect 1393 114576 79120 114856
rect 1393 113904 79567 114576
rect 1393 113624 79120 113904
rect 1393 112952 79567 113624
rect 1393 112672 79120 112952
rect 1393 112000 79567 112672
rect 1393 111720 79120 112000
rect 1393 111184 79567 111720
rect 1393 110904 79120 111184
rect 1393 110232 79567 110904
rect 1393 109952 79120 110232
rect 1393 109280 79567 109952
rect 1393 109000 79120 109280
rect 1393 108328 79567 109000
rect 1393 108048 79120 108328
rect 1393 107376 79567 108048
rect 1393 107096 79120 107376
rect 1393 106424 79567 107096
rect 1393 106144 79120 106424
rect 1393 105472 79567 106144
rect 1393 105192 79120 105472
rect 1393 104520 79567 105192
rect 1393 104240 79120 104520
rect 1393 103568 79567 104240
rect 1393 103288 79120 103568
rect 1393 102752 79567 103288
rect 1393 102472 79120 102752
rect 1393 101800 79567 102472
rect 1393 101520 79120 101800
rect 1393 100848 79567 101520
rect 1393 100568 79120 100848
rect 1393 99896 79567 100568
rect 1393 99616 79120 99896
rect 1393 98944 79567 99616
rect 1393 98664 79120 98944
rect 1393 97992 79567 98664
rect 1393 97712 79120 97992
rect 1393 97040 79567 97712
rect 1393 96760 79120 97040
rect 1393 96088 79567 96760
rect 1393 95808 79120 96088
rect 1393 95136 79567 95808
rect 1393 94856 79120 95136
rect 1393 94320 79567 94856
rect 1393 94040 79120 94320
rect 1393 93368 79567 94040
rect 1393 93088 79120 93368
rect 1393 92416 79567 93088
rect 1393 92136 79120 92416
rect 1393 91464 79567 92136
rect 1393 91184 79120 91464
rect 1393 90512 79567 91184
rect 1393 90232 79120 90512
rect 1393 89560 79567 90232
rect 1393 89280 79120 89560
rect 1393 88608 79567 89280
rect 1393 88328 79120 88608
rect 1393 87656 79567 88328
rect 1393 87376 79120 87656
rect 1393 86704 79567 87376
rect 1393 86424 79120 86704
rect 1393 85888 79567 86424
rect 1393 85608 79120 85888
rect 1393 84936 79567 85608
rect 1393 84656 79120 84936
rect 1393 83984 79567 84656
rect 1393 83704 79120 83984
rect 1393 83032 79567 83704
rect 1393 82752 79120 83032
rect 1393 82080 79567 82752
rect 1393 81800 79120 82080
rect 1393 81128 79567 81800
rect 1393 80848 79120 81128
rect 1393 80176 79567 80848
rect 1393 79896 79120 80176
rect 1393 79224 79567 79896
rect 1393 78944 79120 79224
rect 1393 78272 79567 78944
rect 1393 77992 79120 78272
rect 1393 77456 79567 77992
rect 1393 77176 79120 77456
rect 1393 76504 79567 77176
rect 1393 76224 79120 76504
rect 1393 75552 79567 76224
rect 1393 75272 79120 75552
rect 1393 74600 79567 75272
rect 1393 74320 79120 74600
rect 1393 73648 79567 74320
rect 1393 73368 79120 73648
rect 1393 72696 79567 73368
rect 1393 72416 79120 72696
rect 1393 71744 79567 72416
rect 1393 71464 79120 71744
rect 1393 70792 79567 71464
rect 1393 70512 79120 70792
rect 1393 69840 79567 70512
rect 1393 69560 79120 69840
rect 1393 69024 79567 69560
rect 1393 68744 79120 69024
rect 1393 68072 79567 68744
rect 1393 67792 79120 68072
rect 1393 67120 79567 67792
rect 1393 66840 79120 67120
rect 1393 66168 79567 66840
rect 1393 65888 79120 66168
rect 1393 65216 79567 65888
rect 1393 64936 79120 65216
rect 1393 64264 79567 64936
rect 1393 63984 79120 64264
rect 1393 63312 79567 63984
rect 1393 63032 79120 63312
rect 1393 62360 79567 63032
rect 1393 62080 79120 62360
rect 1393 61408 79567 62080
rect 1393 61128 79120 61408
rect 1393 60592 79567 61128
rect 1393 60312 79120 60592
rect 1393 59640 79567 60312
rect 1393 59360 79120 59640
rect 1393 58688 79567 59360
rect 1393 58408 79120 58688
rect 1393 57736 79567 58408
rect 1393 57456 79120 57736
rect 1393 56784 79567 57456
rect 1393 56504 79120 56784
rect 1393 55832 79567 56504
rect 1393 55552 79120 55832
rect 1393 54880 79567 55552
rect 1393 54600 79120 54880
rect 1393 53928 79567 54600
rect 1393 53648 79120 53928
rect 1393 52976 79567 53648
rect 1393 52696 79120 52976
rect 1393 52024 79567 52696
rect 1393 51744 79120 52024
rect 1393 51208 79567 51744
rect 1393 50928 79120 51208
rect 1393 50256 79567 50928
rect 1393 49976 79120 50256
rect 1393 49304 79567 49976
rect 1393 49024 79120 49304
rect 1393 48352 79567 49024
rect 1393 48072 79120 48352
rect 1393 47400 79567 48072
rect 1393 47120 79120 47400
rect 1393 46448 79567 47120
rect 1393 46168 79120 46448
rect 1393 45496 79567 46168
rect 1393 45216 79120 45496
rect 1393 44544 79567 45216
rect 1393 44264 79120 44544
rect 1393 43592 79567 44264
rect 1393 43312 79120 43592
rect 1393 42776 79567 43312
rect 1393 42496 79120 42776
rect 1393 41824 79567 42496
rect 1393 41544 79120 41824
rect 1393 40872 79567 41544
rect 1393 40592 79120 40872
rect 1393 39920 79567 40592
rect 1393 39640 79120 39920
rect 1393 38968 79567 39640
rect 1393 38688 79120 38968
rect 1393 38016 79567 38688
rect 1393 37736 79120 38016
rect 1393 37064 79567 37736
rect 1393 36784 79120 37064
rect 1393 36112 79567 36784
rect 1393 35832 79120 36112
rect 1393 35160 79567 35832
rect 1393 34880 79120 35160
rect 1393 34344 79567 34880
rect 1393 34064 79120 34344
rect 1393 33392 79567 34064
rect 1393 33112 79120 33392
rect 1393 32440 79567 33112
rect 1393 32160 79120 32440
rect 1393 31488 79567 32160
rect 1393 31208 79120 31488
rect 1393 30536 79567 31208
rect 1393 30256 79120 30536
rect 1393 29584 79567 30256
rect 1393 29304 79120 29584
rect 1393 28632 79567 29304
rect 1393 28352 79120 28632
rect 1393 27680 79567 28352
rect 1393 27400 79120 27680
rect 1393 26728 79567 27400
rect 1393 26448 79120 26728
rect 1393 25912 79567 26448
rect 1393 25632 79120 25912
rect 1393 24960 79567 25632
rect 1393 24680 79120 24960
rect 1393 24008 79567 24680
rect 1393 23728 79120 24008
rect 1393 23056 79567 23728
rect 1393 22776 79120 23056
rect 1393 22104 79567 22776
rect 1393 21824 79120 22104
rect 1393 21152 79567 21824
rect 1393 20872 79120 21152
rect 1393 20200 79567 20872
rect 1393 19920 79120 20200
rect 1393 19248 79567 19920
rect 1393 18968 79120 19248
rect 1393 18296 79567 18968
rect 1393 18016 79120 18296
rect 1393 17480 79567 18016
rect 1393 17200 79120 17480
rect 1393 16528 79567 17200
rect 1393 16248 79120 16528
rect 1393 15576 79567 16248
rect 1393 15296 79120 15576
rect 1393 14624 79567 15296
rect 1393 14344 79120 14624
rect 1393 13672 79567 14344
rect 1393 13392 79120 13672
rect 1393 12720 79567 13392
rect 1393 12440 79120 12720
rect 1393 11768 79567 12440
rect 1393 11488 79120 11768
rect 1393 10816 79567 11488
rect 1393 10536 79120 10816
rect 1393 9864 79567 10536
rect 1393 9584 79120 9864
rect 1393 9048 79567 9584
rect 1393 8768 79120 9048
rect 1393 8096 79567 8768
rect 1393 7816 79120 8096
rect 1393 7144 79567 7816
rect 1393 6864 79120 7144
rect 1393 6192 79567 6864
rect 1393 5912 79120 6192
rect 1393 5240 79567 5912
rect 1393 4960 79120 5240
rect 1393 4288 79567 4960
rect 1393 4008 79120 4288
rect 1393 3336 79567 4008
rect 1393 3056 79120 3336
rect 1393 2384 79567 3056
rect 1393 2104 79120 2384
rect 1393 1432 79567 2104
rect 1393 1152 79120 1432
rect 1393 616 79567 1152
rect 1393 443 79120 616
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
<< obsm4 >>
rect 8155 6155 19488 117061
rect 19968 6155 34848 117061
rect 35328 6155 50208 117061
rect 50688 6155 65568 117061
rect 66048 6155 73725 117061
<< labels >>
rlabel metal2 s 478 119200 534 120000 6 A[0]
port 1 nsew signal input
rlabel metal2 s 10414 119200 10470 120000 6 A[10]
port 2 nsew signal input
rlabel metal2 s 11426 119200 11482 120000 6 A[11]
port 3 nsew signal input
rlabel metal2 s 12438 119200 12494 120000 6 A[12]
port 4 nsew signal input
rlabel metal2 s 13450 119200 13506 120000 6 A[13]
port 5 nsew signal input
rlabel metal2 s 14462 119200 14518 120000 6 A[14]
port 6 nsew signal input
rlabel metal2 s 15474 119200 15530 120000 6 A[15]
port 7 nsew signal input
rlabel metal2 s 16486 119200 16542 120000 6 A[16]
port 8 nsew signal input
rlabel metal2 s 17406 119200 17462 120000 6 A[17]
port 9 nsew signal input
rlabel metal2 s 18418 119200 18474 120000 6 A[18]
port 10 nsew signal input
rlabel metal2 s 19430 119200 19486 120000 6 A[19]
port 11 nsew signal input
rlabel metal2 s 1398 119200 1454 120000 6 A[1]
port 12 nsew signal input
rlabel metal2 s 20442 119200 20498 120000 6 A[20]
port 13 nsew signal input
rlabel metal2 s 21454 119200 21510 120000 6 A[21]
port 14 nsew signal input
rlabel metal2 s 22466 119200 22522 120000 6 A[22]
port 15 nsew signal input
rlabel metal2 s 23478 119200 23534 120000 6 A[23]
port 16 nsew signal input
rlabel metal2 s 2410 119200 2466 120000 6 A[2]
port 17 nsew signal input
rlabel metal2 s 3422 119200 3478 120000 6 A[3]
port 18 nsew signal input
rlabel metal2 s 4434 119200 4490 120000 6 A[4]
port 19 nsew signal input
rlabel metal2 s 5446 119200 5502 120000 6 A[5]
port 20 nsew signal input
rlabel metal2 s 6458 119200 6514 120000 6 A[6]
port 21 nsew signal input
rlabel metal2 s 7470 119200 7526 120000 6 A[7]
port 22 nsew signal input
rlabel metal2 s 8482 119200 8538 120000 6 A[8]
port 23 nsew signal input
rlabel metal2 s 9402 119200 9458 120000 6 A[9]
port 24 nsew signal input
rlabel metal2 s 24490 119200 24546 120000 6 A_h[0]
port 25 nsew signal input
rlabel metal2 s 34426 119200 34482 120000 6 A_h[10]
port 26 nsew signal input
rlabel metal2 s 35438 119200 35494 120000 6 A_h[11]
port 27 nsew signal input
rlabel metal2 s 36450 119200 36506 120000 6 A_h[12]
port 28 nsew signal input
rlabel metal2 s 37462 119200 37518 120000 6 A_h[13]
port 29 nsew signal input
rlabel metal2 s 38474 119200 38530 120000 6 A_h[14]
port 30 nsew signal input
rlabel metal2 s 39486 119200 39542 120000 6 A_h[15]
port 31 nsew signal input
rlabel metal2 s 40498 119200 40554 120000 6 A_h[16]
port 32 nsew signal input
rlabel metal2 s 41418 119200 41474 120000 6 A_h[17]
port 33 nsew signal input
rlabel metal2 s 42430 119200 42486 120000 6 A_h[18]
port 34 nsew signal input
rlabel metal2 s 43442 119200 43498 120000 6 A_h[19]
port 35 nsew signal input
rlabel metal2 s 25410 119200 25466 120000 6 A_h[1]
port 36 nsew signal input
rlabel metal2 s 44454 119200 44510 120000 6 A_h[20]
port 37 nsew signal input
rlabel metal2 s 45466 119200 45522 120000 6 A_h[21]
port 38 nsew signal input
rlabel metal2 s 46478 119200 46534 120000 6 A_h[22]
port 39 nsew signal input
rlabel metal2 s 47490 119200 47546 120000 6 A_h[23]
port 40 nsew signal input
rlabel metal2 s 26422 119200 26478 120000 6 A_h[2]
port 41 nsew signal input
rlabel metal2 s 27434 119200 27490 120000 6 A_h[3]
port 42 nsew signal input
rlabel metal2 s 28446 119200 28502 120000 6 A_h[4]
port 43 nsew signal input
rlabel metal2 s 29458 119200 29514 120000 6 A_h[5]
port 44 nsew signal input
rlabel metal2 s 30470 119200 30526 120000 6 A_h[6]
port 45 nsew signal input
rlabel metal2 s 31482 119200 31538 120000 6 A_h[7]
port 46 nsew signal input
rlabel metal2 s 32494 119200 32550 120000 6 A_h[8]
port 47 nsew signal input
rlabel metal2 s 33414 119200 33470 120000 6 A_h[9]
port 48 nsew signal input
rlabel metal2 s 48502 119200 48558 120000 6 Do[0]
port 49 nsew signal output
rlabel metal2 s 58438 119200 58494 120000 6 Do[10]
port 50 nsew signal output
rlabel metal2 s 59450 119200 59506 120000 6 Do[11]
port 51 nsew signal output
rlabel metal2 s 60462 119200 60518 120000 6 Do[12]
port 52 nsew signal output
rlabel metal2 s 61474 119200 61530 120000 6 Do[13]
port 53 nsew signal output
rlabel metal2 s 62486 119200 62542 120000 6 Do[14]
port 54 nsew signal output
rlabel metal2 s 63498 119200 63554 120000 6 Do[15]
port 55 nsew signal output
rlabel metal2 s 64510 119200 64566 120000 6 Do[16]
port 56 nsew signal output
rlabel metal2 s 65430 119200 65486 120000 6 Do[17]
port 57 nsew signal output
rlabel metal2 s 66442 119200 66498 120000 6 Do[18]
port 58 nsew signal output
rlabel metal2 s 67454 119200 67510 120000 6 Do[19]
port 59 nsew signal output
rlabel metal2 s 49422 119200 49478 120000 6 Do[1]
port 60 nsew signal output
rlabel metal2 s 68466 119200 68522 120000 6 Do[20]
port 61 nsew signal output
rlabel metal2 s 69478 119200 69534 120000 6 Do[21]
port 62 nsew signal output
rlabel metal2 s 70490 119200 70546 120000 6 Do[22]
port 63 nsew signal output
rlabel metal2 s 71502 119200 71558 120000 6 Do[23]
port 64 nsew signal output
rlabel metal2 s 72514 119200 72570 120000 6 Do[24]
port 65 nsew signal output
rlabel metal2 s 73434 119200 73490 120000 6 Do[25]
port 66 nsew signal output
rlabel metal2 s 74446 119200 74502 120000 6 Do[26]
port 67 nsew signal output
rlabel metal2 s 75458 119200 75514 120000 6 Do[27]
port 68 nsew signal output
rlabel metal2 s 76470 119200 76526 120000 6 Do[28]
port 69 nsew signal output
rlabel metal2 s 77482 119200 77538 120000 6 Do[29]
port 70 nsew signal output
rlabel metal2 s 50434 119200 50490 120000 6 Do[2]
port 71 nsew signal output
rlabel metal2 s 78494 119200 78550 120000 6 Do[30]
port 72 nsew signal output
rlabel metal2 s 79506 119200 79562 120000 6 Do[31]
port 73 nsew signal output
rlabel metal2 s 51446 119200 51502 120000 6 Do[3]
port 74 nsew signal output
rlabel metal2 s 52458 119200 52514 120000 6 Do[4]
port 75 nsew signal output
rlabel metal2 s 53470 119200 53526 120000 6 Do[5]
port 76 nsew signal output
rlabel metal2 s 54482 119200 54538 120000 6 Do[6]
port 77 nsew signal output
rlabel metal2 s 55494 119200 55550 120000 6 Do[7]
port 78 nsew signal output
rlabel metal2 s 56506 119200 56562 120000 6 Do[8]
port 79 nsew signal output
rlabel metal2 s 57426 119200 57482 120000 6 Do[9]
port 80 nsew signal output
rlabel metal2 s 9954 0 10010 800 6 clk
port 81 nsew signal input
rlabel metal2 s 69938 0 69994 800 6 hit
port 82 nsew signal output
rlabel metal3 s 79200 416 80000 536 6 line[0]
port 83 nsew signal input
rlabel metal3 s 79200 94120 80000 94240 6 line[100]
port 84 nsew signal input
rlabel metal3 s 79200 94936 80000 95056 6 line[101]
port 85 nsew signal input
rlabel metal3 s 79200 95888 80000 96008 6 line[102]
port 86 nsew signal input
rlabel metal3 s 79200 96840 80000 96960 6 line[103]
port 87 nsew signal input
rlabel metal3 s 79200 97792 80000 97912 6 line[104]
port 88 nsew signal input
rlabel metal3 s 79200 98744 80000 98864 6 line[105]
port 89 nsew signal input
rlabel metal3 s 79200 99696 80000 99816 6 line[106]
port 90 nsew signal input
rlabel metal3 s 79200 100648 80000 100768 6 line[107]
port 91 nsew signal input
rlabel metal3 s 79200 101600 80000 101720 6 line[108]
port 92 nsew signal input
rlabel metal3 s 79200 102552 80000 102672 6 line[109]
port 93 nsew signal input
rlabel metal3 s 79200 9664 80000 9784 6 line[10]
port 94 nsew signal input
rlabel metal3 s 79200 103368 80000 103488 6 line[110]
port 95 nsew signal input
rlabel metal3 s 79200 104320 80000 104440 6 line[111]
port 96 nsew signal input
rlabel metal3 s 79200 105272 80000 105392 6 line[112]
port 97 nsew signal input
rlabel metal3 s 79200 106224 80000 106344 6 line[113]
port 98 nsew signal input
rlabel metal3 s 79200 107176 80000 107296 6 line[114]
port 99 nsew signal input
rlabel metal3 s 79200 108128 80000 108248 6 line[115]
port 100 nsew signal input
rlabel metal3 s 79200 109080 80000 109200 6 line[116]
port 101 nsew signal input
rlabel metal3 s 79200 110032 80000 110152 6 line[117]
port 102 nsew signal input
rlabel metal3 s 79200 110984 80000 111104 6 line[118]
port 103 nsew signal input
rlabel metal3 s 79200 111800 80000 111920 6 line[119]
port 104 nsew signal input
rlabel metal3 s 79200 10616 80000 10736 6 line[11]
port 105 nsew signal input
rlabel metal3 s 79200 112752 80000 112872 6 line[120]
port 106 nsew signal input
rlabel metal3 s 79200 113704 80000 113824 6 line[121]
port 107 nsew signal input
rlabel metal3 s 79200 114656 80000 114776 6 line[122]
port 108 nsew signal input
rlabel metal3 s 79200 115608 80000 115728 6 line[123]
port 109 nsew signal input
rlabel metal3 s 79200 116560 80000 116680 6 line[124]
port 110 nsew signal input
rlabel metal3 s 79200 117512 80000 117632 6 line[125]
port 111 nsew signal input
rlabel metal3 s 79200 118464 80000 118584 6 line[126]
port 112 nsew signal input
rlabel metal3 s 79200 119416 80000 119536 6 line[127]
port 113 nsew signal input
rlabel metal3 s 79200 11568 80000 11688 6 line[12]
port 114 nsew signal input
rlabel metal3 s 79200 12520 80000 12640 6 line[13]
port 115 nsew signal input
rlabel metal3 s 79200 13472 80000 13592 6 line[14]
port 116 nsew signal input
rlabel metal3 s 79200 14424 80000 14544 6 line[15]
port 117 nsew signal input
rlabel metal3 s 79200 15376 80000 15496 6 line[16]
port 118 nsew signal input
rlabel metal3 s 79200 16328 80000 16448 6 line[17]
port 119 nsew signal input
rlabel metal3 s 79200 17280 80000 17400 6 line[18]
port 120 nsew signal input
rlabel metal3 s 79200 18096 80000 18216 6 line[19]
port 121 nsew signal input
rlabel metal3 s 79200 1232 80000 1352 6 line[1]
port 122 nsew signal input
rlabel metal3 s 79200 19048 80000 19168 6 line[20]
port 123 nsew signal input
rlabel metal3 s 79200 20000 80000 20120 6 line[21]
port 124 nsew signal input
rlabel metal3 s 79200 20952 80000 21072 6 line[22]
port 125 nsew signal input
rlabel metal3 s 79200 21904 80000 22024 6 line[23]
port 126 nsew signal input
rlabel metal3 s 79200 22856 80000 22976 6 line[24]
port 127 nsew signal input
rlabel metal3 s 79200 23808 80000 23928 6 line[25]
port 128 nsew signal input
rlabel metal3 s 79200 24760 80000 24880 6 line[26]
port 129 nsew signal input
rlabel metal3 s 79200 25712 80000 25832 6 line[27]
port 130 nsew signal input
rlabel metal3 s 79200 26528 80000 26648 6 line[28]
port 131 nsew signal input
rlabel metal3 s 79200 27480 80000 27600 6 line[29]
port 132 nsew signal input
rlabel metal3 s 79200 2184 80000 2304 6 line[2]
port 133 nsew signal input
rlabel metal3 s 79200 28432 80000 28552 6 line[30]
port 134 nsew signal input
rlabel metal3 s 79200 29384 80000 29504 6 line[31]
port 135 nsew signal input
rlabel metal3 s 79200 30336 80000 30456 6 line[32]
port 136 nsew signal input
rlabel metal3 s 79200 31288 80000 31408 6 line[33]
port 137 nsew signal input
rlabel metal3 s 79200 32240 80000 32360 6 line[34]
port 138 nsew signal input
rlabel metal3 s 79200 33192 80000 33312 6 line[35]
port 139 nsew signal input
rlabel metal3 s 79200 34144 80000 34264 6 line[36]
port 140 nsew signal input
rlabel metal3 s 79200 34960 80000 35080 6 line[37]
port 141 nsew signal input
rlabel metal3 s 79200 35912 80000 36032 6 line[38]
port 142 nsew signal input
rlabel metal3 s 79200 36864 80000 36984 6 line[39]
port 143 nsew signal input
rlabel metal3 s 79200 3136 80000 3256 6 line[3]
port 144 nsew signal input
rlabel metal3 s 79200 37816 80000 37936 6 line[40]
port 145 nsew signal input
rlabel metal3 s 79200 38768 80000 38888 6 line[41]
port 146 nsew signal input
rlabel metal3 s 79200 39720 80000 39840 6 line[42]
port 147 nsew signal input
rlabel metal3 s 79200 40672 80000 40792 6 line[43]
port 148 nsew signal input
rlabel metal3 s 79200 41624 80000 41744 6 line[44]
port 149 nsew signal input
rlabel metal3 s 79200 42576 80000 42696 6 line[45]
port 150 nsew signal input
rlabel metal3 s 79200 43392 80000 43512 6 line[46]
port 151 nsew signal input
rlabel metal3 s 79200 44344 80000 44464 6 line[47]
port 152 nsew signal input
rlabel metal3 s 79200 45296 80000 45416 6 line[48]
port 153 nsew signal input
rlabel metal3 s 79200 46248 80000 46368 6 line[49]
port 154 nsew signal input
rlabel metal3 s 79200 4088 80000 4208 6 line[4]
port 155 nsew signal input
rlabel metal3 s 79200 47200 80000 47320 6 line[50]
port 156 nsew signal input
rlabel metal3 s 79200 48152 80000 48272 6 line[51]
port 157 nsew signal input
rlabel metal3 s 79200 49104 80000 49224 6 line[52]
port 158 nsew signal input
rlabel metal3 s 79200 50056 80000 50176 6 line[53]
port 159 nsew signal input
rlabel metal3 s 79200 51008 80000 51128 6 line[54]
port 160 nsew signal input
rlabel metal3 s 79200 51824 80000 51944 6 line[55]
port 161 nsew signal input
rlabel metal3 s 79200 52776 80000 52896 6 line[56]
port 162 nsew signal input
rlabel metal3 s 79200 53728 80000 53848 6 line[57]
port 163 nsew signal input
rlabel metal3 s 79200 54680 80000 54800 6 line[58]
port 164 nsew signal input
rlabel metal3 s 79200 55632 80000 55752 6 line[59]
port 165 nsew signal input
rlabel metal3 s 79200 5040 80000 5160 6 line[5]
port 166 nsew signal input
rlabel metal3 s 79200 56584 80000 56704 6 line[60]
port 167 nsew signal input
rlabel metal3 s 79200 57536 80000 57656 6 line[61]
port 168 nsew signal input
rlabel metal3 s 79200 58488 80000 58608 6 line[62]
port 169 nsew signal input
rlabel metal3 s 79200 59440 80000 59560 6 line[63]
port 170 nsew signal input
rlabel metal3 s 79200 60392 80000 60512 6 line[64]
port 171 nsew signal input
rlabel metal3 s 79200 61208 80000 61328 6 line[65]
port 172 nsew signal input
rlabel metal3 s 79200 62160 80000 62280 6 line[66]
port 173 nsew signal input
rlabel metal3 s 79200 63112 80000 63232 6 line[67]
port 174 nsew signal input
rlabel metal3 s 79200 64064 80000 64184 6 line[68]
port 175 nsew signal input
rlabel metal3 s 79200 65016 80000 65136 6 line[69]
port 176 nsew signal input
rlabel metal3 s 79200 5992 80000 6112 6 line[6]
port 177 nsew signal input
rlabel metal3 s 79200 65968 80000 66088 6 line[70]
port 178 nsew signal input
rlabel metal3 s 79200 66920 80000 67040 6 line[71]
port 179 nsew signal input
rlabel metal3 s 79200 67872 80000 67992 6 line[72]
port 180 nsew signal input
rlabel metal3 s 79200 68824 80000 68944 6 line[73]
port 181 nsew signal input
rlabel metal3 s 79200 69640 80000 69760 6 line[74]
port 182 nsew signal input
rlabel metal3 s 79200 70592 80000 70712 6 line[75]
port 183 nsew signal input
rlabel metal3 s 79200 71544 80000 71664 6 line[76]
port 184 nsew signal input
rlabel metal3 s 79200 72496 80000 72616 6 line[77]
port 185 nsew signal input
rlabel metal3 s 79200 73448 80000 73568 6 line[78]
port 186 nsew signal input
rlabel metal3 s 79200 74400 80000 74520 6 line[79]
port 187 nsew signal input
rlabel metal3 s 79200 6944 80000 7064 6 line[7]
port 188 nsew signal input
rlabel metal3 s 79200 75352 80000 75472 6 line[80]
port 189 nsew signal input
rlabel metal3 s 79200 76304 80000 76424 6 line[81]
port 190 nsew signal input
rlabel metal3 s 79200 77256 80000 77376 6 line[82]
port 191 nsew signal input
rlabel metal3 s 79200 78072 80000 78192 6 line[83]
port 192 nsew signal input
rlabel metal3 s 79200 79024 80000 79144 6 line[84]
port 193 nsew signal input
rlabel metal3 s 79200 79976 80000 80096 6 line[85]
port 194 nsew signal input
rlabel metal3 s 79200 80928 80000 81048 6 line[86]
port 195 nsew signal input
rlabel metal3 s 79200 81880 80000 82000 6 line[87]
port 196 nsew signal input
rlabel metal3 s 79200 82832 80000 82952 6 line[88]
port 197 nsew signal input
rlabel metal3 s 79200 83784 80000 83904 6 line[89]
port 198 nsew signal input
rlabel metal3 s 79200 7896 80000 8016 6 line[8]
port 199 nsew signal input
rlabel metal3 s 79200 84736 80000 84856 6 line[90]
port 200 nsew signal input
rlabel metal3 s 79200 85688 80000 85808 6 line[91]
port 201 nsew signal input
rlabel metal3 s 79200 86504 80000 86624 6 line[92]
port 202 nsew signal input
rlabel metal3 s 79200 87456 80000 87576 6 line[93]
port 203 nsew signal input
rlabel metal3 s 79200 88408 80000 88528 6 line[94]
port 204 nsew signal input
rlabel metal3 s 79200 89360 80000 89480 6 line[95]
port 205 nsew signal input
rlabel metal3 s 79200 90312 80000 90432 6 line[96]
port 206 nsew signal input
rlabel metal3 s 79200 91264 80000 91384 6 line[97]
port 207 nsew signal input
rlabel metal3 s 79200 92216 80000 92336 6 line[98]
port 208 nsew signal input
rlabel metal3 s 79200 93168 80000 93288 6 line[99]
port 209 nsew signal input
rlabel metal3 s 79200 8848 80000 8968 6 line[9]
port 210 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 rst_n
port 211 nsew signal input
rlabel metal2 s 49974 0 50030 800 6 wr
port 212 nsew signal input
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 213 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 214 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 215 nsew power bidirectional
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 216 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 217 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 80000 120000
string LEFview TRUE
string GDS_FILE /project/openlane/DMC_32x16HC/runs/DMC_32x16HC/results/magic/DMC_32x16HC.gds
string GDS_END 28483382
string GDS_START 234392
<< end >>

