magic
tech sky130A
magscale 1 2
timestamp 1621729262
<< obsli1 >>
rect 1104 2159 79091 117521
<< obsm1 >>
rect 1104 1232 79474 117552
<< metal2 >>
rect 478 119200 534 120000
rect 1490 119200 1546 120000
rect 2594 119200 2650 120000
rect 3698 119200 3754 120000
rect 4802 119200 4858 120000
rect 5814 119200 5870 120000
rect 6918 119200 6974 120000
rect 8022 119200 8078 120000
rect 9126 119200 9182 120000
rect 10138 119200 10194 120000
rect 11242 119200 11298 120000
rect 12346 119200 12402 120000
rect 13450 119200 13506 120000
rect 14462 119200 14518 120000
rect 15566 119200 15622 120000
rect 16670 119200 16726 120000
rect 17774 119200 17830 120000
rect 18786 119200 18842 120000
rect 19890 119200 19946 120000
rect 20994 119200 21050 120000
rect 22098 119200 22154 120000
rect 23110 119200 23166 120000
rect 24214 119200 24270 120000
rect 25318 119200 25374 120000
rect 26422 119200 26478 120000
rect 27434 119200 27490 120000
rect 28538 119200 28594 120000
rect 29642 119200 29698 120000
rect 30746 119200 30802 120000
rect 31758 119200 31814 120000
rect 32862 119200 32918 120000
rect 33966 119200 34022 120000
rect 35070 119200 35126 120000
rect 36082 119200 36138 120000
rect 37186 119200 37242 120000
rect 38290 119200 38346 120000
rect 39394 119200 39450 120000
rect 40498 119200 40554 120000
rect 41510 119200 41566 120000
rect 42614 119200 42670 120000
rect 43718 119200 43774 120000
rect 44822 119200 44878 120000
rect 45834 119200 45890 120000
rect 46938 119200 46994 120000
rect 48042 119200 48098 120000
rect 49146 119200 49202 120000
rect 50158 119200 50214 120000
rect 51262 119200 51318 120000
rect 52366 119200 52422 120000
rect 53470 119200 53526 120000
rect 54482 119200 54538 120000
rect 55586 119200 55642 120000
rect 56690 119200 56746 120000
rect 57794 119200 57850 120000
rect 58806 119200 58862 120000
rect 59910 119200 59966 120000
rect 61014 119200 61070 120000
rect 62118 119200 62174 120000
rect 63130 119200 63186 120000
rect 64234 119200 64290 120000
rect 65338 119200 65394 120000
rect 66442 119200 66498 120000
rect 67454 119200 67510 120000
rect 68558 119200 68614 120000
rect 69662 119200 69718 120000
rect 70766 119200 70822 120000
rect 71778 119200 71834 120000
rect 72882 119200 72938 120000
rect 73986 119200 74042 120000
rect 75090 119200 75146 120000
rect 76102 119200 76158 120000
rect 77206 119200 77262 120000
rect 78310 119200 78366 120000
rect 79414 119200 79470 120000
rect 9954 0 10010 800
rect 29918 0 29974 800
rect 49974 0 50030 800
rect 69938 0 69994 800
<< obsm2 >>
rect 18 119144 422 119513
rect 590 119144 1434 119513
rect 1602 119144 2538 119513
rect 2706 119144 3642 119513
rect 3810 119144 4746 119513
rect 4914 119144 5758 119513
rect 5926 119144 6862 119513
rect 7030 119144 7966 119513
rect 8134 119144 9070 119513
rect 9238 119144 10082 119513
rect 10250 119144 11186 119513
rect 11354 119144 12290 119513
rect 12458 119144 13394 119513
rect 13562 119144 14406 119513
rect 14574 119144 15510 119513
rect 15678 119144 16614 119513
rect 16782 119144 17718 119513
rect 17886 119144 18730 119513
rect 18898 119144 19834 119513
rect 20002 119144 20938 119513
rect 21106 119144 22042 119513
rect 22210 119144 23054 119513
rect 23222 119144 24158 119513
rect 24326 119144 25262 119513
rect 25430 119144 26366 119513
rect 26534 119144 27378 119513
rect 27546 119144 28482 119513
rect 28650 119144 29586 119513
rect 29754 119144 30690 119513
rect 30858 119144 31702 119513
rect 31870 119144 32806 119513
rect 32974 119144 33910 119513
rect 34078 119144 35014 119513
rect 35182 119144 36026 119513
rect 36194 119144 37130 119513
rect 37298 119144 38234 119513
rect 38402 119144 39338 119513
rect 39506 119144 40442 119513
rect 40610 119144 41454 119513
rect 41622 119144 42558 119513
rect 42726 119144 43662 119513
rect 43830 119144 44766 119513
rect 44934 119144 45778 119513
rect 45946 119144 46882 119513
rect 47050 119144 47986 119513
rect 48154 119144 49090 119513
rect 49258 119144 50102 119513
rect 50270 119144 51206 119513
rect 51374 119144 52310 119513
rect 52478 119144 53414 119513
rect 53582 119144 54426 119513
rect 54594 119144 55530 119513
rect 55698 119144 56634 119513
rect 56802 119144 57738 119513
rect 57906 119144 58750 119513
rect 58918 119144 59854 119513
rect 60022 119144 60958 119513
rect 61126 119144 62062 119513
rect 62230 119144 63074 119513
rect 63242 119144 64178 119513
rect 64346 119144 65282 119513
rect 65450 119144 66386 119513
rect 66554 119144 67398 119513
rect 67566 119144 68502 119513
rect 68670 119144 69606 119513
rect 69774 119144 70710 119513
rect 70878 119144 71722 119513
rect 71890 119144 72826 119513
rect 72994 119144 73930 119513
rect 74098 119144 75034 119513
rect 75202 119144 76046 119513
rect 76214 119144 77150 119513
rect 77318 119144 78254 119513
rect 78422 119144 79358 119513
rect 18 856 79468 119144
rect 18 439 9898 856
rect 10066 439 29862 856
rect 30030 439 49918 856
rect 50086 439 69882 856
rect 70050 439 79468 856
<< metal3 >>
rect 79200 119416 80000 119536
rect 79200 118464 80000 118584
rect 79200 117512 80000 117632
rect 79200 116560 80000 116680
rect 79200 115608 80000 115728
rect 79200 114656 80000 114776
rect 79200 113704 80000 113824
rect 79200 112752 80000 112872
rect 79200 111800 80000 111920
rect 79200 110984 80000 111104
rect 79200 110032 80000 110152
rect 79200 109080 80000 109200
rect 79200 108128 80000 108248
rect 79200 107176 80000 107296
rect 79200 106224 80000 106344
rect 79200 105272 80000 105392
rect 79200 104320 80000 104440
rect 79200 103368 80000 103488
rect 79200 102552 80000 102672
rect 79200 101600 80000 101720
rect 79200 100648 80000 100768
rect 79200 99696 80000 99816
rect 79200 98744 80000 98864
rect 79200 97792 80000 97912
rect 79200 96840 80000 96960
rect 79200 95888 80000 96008
rect 79200 94936 80000 95056
rect 79200 94120 80000 94240
rect 79200 93168 80000 93288
rect 79200 92216 80000 92336
rect 79200 91264 80000 91384
rect 79200 90312 80000 90432
rect 79200 89360 80000 89480
rect 79200 88408 80000 88528
rect 79200 87456 80000 87576
rect 79200 86504 80000 86624
rect 79200 85688 80000 85808
rect 79200 84736 80000 84856
rect 79200 83784 80000 83904
rect 79200 82832 80000 82952
rect 79200 81880 80000 82000
rect 79200 80928 80000 81048
rect 79200 79976 80000 80096
rect 79200 79024 80000 79144
rect 79200 78072 80000 78192
rect 79200 77256 80000 77376
rect 79200 76304 80000 76424
rect 79200 75352 80000 75472
rect 79200 74400 80000 74520
rect 79200 73448 80000 73568
rect 79200 72496 80000 72616
rect 79200 71544 80000 71664
rect 79200 70592 80000 70712
rect 79200 69640 80000 69760
rect 79200 68824 80000 68944
rect 79200 67872 80000 67992
rect 79200 66920 80000 67040
rect 79200 65968 80000 66088
rect 79200 65016 80000 65136
rect 79200 64064 80000 64184
rect 79200 63112 80000 63232
rect 79200 62160 80000 62280
rect 79200 61208 80000 61328
rect 79200 60392 80000 60512
rect 79200 59440 80000 59560
rect 79200 58488 80000 58608
rect 79200 57536 80000 57656
rect 79200 56584 80000 56704
rect 79200 55632 80000 55752
rect 79200 54680 80000 54800
rect 79200 53728 80000 53848
rect 79200 52776 80000 52896
rect 79200 51824 80000 51944
rect 79200 51008 80000 51128
rect 79200 50056 80000 50176
rect 79200 49104 80000 49224
rect 79200 48152 80000 48272
rect 79200 47200 80000 47320
rect 79200 46248 80000 46368
rect 79200 45296 80000 45416
rect 79200 44344 80000 44464
rect 79200 43392 80000 43512
rect 79200 42576 80000 42696
rect 79200 41624 80000 41744
rect 79200 40672 80000 40792
rect 79200 39720 80000 39840
rect 79200 38768 80000 38888
rect 79200 37816 80000 37936
rect 79200 36864 80000 36984
rect 79200 35912 80000 36032
rect 79200 34960 80000 35080
rect 79200 34144 80000 34264
rect 79200 33192 80000 33312
rect 79200 32240 80000 32360
rect 79200 31288 80000 31408
rect 79200 30336 80000 30456
rect 79200 29384 80000 29504
rect 79200 28432 80000 28552
rect 79200 27480 80000 27600
rect 79200 26528 80000 26648
rect 79200 25712 80000 25832
rect 79200 24760 80000 24880
rect 79200 23808 80000 23928
rect 79200 22856 80000 22976
rect 79200 21904 80000 22024
rect 79200 20952 80000 21072
rect 79200 20000 80000 20120
rect 79200 19048 80000 19168
rect 79200 18096 80000 18216
rect 79200 17280 80000 17400
rect 79200 16328 80000 16448
rect 79200 15376 80000 15496
rect 79200 14424 80000 14544
rect 79200 13472 80000 13592
rect 79200 12520 80000 12640
rect 79200 11568 80000 11688
rect 79200 10616 80000 10736
rect 79200 9664 80000 9784
rect 79200 8848 80000 8968
rect 79200 7896 80000 8016
rect 79200 6944 80000 7064
rect 79200 5992 80000 6112
rect 79200 5040 80000 5160
rect 79200 4088 80000 4208
rect 79200 3136 80000 3256
rect 79200 2184 80000 2304
rect 79200 1232 80000 1352
rect 79200 416 80000 536
<< obsm3 >>
rect 13 119336 79120 119509
rect 13 118664 79200 119336
rect 13 118384 79120 118664
rect 13 117712 79200 118384
rect 13 117432 79120 117712
rect 13 116760 79200 117432
rect 13 116480 79120 116760
rect 13 115808 79200 116480
rect 13 115528 79120 115808
rect 13 114856 79200 115528
rect 13 114576 79120 114856
rect 13 113904 79200 114576
rect 13 113624 79120 113904
rect 13 112952 79200 113624
rect 13 112672 79120 112952
rect 13 112000 79200 112672
rect 13 111720 79120 112000
rect 13 111184 79200 111720
rect 13 110904 79120 111184
rect 13 110232 79200 110904
rect 13 109952 79120 110232
rect 13 109280 79200 109952
rect 13 109000 79120 109280
rect 13 108328 79200 109000
rect 13 108048 79120 108328
rect 13 107376 79200 108048
rect 13 107096 79120 107376
rect 13 106424 79200 107096
rect 13 106144 79120 106424
rect 13 105472 79200 106144
rect 13 105192 79120 105472
rect 13 104520 79200 105192
rect 13 104240 79120 104520
rect 13 103568 79200 104240
rect 13 103288 79120 103568
rect 13 102752 79200 103288
rect 13 102472 79120 102752
rect 13 101800 79200 102472
rect 13 101520 79120 101800
rect 13 100848 79200 101520
rect 13 100568 79120 100848
rect 13 99896 79200 100568
rect 13 99616 79120 99896
rect 13 98944 79200 99616
rect 13 98664 79120 98944
rect 13 97992 79200 98664
rect 13 97712 79120 97992
rect 13 97040 79200 97712
rect 13 96760 79120 97040
rect 13 96088 79200 96760
rect 13 95808 79120 96088
rect 13 95136 79200 95808
rect 13 94856 79120 95136
rect 13 94320 79200 94856
rect 13 94040 79120 94320
rect 13 93368 79200 94040
rect 13 93088 79120 93368
rect 13 92416 79200 93088
rect 13 92136 79120 92416
rect 13 91464 79200 92136
rect 13 91184 79120 91464
rect 13 90512 79200 91184
rect 13 90232 79120 90512
rect 13 89560 79200 90232
rect 13 89280 79120 89560
rect 13 88608 79200 89280
rect 13 88328 79120 88608
rect 13 87656 79200 88328
rect 13 87376 79120 87656
rect 13 86704 79200 87376
rect 13 86424 79120 86704
rect 13 85888 79200 86424
rect 13 85608 79120 85888
rect 13 84936 79200 85608
rect 13 84656 79120 84936
rect 13 83984 79200 84656
rect 13 83704 79120 83984
rect 13 83032 79200 83704
rect 13 82752 79120 83032
rect 13 82080 79200 82752
rect 13 81800 79120 82080
rect 13 81128 79200 81800
rect 13 80848 79120 81128
rect 13 80176 79200 80848
rect 13 79896 79120 80176
rect 13 79224 79200 79896
rect 13 78944 79120 79224
rect 13 78272 79200 78944
rect 13 77992 79120 78272
rect 13 77456 79200 77992
rect 13 77176 79120 77456
rect 13 76504 79200 77176
rect 13 76224 79120 76504
rect 13 75552 79200 76224
rect 13 75272 79120 75552
rect 13 74600 79200 75272
rect 13 74320 79120 74600
rect 13 73648 79200 74320
rect 13 73368 79120 73648
rect 13 72696 79200 73368
rect 13 72416 79120 72696
rect 13 71744 79200 72416
rect 13 71464 79120 71744
rect 13 70792 79200 71464
rect 13 70512 79120 70792
rect 13 69840 79200 70512
rect 13 69560 79120 69840
rect 13 69024 79200 69560
rect 13 68744 79120 69024
rect 13 68072 79200 68744
rect 13 67792 79120 68072
rect 13 67120 79200 67792
rect 13 66840 79120 67120
rect 13 66168 79200 66840
rect 13 65888 79120 66168
rect 13 65216 79200 65888
rect 13 64936 79120 65216
rect 13 64264 79200 64936
rect 13 63984 79120 64264
rect 13 63312 79200 63984
rect 13 63032 79120 63312
rect 13 62360 79200 63032
rect 13 62080 79120 62360
rect 13 61408 79200 62080
rect 13 61128 79120 61408
rect 13 60592 79200 61128
rect 13 60312 79120 60592
rect 13 59640 79200 60312
rect 13 59360 79120 59640
rect 13 58688 79200 59360
rect 13 58408 79120 58688
rect 13 57736 79200 58408
rect 13 57456 79120 57736
rect 13 56784 79200 57456
rect 13 56504 79120 56784
rect 13 55832 79200 56504
rect 13 55552 79120 55832
rect 13 54880 79200 55552
rect 13 54600 79120 54880
rect 13 53928 79200 54600
rect 13 53648 79120 53928
rect 13 52976 79200 53648
rect 13 52696 79120 52976
rect 13 52024 79200 52696
rect 13 51744 79120 52024
rect 13 51208 79200 51744
rect 13 50928 79120 51208
rect 13 50256 79200 50928
rect 13 49976 79120 50256
rect 13 49304 79200 49976
rect 13 49024 79120 49304
rect 13 48352 79200 49024
rect 13 48072 79120 48352
rect 13 47400 79200 48072
rect 13 47120 79120 47400
rect 13 46448 79200 47120
rect 13 46168 79120 46448
rect 13 45496 79200 46168
rect 13 45216 79120 45496
rect 13 44544 79200 45216
rect 13 44264 79120 44544
rect 13 43592 79200 44264
rect 13 43312 79120 43592
rect 13 42776 79200 43312
rect 13 42496 79120 42776
rect 13 41824 79200 42496
rect 13 41544 79120 41824
rect 13 40872 79200 41544
rect 13 40592 79120 40872
rect 13 39920 79200 40592
rect 13 39640 79120 39920
rect 13 38968 79200 39640
rect 13 38688 79120 38968
rect 13 38016 79200 38688
rect 13 37736 79120 38016
rect 13 37064 79200 37736
rect 13 36784 79120 37064
rect 13 36112 79200 36784
rect 13 35832 79120 36112
rect 13 35160 79200 35832
rect 13 34880 79120 35160
rect 13 34344 79200 34880
rect 13 34064 79120 34344
rect 13 33392 79200 34064
rect 13 33112 79120 33392
rect 13 32440 79200 33112
rect 13 32160 79120 32440
rect 13 31488 79200 32160
rect 13 31208 79120 31488
rect 13 30536 79200 31208
rect 13 30256 79120 30536
rect 13 29584 79200 30256
rect 13 29304 79120 29584
rect 13 28632 79200 29304
rect 13 28352 79120 28632
rect 13 27680 79200 28352
rect 13 27400 79120 27680
rect 13 26728 79200 27400
rect 13 26448 79120 26728
rect 13 25912 79200 26448
rect 13 25632 79120 25912
rect 13 24960 79200 25632
rect 13 24680 79120 24960
rect 13 24008 79200 24680
rect 13 23728 79120 24008
rect 13 23056 79200 23728
rect 13 22776 79120 23056
rect 13 22104 79200 22776
rect 13 21824 79120 22104
rect 13 21152 79200 21824
rect 13 20872 79120 21152
rect 13 20200 79200 20872
rect 13 19920 79120 20200
rect 13 19248 79200 19920
rect 13 18968 79120 19248
rect 13 18296 79200 18968
rect 13 18016 79120 18296
rect 13 17480 79200 18016
rect 13 17200 79120 17480
rect 13 16528 79200 17200
rect 13 16248 79120 16528
rect 13 15576 79200 16248
rect 13 15296 79120 15576
rect 13 14624 79200 15296
rect 13 14344 79120 14624
rect 13 13672 79200 14344
rect 13 13392 79120 13672
rect 13 12720 79200 13392
rect 13 12440 79120 12720
rect 13 11768 79200 12440
rect 13 11488 79120 11768
rect 13 10816 79200 11488
rect 13 10536 79120 10816
rect 13 9864 79200 10536
rect 13 9584 79120 9864
rect 13 9048 79200 9584
rect 13 8768 79120 9048
rect 13 8096 79200 8768
rect 13 7816 79120 8096
rect 13 7144 79200 7816
rect 13 6864 79120 7144
rect 13 6192 79200 6864
rect 13 5912 79120 6192
rect 13 5240 79200 5912
rect 13 4960 79120 5240
rect 13 4288 79200 4960
rect 13 4008 79120 4288
rect 13 3336 79200 4008
rect 13 3056 79120 3336
rect 13 2384 79200 3056
rect 13 2104 79120 2384
rect 13 1432 79200 2104
rect 13 1152 79120 1432
rect 13 616 79200 1152
rect 13 443 79120 616
<< metal4 >>
rect 4208 2128 4528 117552
rect 19568 2128 19888 117552
rect 34928 2128 35248 117552
rect 50288 2128 50608 117552
rect 65648 2128 65968 117552
<< obsm4 >>
rect 14227 5203 19488 114613
rect 19968 5203 34848 114613
rect 35328 5203 50208 114613
rect 50688 5203 65568 114613
rect 66048 5203 74645 114613
<< labels >>
rlabel metal2 s 478 119200 534 120000 6 A[0]
port 1 nsew signal input
rlabel metal2 s 11242 119200 11298 120000 6 A[10]
port 2 nsew signal input
rlabel metal2 s 12346 119200 12402 120000 6 A[11]
port 3 nsew signal input
rlabel metal2 s 13450 119200 13506 120000 6 A[12]
port 4 nsew signal input
rlabel metal2 s 14462 119200 14518 120000 6 A[13]
port 5 nsew signal input
rlabel metal2 s 15566 119200 15622 120000 6 A[14]
port 6 nsew signal input
rlabel metal2 s 16670 119200 16726 120000 6 A[15]
port 7 nsew signal input
rlabel metal2 s 17774 119200 17830 120000 6 A[16]
port 8 nsew signal input
rlabel metal2 s 18786 119200 18842 120000 6 A[17]
port 9 nsew signal input
rlabel metal2 s 19890 119200 19946 120000 6 A[18]
port 10 nsew signal input
rlabel metal2 s 20994 119200 21050 120000 6 A[19]
port 11 nsew signal input
rlabel metal2 s 1490 119200 1546 120000 6 A[1]
port 12 nsew signal input
rlabel metal2 s 22098 119200 22154 120000 6 A[20]
port 13 nsew signal input
rlabel metal2 s 23110 119200 23166 120000 6 A[21]
port 14 nsew signal input
rlabel metal2 s 2594 119200 2650 120000 6 A[2]
port 15 nsew signal input
rlabel metal2 s 3698 119200 3754 120000 6 A[3]
port 16 nsew signal input
rlabel metal2 s 4802 119200 4858 120000 6 A[4]
port 17 nsew signal input
rlabel metal2 s 5814 119200 5870 120000 6 A[5]
port 18 nsew signal input
rlabel metal2 s 6918 119200 6974 120000 6 A[6]
port 19 nsew signal input
rlabel metal2 s 8022 119200 8078 120000 6 A[7]
port 20 nsew signal input
rlabel metal2 s 9126 119200 9182 120000 6 A[8]
port 21 nsew signal input
rlabel metal2 s 10138 119200 10194 120000 6 A[9]
port 22 nsew signal input
rlabel metal2 s 24214 119200 24270 120000 6 A_h[0]
port 23 nsew signal input
rlabel metal2 s 35070 119200 35126 120000 6 A_h[10]
port 24 nsew signal input
rlabel metal2 s 36082 119200 36138 120000 6 A_h[11]
port 25 nsew signal input
rlabel metal2 s 37186 119200 37242 120000 6 A_h[12]
port 26 nsew signal input
rlabel metal2 s 38290 119200 38346 120000 6 A_h[13]
port 27 nsew signal input
rlabel metal2 s 39394 119200 39450 120000 6 A_h[14]
port 28 nsew signal input
rlabel metal2 s 40498 119200 40554 120000 6 A_h[15]
port 29 nsew signal input
rlabel metal2 s 41510 119200 41566 120000 6 A_h[16]
port 30 nsew signal input
rlabel metal2 s 42614 119200 42670 120000 6 A_h[17]
port 31 nsew signal input
rlabel metal2 s 43718 119200 43774 120000 6 A_h[18]
port 32 nsew signal input
rlabel metal2 s 44822 119200 44878 120000 6 A_h[19]
port 33 nsew signal input
rlabel metal2 s 25318 119200 25374 120000 6 A_h[1]
port 34 nsew signal input
rlabel metal2 s 26422 119200 26478 120000 6 A_h[2]
port 35 nsew signal input
rlabel metal2 s 27434 119200 27490 120000 6 A_h[3]
port 36 nsew signal input
rlabel metal2 s 28538 119200 28594 120000 6 A_h[4]
port 37 nsew signal input
rlabel metal2 s 29642 119200 29698 120000 6 A_h[5]
port 38 nsew signal input
rlabel metal2 s 30746 119200 30802 120000 6 A_h[6]
port 39 nsew signal input
rlabel metal2 s 31758 119200 31814 120000 6 A_h[7]
port 40 nsew signal input
rlabel metal2 s 32862 119200 32918 120000 6 A_h[8]
port 41 nsew signal input
rlabel metal2 s 33966 119200 34022 120000 6 A_h[9]
port 42 nsew signal input
rlabel metal2 s 45834 119200 45890 120000 6 Do[0]
port 43 nsew signal output
rlabel metal2 s 56690 119200 56746 120000 6 Do[10]
port 44 nsew signal output
rlabel metal2 s 57794 119200 57850 120000 6 Do[11]
port 45 nsew signal output
rlabel metal2 s 58806 119200 58862 120000 6 Do[12]
port 46 nsew signal output
rlabel metal2 s 59910 119200 59966 120000 6 Do[13]
port 47 nsew signal output
rlabel metal2 s 61014 119200 61070 120000 6 Do[14]
port 48 nsew signal output
rlabel metal2 s 62118 119200 62174 120000 6 Do[15]
port 49 nsew signal output
rlabel metal2 s 63130 119200 63186 120000 6 Do[16]
port 50 nsew signal output
rlabel metal2 s 64234 119200 64290 120000 6 Do[17]
port 51 nsew signal output
rlabel metal2 s 65338 119200 65394 120000 6 Do[18]
port 52 nsew signal output
rlabel metal2 s 66442 119200 66498 120000 6 Do[19]
port 53 nsew signal output
rlabel metal2 s 46938 119200 46994 120000 6 Do[1]
port 54 nsew signal output
rlabel metal2 s 67454 119200 67510 120000 6 Do[20]
port 55 nsew signal output
rlabel metal2 s 68558 119200 68614 120000 6 Do[21]
port 56 nsew signal output
rlabel metal2 s 69662 119200 69718 120000 6 Do[22]
port 57 nsew signal output
rlabel metal2 s 70766 119200 70822 120000 6 Do[23]
port 58 nsew signal output
rlabel metal2 s 71778 119200 71834 120000 6 Do[24]
port 59 nsew signal output
rlabel metal2 s 72882 119200 72938 120000 6 Do[25]
port 60 nsew signal output
rlabel metal2 s 73986 119200 74042 120000 6 Do[26]
port 61 nsew signal output
rlabel metal2 s 75090 119200 75146 120000 6 Do[27]
port 62 nsew signal output
rlabel metal2 s 76102 119200 76158 120000 6 Do[28]
port 63 nsew signal output
rlabel metal2 s 77206 119200 77262 120000 6 Do[29]
port 64 nsew signal output
rlabel metal2 s 48042 119200 48098 120000 6 Do[2]
port 65 nsew signal output
rlabel metal2 s 78310 119200 78366 120000 6 Do[30]
port 66 nsew signal output
rlabel metal2 s 79414 119200 79470 120000 6 Do[31]
port 67 nsew signal output
rlabel metal2 s 49146 119200 49202 120000 6 Do[3]
port 68 nsew signal output
rlabel metal2 s 50158 119200 50214 120000 6 Do[4]
port 69 nsew signal output
rlabel metal2 s 51262 119200 51318 120000 6 Do[5]
port 70 nsew signal output
rlabel metal2 s 52366 119200 52422 120000 6 Do[6]
port 71 nsew signal output
rlabel metal2 s 53470 119200 53526 120000 6 Do[7]
port 72 nsew signal output
rlabel metal2 s 54482 119200 54538 120000 6 Do[8]
port 73 nsew signal output
rlabel metal2 s 55586 119200 55642 120000 6 Do[9]
port 74 nsew signal output
rlabel metal2 s 9954 0 10010 800 6 clk
port 75 nsew signal input
rlabel metal2 s 69938 0 69994 800 6 hit
port 76 nsew signal output
rlabel metal3 s 79200 416 80000 536 6 line[0]
port 77 nsew signal input
rlabel metal3 s 79200 94120 80000 94240 6 line[100]
port 78 nsew signal input
rlabel metal3 s 79200 94936 80000 95056 6 line[101]
port 79 nsew signal input
rlabel metal3 s 79200 95888 80000 96008 6 line[102]
port 80 nsew signal input
rlabel metal3 s 79200 96840 80000 96960 6 line[103]
port 81 nsew signal input
rlabel metal3 s 79200 97792 80000 97912 6 line[104]
port 82 nsew signal input
rlabel metal3 s 79200 98744 80000 98864 6 line[105]
port 83 nsew signal input
rlabel metal3 s 79200 99696 80000 99816 6 line[106]
port 84 nsew signal input
rlabel metal3 s 79200 100648 80000 100768 6 line[107]
port 85 nsew signal input
rlabel metal3 s 79200 101600 80000 101720 6 line[108]
port 86 nsew signal input
rlabel metal3 s 79200 102552 80000 102672 6 line[109]
port 87 nsew signal input
rlabel metal3 s 79200 9664 80000 9784 6 line[10]
port 88 nsew signal input
rlabel metal3 s 79200 103368 80000 103488 6 line[110]
port 89 nsew signal input
rlabel metal3 s 79200 104320 80000 104440 6 line[111]
port 90 nsew signal input
rlabel metal3 s 79200 105272 80000 105392 6 line[112]
port 91 nsew signal input
rlabel metal3 s 79200 106224 80000 106344 6 line[113]
port 92 nsew signal input
rlabel metal3 s 79200 107176 80000 107296 6 line[114]
port 93 nsew signal input
rlabel metal3 s 79200 108128 80000 108248 6 line[115]
port 94 nsew signal input
rlabel metal3 s 79200 109080 80000 109200 6 line[116]
port 95 nsew signal input
rlabel metal3 s 79200 110032 80000 110152 6 line[117]
port 96 nsew signal input
rlabel metal3 s 79200 110984 80000 111104 6 line[118]
port 97 nsew signal input
rlabel metal3 s 79200 111800 80000 111920 6 line[119]
port 98 nsew signal input
rlabel metal3 s 79200 10616 80000 10736 6 line[11]
port 99 nsew signal input
rlabel metal3 s 79200 112752 80000 112872 6 line[120]
port 100 nsew signal input
rlabel metal3 s 79200 113704 80000 113824 6 line[121]
port 101 nsew signal input
rlabel metal3 s 79200 114656 80000 114776 6 line[122]
port 102 nsew signal input
rlabel metal3 s 79200 115608 80000 115728 6 line[123]
port 103 nsew signal input
rlabel metal3 s 79200 116560 80000 116680 6 line[124]
port 104 nsew signal input
rlabel metal3 s 79200 117512 80000 117632 6 line[125]
port 105 nsew signal input
rlabel metal3 s 79200 118464 80000 118584 6 line[126]
port 106 nsew signal input
rlabel metal3 s 79200 119416 80000 119536 6 line[127]
port 107 nsew signal input
rlabel metal3 s 79200 11568 80000 11688 6 line[12]
port 108 nsew signal input
rlabel metal3 s 79200 12520 80000 12640 6 line[13]
port 109 nsew signal input
rlabel metal3 s 79200 13472 80000 13592 6 line[14]
port 110 nsew signal input
rlabel metal3 s 79200 14424 80000 14544 6 line[15]
port 111 nsew signal input
rlabel metal3 s 79200 15376 80000 15496 6 line[16]
port 112 nsew signal input
rlabel metal3 s 79200 16328 80000 16448 6 line[17]
port 113 nsew signal input
rlabel metal3 s 79200 17280 80000 17400 6 line[18]
port 114 nsew signal input
rlabel metal3 s 79200 18096 80000 18216 6 line[19]
port 115 nsew signal input
rlabel metal3 s 79200 1232 80000 1352 6 line[1]
port 116 nsew signal input
rlabel metal3 s 79200 19048 80000 19168 6 line[20]
port 117 nsew signal input
rlabel metal3 s 79200 20000 80000 20120 6 line[21]
port 118 nsew signal input
rlabel metal3 s 79200 20952 80000 21072 6 line[22]
port 119 nsew signal input
rlabel metal3 s 79200 21904 80000 22024 6 line[23]
port 120 nsew signal input
rlabel metal3 s 79200 22856 80000 22976 6 line[24]
port 121 nsew signal input
rlabel metal3 s 79200 23808 80000 23928 6 line[25]
port 122 nsew signal input
rlabel metal3 s 79200 24760 80000 24880 6 line[26]
port 123 nsew signal input
rlabel metal3 s 79200 25712 80000 25832 6 line[27]
port 124 nsew signal input
rlabel metal3 s 79200 26528 80000 26648 6 line[28]
port 125 nsew signal input
rlabel metal3 s 79200 27480 80000 27600 6 line[29]
port 126 nsew signal input
rlabel metal3 s 79200 2184 80000 2304 6 line[2]
port 127 nsew signal input
rlabel metal3 s 79200 28432 80000 28552 6 line[30]
port 128 nsew signal input
rlabel metal3 s 79200 29384 80000 29504 6 line[31]
port 129 nsew signal input
rlabel metal3 s 79200 30336 80000 30456 6 line[32]
port 130 nsew signal input
rlabel metal3 s 79200 31288 80000 31408 6 line[33]
port 131 nsew signal input
rlabel metal3 s 79200 32240 80000 32360 6 line[34]
port 132 nsew signal input
rlabel metal3 s 79200 33192 80000 33312 6 line[35]
port 133 nsew signal input
rlabel metal3 s 79200 34144 80000 34264 6 line[36]
port 134 nsew signal input
rlabel metal3 s 79200 34960 80000 35080 6 line[37]
port 135 nsew signal input
rlabel metal3 s 79200 35912 80000 36032 6 line[38]
port 136 nsew signal input
rlabel metal3 s 79200 36864 80000 36984 6 line[39]
port 137 nsew signal input
rlabel metal3 s 79200 3136 80000 3256 6 line[3]
port 138 nsew signal input
rlabel metal3 s 79200 37816 80000 37936 6 line[40]
port 139 nsew signal input
rlabel metal3 s 79200 38768 80000 38888 6 line[41]
port 140 nsew signal input
rlabel metal3 s 79200 39720 80000 39840 6 line[42]
port 141 nsew signal input
rlabel metal3 s 79200 40672 80000 40792 6 line[43]
port 142 nsew signal input
rlabel metal3 s 79200 41624 80000 41744 6 line[44]
port 143 nsew signal input
rlabel metal3 s 79200 42576 80000 42696 6 line[45]
port 144 nsew signal input
rlabel metal3 s 79200 43392 80000 43512 6 line[46]
port 145 nsew signal input
rlabel metal3 s 79200 44344 80000 44464 6 line[47]
port 146 nsew signal input
rlabel metal3 s 79200 45296 80000 45416 6 line[48]
port 147 nsew signal input
rlabel metal3 s 79200 46248 80000 46368 6 line[49]
port 148 nsew signal input
rlabel metal3 s 79200 4088 80000 4208 6 line[4]
port 149 nsew signal input
rlabel metal3 s 79200 47200 80000 47320 6 line[50]
port 150 nsew signal input
rlabel metal3 s 79200 48152 80000 48272 6 line[51]
port 151 nsew signal input
rlabel metal3 s 79200 49104 80000 49224 6 line[52]
port 152 nsew signal input
rlabel metal3 s 79200 50056 80000 50176 6 line[53]
port 153 nsew signal input
rlabel metal3 s 79200 51008 80000 51128 6 line[54]
port 154 nsew signal input
rlabel metal3 s 79200 51824 80000 51944 6 line[55]
port 155 nsew signal input
rlabel metal3 s 79200 52776 80000 52896 6 line[56]
port 156 nsew signal input
rlabel metal3 s 79200 53728 80000 53848 6 line[57]
port 157 nsew signal input
rlabel metal3 s 79200 54680 80000 54800 6 line[58]
port 158 nsew signal input
rlabel metal3 s 79200 55632 80000 55752 6 line[59]
port 159 nsew signal input
rlabel metal3 s 79200 5040 80000 5160 6 line[5]
port 160 nsew signal input
rlabel metal3 s 79200 56584 80000 56704 6 line[60]
port 161 nsew signal input
rlabel metal3 s 79200 57536 80000 57656 6 line[61]
port 162 nsew signal input
rlabel metal3 s 79200 58488 80000 58608 6 line[62]
port 163 nsew signal input
rlabel metal3 s 79200 59440 80000 59560 6 line[63]
port 164 nsew signal input
rlabel metal3 s 79200 60392 80000 60512 6 line[64]
port 165 nsew signal input
rlabel metal3 s 79200 61208 80000 61328 6 line[65]
port 166 nsew signal input
rlabel metal3 s 79200 62160 80000 62280 6 line[66]
port 167 nsew signal input
rlabel metal3 s 79200 63112 80000 63232 6 line[67]
port 168 nsew signal input
rlabel metal3 s 79200 64064 80000 64184 6 line[68]
port 169 nsew signal input
rlabel metal3 s 79200 65016 80000 65136 6 line[69]
port 170 nsew signal input
rlabel metal3 s 79200 5992 80000 6112 6 line[6]
port 171 nsew signal input
rlabel metal3 s 79200 65968 80000 66088 6 line[70]
port 172 nsew signal input
rlabel metal3 s 79200 66920 80000 67040 6 line[71]
port 173 nsew signal input
rlabel metal3 s 79200 67872 80000 67992 6 line[72]
port 174 nsew signal input
rlabel metal3 s 79200 68824 80000 68944 6 line[73]
port 175 nsew signal input
rlabel metal3 s 79200 69640 80000 69760 6 line[74]
port 176 nsew signal input
rlabel metal3 s 79200 70592 80000 70712 6 line[75]
port 177 nsew signal input
rlabel metal3 s 79200 71544 80000 71664 6 line[76]
port 178 nsew signal input
rlabel metal3 s 79200 72496 80000 72616 6 line[77]
port 179 nsew signal input
rlabel metal3 s 79200 73448 80000 73568 6 line[78]
port 180 nsew signal input
rlabel metal3 s 79200 74400 80000 74520 6 line[79]
port 181 nsew signal input
rlabel metal3 s 79200 6944 80000 7064 6 line[7]
port 182 nsew signal input
rlabel metal3 s 79200 75352 80000 75472 6 line[80]
port 183 nsew signal input
rlabel metal3 s 79200 76304 80000 76424 6 line[81]
port 184 nsew signal input
rlabel metal3 s 79200 77256 80000 77376 6 line[82]
port 185 nsew signal input
rlabel metal3 s 79200 78072 80000 78192 6 line[83]
port 186 nsew signal input
rlabel metal3 s 79200 79024 80000 79144 6 line[84]
port 187 nsew signal input
rlabel metal3 s 79200 79976 80000 80096 6 line[85]
port 188 nsew signal input
rlabel metal3 s 79200 80928 80000 81048 6 line[86]
port 189 nsew signal input
rlabel metal3 s 79200 81880 80000 82000 6 line[87]
port 190 nsew signal input
rlabel metal3 s 79200 82832 80000 82952 6 line[88]
port 191 nsew signal input
rlabel metal3 s 79200 83784 80000 83904 6 line[89]
port 192 nsew signal input
rlabel metal3 s 79200 7896 80000 8016 6 line[8]
port 193 nsew signal input
rlabel metal3 s 79200 84736 80000 84856 6 line[90]
port 194 nsew signal input
rlabel metal3 s 79200 85688 80000 85808 6 line[91]
port 195 nsew signal input
rlabel metal3 s 79200 86504 80000 86624 6 line[92]
port 196 nsew signal input
rlabel metal3 s 79200 87456 80000 87576 6 line[93]
port 197 nsew signal input
rlabel metal3 s 79200 88408 80000 88528 6 line[94]
port 198 nsew signal input
rlabel metal3 s 79200 89360 80000 89480 6 line[95]
port 199 nsew signal input
rlabel metal3 s 79200 90312 80000 90432 6 line[96]
port 200 nsew signal input
rlabel metal3 s 79200 91264 80000 91384 6 line[97]
port 201 nsew signal input
rlabel metal3 s 79200 92216 80000 92336 6 line[98]
port 202 nsew signal input
rlabel metal3 s 79200 93168 80000 93288 6 line[99]
port 203 nsew signal input
rlabel metal3 s 79200 8848 80000 8968 6 line[9]
port 204 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 rst_n
port 205 nsew signal input
rlabel metal2 s 49974 0 50030 800 6 wr
port 206 nsew signal input
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 207 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 208 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 209 nsew power bidirectional
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 210 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 211 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 80000 120000
string LEFview TRUE
string GDS_FILE /project/openlane/DMC_32x16HC/runs/DMC_32x16HC/results/magic/DMC_32x16HC.gds
string GDS_END 28100238
string GDS_START 234392
<< end >>

