VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO DFFRAM_1Kx32
  CLASS BLOCK ;
  FOREIGN DFFRAM_1Kx32 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1100.000 BY 1400.000 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.290 1396.000 446.570 1400.000 ;
    END
  END A[0]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.090 1396.000 460.370 1400.000 ;
    END
  END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.890 1396.000 474.170 1400.000 ;
    END
  END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.690 1396.000 487.970 1400.000 ;
    END
  END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.030 1396.000 501.310 1400.000 ;
    END
  END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.830 1396.000 515.110 1400.000 ;
    END
  END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.630 1396.000 528.910 1400.000 ;
    END
  END A[6]
  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.430 1396.000 542.710 1400.000 ;
    END
  END A[7]
  PIN A[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.230 1396.000 556.510 1400.000 ;
    END
  END A[8]
  PIN A[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.030 1396.000 570.310 1400.000 ;
    END
  END A[9]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 583.830 1396.000 584.110 1400.000 ;
    END
  END CLK
  PIN Di[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.170 1396.000 666.450 1400.000 ;
    END
  END Di[0]
  PIN Di[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 803.710 1396.000 803.990 1400.000 ;
    END
  END Di[10]
  PIN Di[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.510 1396.000 817.790 1400.000 ;
    END
  END Di[11]
  PIN Di[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 831.310 1396.000 831.590 1400.000 ;
    END
  END Di[12]
  PIN Di[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 845.110 1396.000 845.390 1400.000 ;
    END
  END Di[13]
  PIN Di[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 858.910 1396.000 859.190 1400.000 ;
    END
  END Di[14]
  PIN Di[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 872.250 1396.000 872.530 1400.000 ;
    END
  END Di[15]
  PIN Di[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 886.050 1396.000 886.330 1400.000 ;
    END
  END Di[16]
  PIN Di[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 899.850 1396.000 900.130 1400.000 ;
    END
  END Di[17]
  PIN Di[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 913.650 1396.000 913.930 1400.000 ;
    END
  END Di[18]
  PIN Di[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.450 1396.000 927.730 1400.000 ;
    END
  END Di[19]
  PIN Di[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.970 1396.000 680.250 1400.000 ;
    END
  END Di[1]
  PIN Di[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 941.250 1396.000 941.530 1400.000 ;
    END
  END Di[20]
  PIN Di[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 955.050 1396.000 955.330 1400.000 ;
    END
  END Di[21]
  PIN Di[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 968.850 1396.000 969.130 1400.000 ;
    END
  END Di[22]
  PIN Di[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 982.650 1396.000 982.930 1400.000 ;
    END
  END Di[23]
  PIN Di[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.990 1396.000 996.270 1400.000 ;
    END
  END Di[24]
  PIN Di[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1009.790 1396.000 1010.070 1400.000 ;
    END
  END Di[25]
  PIN Di[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1023.590 1396.000 1023.870 1400.000 ;
    END
  END Di[26]
  PIN Di[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1037.390 1396.000 1037.670 1400.000 ;
    END
  END Di[27]
  PIN Di[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1051.190 1396.000 1051.470 1400.000 ;
    END
  END Di[28]
  PIN Di[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1064.990 1396.000 1065.270 1400.000 ;
    END
  END Di[29]
  PIN Di[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 693.770 1396.000 694.050 1400.000 ;
    END
  END Di[2]
  PIN Di[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1078.790 1396.000 1079.070 1400.000 ;
    END
  END Di[30]
  PIN Di[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1092.590 1396.000 1092.870 1400.000 ;
    END
  END Di[31]
  PIN Di[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.570 1396.000 707.850 1400.000 ;
    END
  END Di[3]
  PIN Di[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.370 1396.000 721.650 1400.000 ;
    END
  END Di[4]
  PIN Di[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.170 1396.000 735.450 1400.000 ;
    END
  END Di[5]
  PIN Di[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.510 1396.000 748.790 1400.000 ;
    END
  END Di[6]
  PIN Di[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 762.310 1396.000 762.590 1400.000 ;
    END
  END Di[7]
  PIN Di[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.110 1396.000 776.390 1400.000 ;
    END
  END Di[8]
  PIN Di[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.910 1396.000 790.190 1400.000 ;
    END
  END Di[9]
  PIN Do[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 1396.000 6.810 1400.000 ;
    END
  END Do[0]
  PIN Do[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 1396.000 143.890 1400.000 ;
    END
  END Do[10]
  PIN Do[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.410 1396.000 157.690 1400.000 ;
    END
  END Do[11]
  PIN Do[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.210 1396.000 171.490 1400.000 ;
    END
  END Do[12]
  PIN Do[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 1396.000 185.290 1400.000 ;
    END
  END Do[13]
  PIN Do[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.810 1396.000 199.090 1400.000 ;
    END
  END Do[14]
  PIN Do[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 1396.000 212.890 1400.000 ;
    END
  END Do[15]
  PIN Do[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 1396.000 226.690 1400.000 ;
    END
  END Do[16]
  PIN Do[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.210 1396.000 240.490 1400.000 ;
    END
  END Do[17]
  PIN Do[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.550 1396.000 253.830 1400.000 ;
    END
  END Do[18]
  PIN Do[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 1396.000 267.630 1400.000 ;
    END
  END Do[19]
  PIN Do[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 1396.000 20.150 1400.000 ;
    END
  END Do[1]
  PIN Do[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.150 1396.000 281.430 1400.000 ;
    END
  END Do[20]
  PIN Do[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.950 1396.000 295.230 1400.000 ;
    END
  END Do[21]
  PIN Do[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.750 1396.000 309.030 1400.000 ;
    END
  END Do[22]
  PIN Do[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.550 1396.000 322.830 1400.000 ;
    END
  END Do[23]
  PIN Do[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.350 1396.000 336.630 1400.000 ;
    END
  END Do[24]
  PIN Do[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.150 1396.000 350.430 1400.000 ;
    END
  END Do[25]
  PIN Do[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 1396.000 364.230 1400.000 ;
    END
  END Do[26]
  PIN Do[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.290 1396.000 377.570 1400.000 ;
    END
  END Do[27]
  PIN Do[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.090 1396.000 391.370 1400.000 ;
    END
  END Do[28]
  PIN Do[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.890 1396.000 405.170 1400.000 ;
    END
  END Do[29]
  PIN Do[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 1396.000 33.950 1400.000 ;
    END
  END Do[2]
  PIN Do[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 1396.000 418.970 1400.000 ;
    END
  END Do[30]
  PIN Do[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.490 1396.000 432.770 1400.000 ;
    END
  END Do[31]
  PIN Do[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 1396.000 47.750 1400.000 ;
    END
  END Do[3]
  PIN Do[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 1396.000 61.550 1400.000 ;
    END
  END Do[4]
  PIN Do[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 1396.000 75.350 1400.000 ;
    END
  END Do[5]
  PIN Do[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 1396.000 89.150 1400.000 ;
    END
  END Do[6]
  PIN Do[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.670 1396.000 102.950 1400.000 ;
    END
  END Do[7]
  PIN Do[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.470 1396.000 116.750 1400.000 ;
    END
  END Do[8]
  PIN Do[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 1396.000 130.090 1400.000 ;
    END
  END Do[9]
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.370 1396.000 652.650 1400.000 ;
    END
  END EN
  PIN WE[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.630 1396.000 597.910 1400.000 ;
    END
  END WE[0]
  PIN WE[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.430 1396.000 611.710 1400.000 ;
    END
  END WE[1]
  PIN WE[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.770 1396.000 625.050 1400.000 ;
    END
  END WE[2]
  PIN WE[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 638.570 1396.000 638.850 1400.000 ;
    END
  END WE[3]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1387.440 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1387.440 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1387.440 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1387.440 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1387.440 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1387.440 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1387.440 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1387.440 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1387.440 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1387.440 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1387.440 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1387.440 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1387.440 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1387.440 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 1385.785 1094.530 1387.390 ;
        RECT 5.330 1380.345 1094.530 1383.175 ;
        RECT 5.330 1374.905 1094.530 1377.735 ;
        RECT 5.330 1369.515 1094.530 1372.295 ;
        RECT 5.330 1369.465 430.240 1369.515 ;
        RECT 5.330 1366.805 111.855 1366.855 ;
        RECT 5.330 1364.075 1094.530 1366.805 ;
        RECT 5.330 1364.025 67.760 1364.075 ;
        RECT 5.330 1361.365 83.795 1361.415 ;
        RECT 5.330 1358.635 1094.530 1361.365 ;
        RECT 5.330 1358.585 72.820 1358.635 ;
        RECT 5.330 1355.925 127.035 1355.975 ;
        RECT 5.330 1353.195 1094.530 1355.925 ;
        RECT 5.330 1353.145 202.935 1353.195 ;
        RECT 5.330 1350.485 615.555 1350.535 ;
        RECT 5.330 1347.755 1094.530 1350.485 ;
        RECT 5.330 1347.705 111.855 1347.755 ;
        RECT 5.330 1345.045 304.200 1345.095 ;
        RECT 5.330 1342.315 1094.530 1345.045 ;
        RECT 5.330 1342.265 260.435 1342.315 ;
        RECT 5.330 1339.605 39.240 1339.655 ;
        RECT 5.330 1336.875 1094.530 1339.605 ;
        RECT 5.330 1336.825 70.980 1336.875 ;
        RECT 5.330 1334.165 33.260 1334.215 ;
        RECT 5.330 1331.435 1094.530 1334.165 ;
        RECT 5.330 1331.385 42.855 1331.435 ;
        RECT 5.330 1328.725 31.880 1328.775 ;
        RECT 5.330 1325.995 1094.530 1328.725 ;
        RECT 5.330 1325.945 78.735 1325.995 ;
        RECT 5.330 1323.285 29.055 1323.335 ;
        RECT 5.330 1320.555 1094.530 1323.285 ;
        RECT 5.330 1320.505 127.955 1320.555 ;
        RECT 5.330 1317.845 30.960 1317.895 ;
        RECT 5.330 1315.115 1094.530 1317.845 ;
        RECT 5.330 1315.065 260.960 1315.115 ;
        RECT 5.330 1312.405 151.875 1312.455 ;
        RECT 5.330 1309.675 1094.530 1312.405 ;
        RECT 5.330 1309.625 183.615 1309.675 ;
        RECT 5.330 1306.965 29.515 1307.015 ;
        RECT 5.330 1304.235 1094.530 1306.965 ;
        RECT 5.330 1304.185 71.375 1304.235 ;
        RECT 5.330 1301.525 75.515 1301.575 ;
        RECT 5.330 1298.795 1094.530 1301.525 ;
        RECT 5.330 1298.745 126.575 1298.795 ;
        RECT 5.330 1296.085 549.380 1296.135 ;
        RECT 5.330 1293.355 1094.530 1296.085 ;
        RECT 5.330 1293.305 283.435 1293.355 ;
        RECT 5.330 1290.645 266.875 1290.695 ;
        RECT 5.330 1287.915 1094.530 1290.645 ;
        RECT 5.330 1287.865 200.635 1287.915 ;
        RECT 5.330 1285.205 32.800 1285.255 ;
        RECT 5.330 1282.475 1094.530 1285.205 ;
        RECT 5.330 1282.425 36.020 1282.475 ;
        RECT 5.330 1279.765 396.135 1279.815 ;
        RECT 5.330 1277.035 1094.530 1279.765 ;
        RECT 5.330 1276.985 52.055 1277.035 ;
        RECT 5.330 1274.325 31.815 1274.375 ;
        RECT 5.330 1271.595 1094.530 1274.325 ;
        RECT 5.330 1271.545 182.695 1271.595 ;
        RECT 5.330 1268.885 34.180 1268.935 ;
        RECT 5.330 1266.155 1094.530 1268.885 ;
        RECT 5.330 1266.105 33.655 1266.155 ;
        RECT 5.330 1263.445 157.855 1263.495 ;
        RECT 5.330 1260.715 1094.530 1263.445 ;
        RECT 5.330 1260.665 36.020 1260.715 ;
        RECT 5.330 1258.005 32.275 1258.055 ;
        RECT 5.330 1255.275 1094.530 1258.005 ;
        RECT 5.330 1255.225 200.175 1255.275 ;
        RECT 5.330 1252.565 31.420 1252.615 ;
        RECT 5.330 1249.835 1094.530 1252.565 ;
        RECT 5.330 1249.785 59.415 1249.835 ;
        RECT 5.330 1247.125 50.675 1247.175 ;
        RECT 5.330 1244.395 1094.530 1247.125 ;
        RECT 5.330 1244.345 50.280 1244.395 ;
        RECT 5.330 1241.685 28.595 1241.735 ;
        RECT 5.330 1238.955 1094.530 1241.685 ;
        RECT 5.330 1238.905 26.295 1238.955 ;
        RECT 5.330 1236.245 91.680 1236.295 ;
        RECT 5.330 1233.515 1094.530 1236.245 ;
        RECT 5.330 1233.465 1025.020 1233.515 ;
        RECT 5.330 1230.805 68.680 1230.855 ;
        RECT 5.330 1228.075 1094.530 1230.805 ;
        RECT 5.330 1228.025 157.395 1228.075 ;
        RECT 5.330 1225.365 81.035 1225.415 ;
        RECT 5.330 1222.635 1094.530 1225.365 ;
        RECT 5.330 1222.585 71.440 1222.635 ;
        RECT 5.330 1219.925 126.115 1219.975 ;
        RECT 5.330 1217.195 1094.530 1219.925 ;
        RECT 5.330 1217.145 69.600 1217.195 ;
        RECT 5.330 1214.485 75.580 1214.535 ;
        RECT 5.330 1211.755 1094.530 1214.485 ;
        RECT 5.330 1211.705 69.075 1211.755 ;
        RECT 5.330 1209.045 317.475 1209.095 ;
        RECT 5.330 1206.315 1094.530 1209.045 ;
        RECT 5.330 1206.265 70.060 1206.315 ;
        RECT 5.330 1203.605 101.800 1203.655 ;
        RECT 5.330 1200.875 1094.530 1203.605 ;
        RECT 5.330 1200.825 71.900 1200.875 ;
        RECT 5.330 1198.165 317.475 1198.215 ;
        RECT 5.330 1195.435 1094.530 1198.165 ;
        RECT 5.330 1195.385 149.115 1195.435 ;
        RECT 5.330 1192.725 548.460 1192.775 ;
        RECT 5.330 1189.995 1094.530 1192.725 ;
        RECT 5.330 1189.945 882.420 1189.995 ;
        RECT 5.330 1184.555 1094.530 1187.335 ;
        RECT 5.330 1184.505 848.840 1184.555 ;
        RECT 5.330 1181.845 283.435 1181.895 ;
        RECT 5.330 1179.115 1094.530 1181.845 ;
        RECT 5.330 1179.065 852.980 1179.115 ;
        RECT 5.330 1176.405 259.120 1176.455 ;
        RECT 5.330 1173.675 1094.530 1176.405 ;
        RECT 5.330 1173.625 299.995 1173.675 ;
        RECT 5.330 1170.965 259.580 1171.015 ;
        RECT 5.330 1168.235 1094.530 1170.965 ;
        RECT 5.330 1168.185 432.540 1168.235 ;
        RECT 5.330 1165.525 28.200 1165.575 ;
        RECT 5.330 1162.795 1094.530 1165.525 ;
        RECT 5.330 1162.745 27.280 1162.795 ;
        RECT 5.330 1160.085 42.460 1160.135 ;
        RECT 5.330 1157.355 1094.530 1160.085 ;
        RECT 5.330 1157.305 59.875 1157.355 ;
        RECT 5.330 1154.645 23.140 1154.695 ;
        RECT 5.330 1151.915 1094.530 1154.645 ;
        RECT 5.330 1151.865 25.440 1151.915 ;
        RECT 5.330 1149.205 56.195 1149.255 ;
        RECT 5.330 1146.475 1094.530 1149.205 ;
        RECT 5.330 1146.425 157.395 1146.475 ;
        RECT 5.330 1143.765 259.120 1143.815 ;
        RECT 5.330 1141.035 1094.530 1143.765 ;
        RECT 5.330 1140.985 259.975 1141.035 ;
        RECT 5.330 1138.325 501.475 1138.375 ;
        RECT 5.330 1135.595 1094.530 1138.325 ;
        RECT 5.330 1135.545 591.635 1135.595 ;
        RECT 5.330 1132.885 770.575 1132.935 ;
        RECT 5.330 1130.155 1094.530 1132.885 ;
        RECT 5.330 1130.105 17.555 1130.155 ;
        RECT 5.330 1127.445 166.135 1127.495 ;
        RECT 5.330 1124.715 1094.530 1127.445 ;
        RECT 5.330 1124.665 299.075 1124.715 ;
        RECT 5.330 1122.005 931.115 1122.055 ;
        RECT 5.330 1119.275 1094.530 1122.005 ;
        RECT 5.330 1119.225 257.740 1119.275 ;
        RECT 5.330 1116.565 241.180 1116.615 ;
        RECT 5.330 1113.835 1094.530 1116.565 ;
        RECT 5.330 1113.785 335.875 1113.835 ;
        RECT 5.330 1111.125 885.575 1111.175 ;
        RECT 5.330 1108.395 1094.530 1111.125 ;
        RECT 5.330 1108.345 94.375 1108.395 ;
        RECT 5.330 1105.685 31.420 1105.735 ;
        RECT 5.330 1102.955 1094.530 1105.685 ;
        RECT 5.330 1102.905 59.415 1102.955 ;
        RECT 5.330 1100.245 32.340 1100.295 ;
        RECT 5.330 1097.515 1094.530 1100.245 ;
        RECT 5.330 1097.465 72.820 1097.515 ;
        RECT 5.330 1094.805 28.135 1094.855 ;
        RECT 5.330 1092.075 1094.530 1094.805 ;
        RECT 5.330 1092.025 156.015 1092.075 ;
        RECT 5.330 1089.365 29.055 1089.415 ;
        RECT 5.330 1086.635 1094.530 1089.365 ;
        RECT 5.330 1086.585 29.120 1086.635 ;
        RECT 5.330 1083.925 153.255 1083.975 ;
        RECT 5.330 1081.195 1094.530 1083.925 ;
        RECT 5.330 1081.145 250.775 1081.195 ;
        RECT 5.330 1078.485 76.500 1078.535 ;
        RECT 5.330 1075.755 1094.530 1078.485 ;
        RECT 5.330 1075.705 183.615 1075.755 ;
        RECT 5.330 1073.045 24.520 1073.095 ;
        RECT 5.330 1070.315 1094.530 1073.045 ;
        RECT 5.330 1070.265 111.855 1070.315 ;
        RECT 5.330 1067.605 244.795 1067.655 ;
        RECT 5.330 1064.875 1094.530 1067.605 ;
        RECT 5.330 1064.825 452.715 1064.875 ;
        RECT 5.330 1062.165 151.415 1062.215 ;
        RECT 5.330 1059.435 1094.530 1062.165 ;
        RECT 5.330 1059.385 145.435 1059.435 ;
        RECT 5.330 1056.725 30.500 1056.775 ;
        RECT 5.330 1053.995 1094.530 1056.725 ;
        RECT 5.330 1053.945 70.980 1053.995 ;
        RECT 5.330 1051.285 39.635 1051.335 ;
        RECT 5.330 1048.555 1094.530 1051.285 ;
        RECT 5.330 1048.505 43.380 1048.555 ;
        RECT 5.330 1045.845 260.040 1045.895 ;
        RECT 5.330 1043.115 1094.530 1045.845 ;
        RECT 5.330 1043.065 172.575 1043.115 ;
        RECT 5.330 1040.405 186.375 1040.455 ;
        RECT 5.330 1037.675 1094.530 1040.405 ;
        RECT 5.330 1037.625 323.455 1037.675 ;
        RECT 5.330 1034.965 593.080 1035.015 ;
        RECT 5.330 1032.235 1094.530 1034.965 ;
        RECT 5.330 1032.185 25.440 1032.235 ;
        RECT 5.330 1029.525 30.500 1029.575 ;
        RECT 5.330 1026.795 1094.530 1029.525 ;
        RECT 5.330 1026.745 28.660 1026.795 ;
        RECT 5.330 1024.085 31.880 1024.135 ;
        RECT 5.330 1021.355 1094.530 1024.085 ;
        RECT 5.330 1021.305 34.575 1021.355 ;
        RECT 5.330 1018.645 46.535 1018.695 ;
        RECT 5.330 1015.915 1094.530 1018.645 ;
        RECT 5.330 1015.865 70.455 1015.915 ;
        RECT 5.330 1013.205 185.915 1013.255 ;
        RECT 5.330 1010.475 1094.530 1013.205 ;
        RECT 5.330 1010.425 452.715 1010.475 ;
        RECT 5.330 1007.765 448.115 1007.815 ;
        RECT 5.330 1005.035 1094.530 1007.765 ;
        RECT 5.330 1004.985 21.300 1005.035 ;
        RECT 5.330 1002.325 159.695 1002.375 ;
        RECT 5.330 999.595 1094.530 1002.325 ;
        RECT 5.330 999.545 177.635 999.595 ;
        RECT 5.330 996.885 84.715 996.935 ;
        RECT 5.330 994.155 1094.530 996.885 ;
        RECT 5.330 994.105 29.120 994.155 ;
        RECT 5.330 991.445 100.815 991.495 ;
        RECT 5.330 988.715 1094.530 991.445 ;
        RECT 5.330 988.665 25.440 988.715 ;
        RECT 5.330 986.005 87.475 986.055 ;
        RECT 5.330 983.275 1094.530 986.005 ;
        RECT 5.330 983.225 72.755 983.275 ;
        RECT 5.330 980.565 118.360 980.615 ;
        RECT 5.330 977.835 1094.530 980.565 ;
        RECT 5.330 977.785 129.335 977.835 ;
        RECT 5.330 975.125 24.980 975.175 ;
        RECT 5.330 972.395 1094.530 975.125 ;
        RECT 5.330 972.345 45.155 972.395 ;
        RECT 5.330 969.685 28.135 969.735 ;
        RECT 5.330 966.955 1094.530 969.685 ;
        RECT 5.330 966.905 60.795 966.955 ;
        RECT 5.330 964.245 158.380 964.295 ;
        RECT 5.330 961.515 1094.530 964.245 ;
        RECT 5.330 961.465 160.220 961.515 ;
        RECT 5.330 958.805 293.095 958.855 ;
        RECT 5.330 956.075 1094.530 958.805 ;
        RECT 5.330 956.025 174.480 956.075 ;
        RECT 5.330 953.365 316.095 953.415 ;
        RECT 5.330 950.635 1094.530 953.365 ;
        RECT 5.330 950.585 157.920 950.635 ;
        RECT 5.330 947.925 243.940 947.975 ;
        RECT 5.330 945.195 1094.530 947.925 ;
        RECT 5.330 945.145 183.615 945.195 ;
        RECT 5.330 942.485 160.680 942.535 ;
        RECT 5.330 939.755 1094.530 942.485 ;
        RECT 5.330 939.705 276.995 939.755 ;
        RECT 5.330 937.045 171.260 937.095 ;
        RECT 5.330 934.315 1094.530 937.045 ;
        RECT 5.330 934.265 33.195 934.315 ;
        RECT 5.330 931.605 20.315 931.655 ;
        RECT 5.330 928.875 1094.530 931.605 ;
        RECT 5.330 928.825 43.775 928.875 ;
        RECT 5.330 926.165 167.515 926.215 ;
        RECT 5.330 923.435 1094.530 926.165 ;
        RECT 5.330 923.385 10.720 923.435 ;
        RECT 5.330 920.725 39.635 920.775 ;
        RECT 5.330 917.995 1094.530 920.725 ;
        RECT 5.330 917.945 41.935 917.995 ;
        RECT 5.330 915.285 39.635 915.335 ;
        RECT 5.330 912.555 1094.530 915.285 ;
        RECT 5.330 912.505 21.760 912.555 ;
        RECT 5.330 909.845 7.895 909.895 ;
        RECT 5.330 907.115 1094.530 909.845 ;
        RECT 5.330 907.065 40.555 907.115 ;
        RECT 5.330 904.405 22.615 904.455 ;
        RECT 5.330 901.675 1094.530 904.405 ;
        RECT 5.330 901.625 78.735 901.675 ;
        RECT 5.330 898.965 39.635 899.015 ;
        RECT 5.330 896.235 1094.530 898.965 ;
        RECT 5.330 896.185 79.720 896.235 ;
        RECT 5.330 893.525 99.435 893.575 ;
        RECT 5.330 890.795 1094.530 893.525 ;
        RECT 5.330 890.745 99.435 890.795 ;
        RECT 5.330 888.085 39.175 888.135 ;
        RECT 5.330 885.355 1094.530 888.085 ;
        RECT 5.330 885.305 209.835 885.355 ;
        RECT 5.330 882.645 191.500 882.695 ;
        RECT 5.330 879.915 1094.530 882.645 ;
        RECT 5.330 879.865 21.300 879.915 ;
        RECT 5.330 877.205 244.400 877.255 ;
        RECT 5.330 874.475 1094.530 877.205 ;
        RECT 5.330 874.425 36.020 874.475 ;
        RECT 5.330 871.765 39.635 871.815 ;
        RECT 5.330 869.035 1094.530 871.765 ;
        RECT 5.330 868.985 90.235 869.035 ;
        RECT 5.330 866.325 56.655 866.375 ;
        RECT 5.330 863.595 1094.530 866.325 ;
        RECT 5.330 863.545 90.235 863.595 ;
        RECT 5.330 860.885 75.055 860.935 ;
        RECT 5.330 858.155 1094.530 860.885 ;
        RECT 5.330 858.105 159.760 858.155 ;
        RECT 5.330 855.445 26.360 855.495 ;
        RECT 5.330 852.715 1094.530 855.445 ;
        RECT 5.330 852.665 43.775 852.715 ;
        RECT 5.330 850.005 49.360 850.055 ;
        RECT 5.330 847.275 1094.530 850.005 ;
        RECT 5.330 847.225 167.975 847.275 ;
        RECT 5.330 844.565 311.035 844.615 ;
        RECT 5.330 841.835 1094.530 844.565 ;
        RECT 5.330 841.785 87.475 841.835 ;
        RECT 5.330 839.125 129.400 839.175 ;
        RECT 5.330 836.395 1094.530 839.125 ;
        RECT 5.330 836.345 85.635 836.395 ;
        RECT 5.330 833.685 196.035 833.735 ;
        RECT 5.330 830.955 1094.530 833.685 ;
        RECT 5.330 830.905 44.300 830.955 ;
        RECT 5.330 828.245 26.820 828.295 ;
        RECT 5.330 825.515 1094.530 828.245 ;
        RECT 5.330 825.465 29.120 825.515 ;
        RECT 5.330 822.805 34.180 822.855 ;
        RECT 5.330 820.075 1094.530 822.805 ;
        RECT 5.330 820.025 37.795 820.075 ;
        RECT 5.330 817.365 429.320 817.415 ;
        RECT 5.330 814.635 1094.530 817.365 ;
        RECT 5.330 814.585 26.295 814.635 ;
        RECT 5.330 811.925 518.495 811.975 ;
        RECT 5.330 809.195 1094.530 811.925 ;
        RECT 5.330 809.145 10.720 809.195 ;
        RECT 5.330 806.485 522.635 806.535 ;
        RECT 5.330 803.755 1094.530 806.485 ;
        RECT 5.330 803.705 41.935 803.755 ;
        RECT 5.330 801.045 151.415 801.095 ;
        RECT 5.330 798.315 1094.530 801.045 ;
        RECT 5.330 798.265 18.080 798.315 ;
        RECT 5.330 795.605 32.275 795.655 ;
        RECT 5.330 792.875 1094.530 795.605 ;
        RECT 5.330 792.825 111.855 792.875 ;
        RECT 5.330 790.165 91.615 790.215 ;
        RECT 5.330 787.435 1094.530 790.165 ;
        RECT 5.330 787.385 8.355 787.435 ;
        RECT 5.330 784.725 133.935 784.775 ;
        RECT 5.330 781.995 1094.530 784.725 ;
        RECT 5.330 781.945 363.015 781.995 ;
        RECT 5.330 779.285 775.700 779.335 ;
        RECT 5.330 776.555 1094.530 779.285 ;
        RECT 5.330 776.505 74.595 776.555 ;
        RECT 5.330 773.845 144.515 773.895 ;
        RECT 5.330 771.115 1094.530 773.845 ;
        RECT 5.330 771.065 76.500 771.115 ;
        RECT 5.330 768.405 46.535 768.455 ;
        RECT 5.330 765.675 1094.530 768.405 ;
        RECT 5.330 765.625 10.720 765.675 ;
        RECT 5.330 762.965 31.355 763.015 ;
        RECT 5.330 760.235 1094.530 762.965 ;
        RECT 5.330 760.185 88.460 760.235 ;
        RECT 5.330 757.525 10.720 757.575 ;
        RECT 5.330 754.795 1094.530 757.525 ;
        RECT 5.330 754.745 470.195 754.795 ;
        RECT 5.330 752.085 128.875 752.135 ;
        RECT 5.330 749.355 1094.530 752.085 ;
        RECT 5.330 749.305 26.295 749.355 ;
        RECT 5.330 746.645 301.835 746.695 ;
        RECT 5.330 743.915 1094.530 746.645 ;
        RECT 5.330 743.865 107.780 743.915 ;
        RECT 5.330 741.205 30.500 741.255 ;
        RECT 5.330 738.475 1094.530 741.205 ;
        RECT 5.330 738.425 128.480 738.475 ;
        RECT 5.330 735.765 131.175 735.815 ;
        RECT 5.330 733.035 1094.530 735.765 ;
        RECT 5.330 732.985 132.620 733.035 ;
        RECT 5.330 730.325 10.720 730.375 ;
        RECT 5.330 727.595 1094.530 730.325 ;
        RECT 5.330 727.545 18.935 727.595 ;
        RECT 5.330 724.885 77.420 724.935 ;
        RECT 5.330 722.155 1094.530 724.885 ;
        RECT 5.330 722.105 7.895 722.155 ;
        RECT 5.330 719.445 83.860 719.495 ;
        RECT 5.330 716.715 1094.530 719.445 ;
        RECT 5.330 716.665 23.140 716.715 ;
        RECT 5.330 714.005 10.720 714.055 ;
        RECT 5.330 711.275 1094.530 714.005 ;
        RECT 5.330 711.225 302.755 711.275 ;
        RECT 5.330 708.565 461.520 708.615 ;
        RECT 5.330 705.835 1094.530 708.565 ;
        RECT 5.330 705.785 489.515 705.835 ;
        RECT 5.330 703.125 31.880 703.175 ;
        RECT 5.330 700.395 1094.530 703.125 ;
        RECT 5.330 700.345 245.780 700.395 ;
        RECT 5.330 697.685 340.935 697.735 ;
        RECT 5.330 694.955 1094.530 697.685 ;
        RECT 5.330 694.905 18.080 694.955 ;
        RECT 5.330 692.245 242.035 692.295 ;
        RECT 5.330 689.515 1094.530 692.245 ;
        RECT 5.330 689.465 273.315 689.515 ;
        RECT 5.330 686.805 294.540 686.855 ;
        RECT 5.330 684.075 1094.530 686.805 ;
        RECT 5.330 684.025 52.515 684.075 ;
        RECT 5.330 681.365 252.220 681.415 ;
        RECT 5.330 678.635 1094.530 681.365 ;
        RECT 5.330 678.585 272.000 678.635 ;
        RECT 5.330 675.925 144.515 675.975 ;
        RECT 5.330 673.195 1094.530 675.925 ;
        RECT 5.330 673.145 44.235 673.195 ;
        RECT 5.330 670.485 26.820 670.535 ;
        RECT 5.330 667.755 1094.530 670.485 ;
        RECT 5.330 667.705 24.455 667.755 ;
        RECT 5.330 665.045 537.815 665.095 ;
        RECT 5.330 662.315 1094.530 665.045 ;
        RECT 5.330 662.265 289.940 662.315 ;
        RECT 5.330 659.605 572.315 659.655 ;
        RECT 5.330 656.875 1094.530 659.605 ;
        RECT 5.330 656.825 121.580 656.875 ;
        RECT 5.330 654.165 135.775 654.215 ;
        RECT 5.330 651.435 1094.530 654.165 ;
        RECT 5.330 651.385 117.440 651.435 ;
        RECT 5.330 648.725 186.375 648.775 ;
        RECT 5.330 645.995 1094.530 648.725 ;
        RECT 5.330 645.945 120.595 645.995 ;
        RECT 5.330 643.285 169.815 643.335 ;
        RECT 5.330 640.555 1094.530 643.285 ;
        RECT 5.330 640.505 100.420 640.555 ;
        RECT 5.330 637.845 126.575 637.895 ;
        RECT 5.330 635.115 1094.530 637.845 ;
        RECT 5.330 635.065 104.100 635.115 ;
        RECT 5.330 632.405 120.200 632.455 ;
        RECT 5.330 629.675 1094.530 632.405 ;
        RECT 5.330 629.625 103.180 629.675 ;
        RECT 5.330 626.965 262.800 627.015 ;
        RECT 5.330 624.235 1094.530 626.965 ;
        RECT 5.330 624.185 142.740 624.235 ;
        RECT 5.330 621.525 140.835 621.575 ;
        RECT 5.330 618.795 1094.530 621.525 ;
        RECT 5.330 618.745 94.835 618.795 ;
        RECT 5.330 616.085 101.800 616.135 ;
        RECT 5.330 613.355 1094.530 616.085 ;
        RECT 5.330 613.305 383.715 613.355 ;
        RECT 5.330 610.645 65.855 610.695 ;
        RECT 5.330 607.915 1094.530 610.645 ;
        RECT 5.330 607.865 50.675 607.915 ;
        RECT 5.330 605.205 49.360 605.255 ;
        RECT 5.330 602.475 1094.530 605.205 ;
        RECT 5.330 602.425 50.740 602.475 ;
        RECT 5.330 599.765 51.660 599.815 ;
        RECT 5.330 597.035 1094.530 599.765 ;
        RECT 5.330 596.985 51.135 597.035 ;
        RECT 5.330 594.325 50.280 594.375 ;
        RECT 5.330 591.595 1094.530 594.325 ;
        RECT 5.330 591.545 69.535 591.595 ;
        RECT 5.330 588.885 50.280 588.935 ;
        RECT 5.330 586.155 1094.530 588.885 ;
        RECT 5.330 586.105 51.200 586.155 ;
        RECT 5.330 583.445 51.200 583.495 ;
        RECT 5.330 580.715 1094.530 583.445 ;
        RECT 5.330 580.665 51.595 580.715 ;
        RECT 5.330 578.005 50.740 578.055 ;
        RECT 5.330 575.275 1094.530 578.005 ;
        RECT 5.330 575.225 52.055 575.275 ;
        RECT 5.330 572.565 130.715 572.615 ;
        RECT 5.330 569.835 1094.530 572.565 ;
        RECT 5.330 569.785 164.295 569.835 ;
        RECT 5.330 567.125 616.475 567.175 ;
        RECT 5.330 564.395 1094.530 567.125 ;
        RECT 5.330 564.345 586.640 564.395 ;
        RECT 5.330 561.685 599.980 561.735 ;
        RECT 5.330 558.955 1094.530 561.685 ;
        RECT 5.330 558.905 97.595 558.955 ;
        RECT 5.330 556.245 82.020 556.295 ;
        RECT 5.330 553.515 1094.530 556.245 ;
        RECT 5.330 553.465 77.880 553.515 ;
        RECT 5.330 550.805 75.580 550.855 ;
        RECT 5.330 548.075 1094.530 550.805 ;
        RECT 5.330 548.025 138.075 548.075 ;
        RECT 5.330 545.365 76.040 545.415 ;
        RECT 5.330 542.635 1094.530 545.365 ;
        RECT 5.330 542.585 78.735 542.635 ;
        RECT 5.330 539.925 244.795 539.975 ;
        RECT 5.330 537.195 1094.530 539.925 ;
        RECT 5.330 537.145 140.835 537.195 ;
        RECT 5.330 534.485 92.075 534.535 ;
        RECT 5.330 531.755 1094.530 534.485 ;
        RECT 5.330 531.705 80.180 531.755 ;
        RECT 5.330 529.045 118.295 529.095 ;
        RECT 5.330 526.315 1094.530 529.045 ;
        RECT 5.330 526.265 80.640 526.315 ;
        RECT 5.330 523.605 154.635 523.655 ;
        RECT 5.330 520.875 1094.530 523.605 ;
        RECT 5.330 520.825 88.460 520.875 ;
        RECT 5.330 518.165 77.420 518.215 ;
        RECT 5.330 515.435 1094.530 518.165 ;
        RECT 5.330 515.385 127.495 515.435 ;
        RECT 5.330 512.725 76.960 512.775 ;
        RECT 5.330 509.995 1094.530 512.725 ;
        RECT 5.330 509.945 92.995 509.995 ;
        RECT 5.330 507.285 248.015 507.335 ;
        RECT 5.330 504.555 1094.530 507.285 ;
        RECT 5.330 504.505 456.460 504.555 ;
        RECT 5.330 501.845 37.400 501.895 ;
        RECT 5.330 499.115 1094.530 501.845 ;
        RECT 5.330 499.065 26.360 499.115 ;
        RECT 5.330 496.405 156.015 496.455 ;
        RECT 5.330 493.675 1094.530 496.405 ;
        RECT 5.330 493.625 366.235 493.675 ;
        RECT 5.330 490.965 27.740 491.015 ;
        RECT 5.330 488.235 1094.530 490.965 ;
        RECT 5.330 488.185 48.900 488.235 ;
        RECT 5.330 485.525 80.575 485.575 ;
        RECT 5.330 482.795 1094.530 485.525 ;
        RECT 5.330 482.745 38.320 482.795 ;
        RECT 5.330 480.085 155.555 480.135 ;
        RECT 5.330 477.355 1094.530 480.085 ;
        RECT 5.330 477.305 164.295 477.355 ;
        RECT 5.330 474.645 157.855 474.695 ;
        RECT 5.330 471.915 1094.530 474.645 ;
        RECT 5.330 471.865 92.995 471.915 ;
        RECT 5.330 469.205 75.580 469.255 ;
        RECT 5.330 466.475 1094.530 469.205 ;
        RECT 5.330 466.425 289.020 466.475 ;
        RECT 5.330 463.765 160.155 463.815 ;
        RECT 5.330 461.035 1094.530 463.765 ;
        RECT 5.330 460.985 145.895 461.035 ;
        RECT 5.330 458.325 234.280 458.375 ;
        RECT 5.330 455.595 1094.530 458.325 ;
        RECT 5.330 455.545 598.535 455.595 ;
        RECT 5.330 452.885 118.295 452.935 ;
        RECT 5.330 450.155 1094.530 452.885 ;
        RECT 5.330 450.105 245.780 450.155 ;
        RECT 5.330 447.445 293.160 447.495 ;
        RECT 5.330 444.715 1094.530 447.445 ;
        RECT 5.330 444.665 22.155 444.715 ;
        RECT 5.330 442.005 49.360 442.055 ;
        RECT 5.330 439.275 1094.530 442.005 ;
        RECT 5.330 439.225 21.300 439.275 ;
        RECT 5.330 436.565 24.520 436.615 ;
        RECT 5.330 433.835 1094.530 436.565 ;
        RECT 5.330 433.785 350.135 433.835 ;
        RECT 5.330 431.125 423.800 431.175 ;
        RECT 5.330 428.395 1094.530 431.125 ;
        RECT 5.330 428.345 24.980 428.395 ;
        RECT 5.330 425.685 21.695 425.735 ;
        RECT 5.330 422.955 1094.530 425.685 ;
        RECT 5.330 422.905 507.455 422.955 ;
        RECT 5.330 420.245 226.000 420.295 ;
        RECT 5.330 417.515 1094.530 420.245 ;
        RECT 5.330 417.465 272.000 417.515 ;
        RECT 5.330 414.805 38.780 414.855 ;
        RECT 5.330 412.075 1094.530 414.805 ;
        RECT 5.330 412.025 26.820 412.075 ;
        RECT 5.330 409.365 223.175 409.415 ;
        RECT 5.330 406.635 1094.530 409.365 ;
        RECT 5.330 406.585 269.175 406.635 ;
        RECT 5.330 403.925 33.720 403.975 ;
        RECT 5.330 401.195 1094.530 403.925 ;
        RECT 5.330 401.145 229.220 401.195 ;
        RECT 5.330 398.485 120.200 398.535 ;
        RECT 5.330 395.755 1094.530 398.485 ;
        RECT 5.330 395.705 144.055 395.755 ;
        RECT 5.330 393.045 74.135 393.095 ;
        RECT 5.330 390.315 1094.530 393.045 ;
        RECT 5.330 390.265 49.755 390.315 ;
        RECT 5.330 387.605 158.775 387.655 ;
        RECT 5.330 384.875 1094.530 387.605 ;
        RECT 5.330 384.825 24.060 384.875 ;
        RECT 5.330 382.165 249.460 382.215 ;
        RECT 5.330 379.435 1094.530 382.165 ;
        RECT 5.330 379.385 28.660 379.435 ;
        RECT 5.330 376.725 110.015 376.775 ;
        RECT 5.330 373.995 1094.530 376.725 ;
        RECT 5.330 373.945 26.820 373.995 ;
        RECT 5.330 371.285 39.635 371.335 ;
        RECT 5.330 368.555 1094.530 371.285 ;
        RECT 5.330 368.505 172.575 368.555 ;
        RECT 5.330 365.845 282.515 365.895 ;
        RECT 5.330 363.115 1094.530 365.845 ;
        RECT 5.330 363.065 154.175 363.115 ;
        RECT 5.330 360.405 38.320 360.455 ;
        RECT 5.330 357.675 1094.530 360.405 ;
        RECT 5.330 357.625 157.395 357.675 ;
        RECT 5.330 354.965 76.895 355.015 ;
        RECT 5.330 352.235 1094.530 354.965 ;
        RECT 5.330 352.185 39.240 352.235 ;
        RECT 5.330 349.525 39.635 349.575 ;
        RECT 5.330 346.795 1094.530 349.525 ;
        RECT 5.330 346.745 124.735 346.795 ;
        RECT 5.330 344.085 121.120 344.135 ;
        RECT 5.330 341.355 1094.530 344.085 ;
        RECT 5.330 341.305 87.475 341.355 ;
        RECT 5.330 338.645 85.635 338.695 ;
        RECT 5.330 335.915 1094.530 338.645 ;
        RECT 5.330 335.865 10.720 335.915 ;
        RECT 5.330 333.205 51.135 333.255 ;
        RECT 5.330 330.475 1094.530 333.205 ;
        RECT 5.330 330.425 157.395 330.475 ;
        RECT 5.330 327.765 485.375 327.815 ;
        RECT 5.330 325.035 1094.530 327.765 ;
        RECT 5.330 324.985 50.675 325.035 ;
        RECT 5.330 322.325 327.595 322.375 ;
        RECT 5.330 319.595 1094.530 322.325 ;
        RECT 5.330 319.545 416.900 319.595 ;
        RECT 5.330 316.885 50.215 316.935 ;
        RECT 5.330 314.155 1094.530 316.885 ;
        RECT 5.330 314.105 10.720 314.155 ;
        RECT 5.330 311.445 24.060 311.495 ;
        RECT 5.330 308.715 1094.530 311.445 ;
        RECT 5.330 308.665 78.735 308.715 ;
        RECT 5.330 306.005 80.115 306.055 ;
        RECT 5.330 303.275 1094.530 306.005 ;
        RECT 5.330 303.225 34.575 303.275 ;
        RECT 5.330 300.565 50.215 300.615 ;
        RECT 5.330 297.785 1094.530 300.565 ;
        RECT 5.330 295.125 417.360 295.175 ;
        RECT 5.330 292.395 1094.530 295.125 ;
        RECT 5.330 292.345 26.360 292.395 ;
        RECT 5.330 289.685 49.295 289.735 ;
        RECT 5.330 286.955 1094.530 289.685 ;
        RECT 5.330 286.905 7.895 286.955 ;
        RECT 5.330 284.245 492.275 284.295 ;
        RECT 5.330 281.515 1094.530 284.245 ;
        RECT 5.330 281.465 33.655 281.515 ;
        RECT 5.330 278.805 275.615 278.855 ;
        RECT 5.330 276.075 1094.530 278.805 ;
        RECT 5.330 276.025 269.175 276.075 ;
        RECT 5.330 273.365 246.635 273.415 ;
        RECT 5.330 270.635 1094.530 273.365 ;
        RECT 5.330 270.585 21.235 270.635 ;
        RECT 5.330 267.925 115.075 267.975 ;
        RECT 5.330 265.195 1094.530 267.925 ;
        RECT 5.330 265.145 76.435 265.195 ;
        RECT 5.330 262.485 125.195 262.535 ;
        RECT 5.330 259.755 1094.530 262.485 ;
        RECT 5.330 259.705 19.000 259.755 ;
        RECT 5.330 257.045 56.655 257.095 ;
        RECT 5.330 254.315 1094.530 257.045 ;
        RECT 5.330 254.265 20.380 254.315 ;
        RECT 5.330 251.605 37.335 251.655 ;
        RECT 5.330 248.875 1094.530 251.605 ;
        RECT 5.330 248.825 18.475 248.875 ;
        RECT 5.330 246.165 73.215 246.215 ;
        RECT 5.330 243.435 1094.530 246.165 ;
        RECT 5.330 243.385 42.395 243.435 ;
        RECT 5.330 240.725 147.340 240.775 ;
        RECT 5.330 237.995 1094.530 240.725 ;
        RECT 5.330 237.945 69.995 237.995 ;
        RECT 5.330 235.285 290.335 235.335 ;
        RECT 5.330 232.555 1094.530 235.285 ;
        RECT 5.330 232.505 272.460 232.555 ;
        RECT 5.330 229.845 146.420 229.895 ;
        RECT 5.330 227.115 1094.530 229.845 ;
        RECT 5.330 227.065 190.515 227.115 ;
        RECT 5.330 224.405 416.440 224.455 ;
        RECT 5.330 221.675 1094.530 224.405 ;
        RECT 5.330 221.625 44.235 221.675 ;
        RECT 5.330 218.965 245.320 219.015 ;
        RECT 5.330 216.235 1094.530 218.965 ;
        RECT 5.330 216.185 146.420 216.235 ;
        RECT 5.330 213.525 343.235 213.575 ;
        RECT 5.330 210.795 1094.530 213.525 ;
        RECT 5.330 210.745 237.960 210.795 ;
        RECT 5.330 208.085 146.880 208.135 ;
        RECT 5.330 205.355 1094.530 208.085 ;
        RECT 5.330 205.305 10.720 205.355 ;
        RECT 5.330 202.645 342.315 202.695 ;
        RECT 5.330 199.915 1094.530 202.645 ;
        RECT 5.330 199.865 27.740 199.915 ;
        RECT 5.330 197.205 57.575 197.255 ;
        RECT 5.330 194.475 1094.530 197.205 ;
        RECT 5.330 194.425 23.140 194.475 ;
        RECT 5.330 191.765 23.140 191.815 ;
        RECT 5.330 189.035 1094.530 191.765 ;
        RECT 5.330 188.985 37.400 189.035 ;
        RECT 5.330 186.325 115.600 186.375 ;
        RECT 5.330 183.595 1094.530 186.325 ;
        RECT 5.330 183.545 297.695 183.595 ;
        RECT 5.330 180.885 178.555 180.935 ;
        RECT 5.330 178.155 1094.530 180.885 ;
        RECT 5.330 178.105 629.420 178.155 ;
        RECT 5.330 175.445 46.535 175.495 ;
        RECT 5.330 172.715 1094.530 175.445 ;
        RECT 5.330 172.665 73.215 172.715 ;
        RECT 5.330 170.005 135.775 170.055 ;
        RECT 5.330 167.275 1094.530 170.005 ;
        RECT 5.330 167.225 116.060 167.275 ;
        RECT 5.330 164.565 117.440 164.615 ;
        RECT 5.330 161.835 1094.530 164.565 ;
        RECT 5.330 161.785 178.555 161.835 ;
        RECT 5.330 159.125 275.155 159.175 ;
        RECT 5.330 156.395 1094.530 159.125 ;
        RECT 5.330 156.345 242.955 156.395 ;
        RECT 5.330 153.685 241.180 153.735 ;
        RECT 5.330 150.955 1094.530 153.685 ;
        RECT 5.330 150.905 19.920 150.955 ;
        RECT 5.330 148.245 49.360 148.295 ;
        RECT 5.330 145.515 1094.530 148.245 ;
        RECT 5.330 145.465 384.700 145.515 ;
        RECT 5.330 142.805 818.415 142.855 ;
        RECT 5.330 140.075 1094.530 142.805 ;
        RECT 5.330 140.025 19.460 140.075 ;
        RECT 5.330 137.365 37.860 137.415 ;
        RECT 5.330 134.635 1094.530 137.365 ;
        RECT 5.330 134.585 50.215 134.635 ;
        RECT 5.330 131.925 81.955 131.975 ;
        RECT 5.330 129.195 1094.530 131.925 ;
        RECT 5.330 129.145 130.320 129.195 ;
        RECT 5.330 126.485 137.220 126.535 ;
        RECT 5.330 123.755 1094.530 126.485 ;
        RECT 5.330 123.705 70.455 123.755 ;
        RECT 5.330 121.045 135.775 121.095 ;
        RECT 5.330 118.315 1094.530 121.045 ;
        RECT 5.330 118.265 36.020 118.315 ;
        RECT 5.330 115.605 226.000 115.655 ;
        RECT 5.330 112.875 1094.530 115.605 ;
        RECT 5.330 112.825 21.760 112.875 ;
        RECT 5.330 110.165 263.260 110.215 ;
        RECT 5.330 107.435 1094.530 110.165 ;
        RECT 5.330 107.385 47.520 107.435 ;
        RECT 5.330 104.725 36.480 104.775 ;
        RECT 5.330 101.995 1094.530 104.725 ;
        RECT 5.330 101.945 74.595 101.995 ;
        RECT 5.330 99.285 7.895 99.335 ;
        RECT 5.330 96.555 1094.530 99.285 ;
        RECT 5.330 96.505 120.200 96.555 ;
        RECT 5.330 93.845 23.600 93.895 ;
        RECT 5.330 91.115 1094.530 93.845 ;
        RECT 5.330 91.065 24.980 91.115 ;
        RECT 5.330 88.405 156.475 88.455 ;
        RECT 5.330 85.675 1094.530 88.405 ;
        RECT 5.330 85.625 125.260 85.675 ;
        RECT 5.330 82.965 119.740 83.015 ;
        RECT 5.330 80.235 1094.530 82.965 ;
        RECT 5.330 80.185 440.820 80.235 ;
        RECT 5.330 77.525 261.815 77.575 ;
        RECT 5.330 74.795 1094.530 77.525 ;
        RECT 5.330 74.745 229.680 74.795 ;
        RECT 5.330 72.085 65.920 72.135 ;
        RECT 5.330 69.355 1094.530 72.085 ;
        RECT 5.330 69.305 24.915 69.355 ;
        RECT 5.330 66.645 139.060 66.695 ;
        RECT 5.330 63.915 1094.530 66.645 ;
        RECT 5.330 63.865 77.355 63.915 ;
        RECT 5.330 61.205 23.140 61.255 ;
        RECT 5.330 58.475 1094.530 61.205 ;
        RECT 5.330 58.425 35.955 58.475 ;
        RECT 5.330 55.765 64.475 55.815 ;
        RECT 5.330 53.035 1094.530 55.765 ;
        RECT 5.330 52.985 150.035 53.035 ;
        RECT 5.330 50.325 120.660 50.375 ;
        RECT 5.330 47.595 1094.530 50.325 ;
        RECT 5.330 47.545 138.075 47.595 ;
        RECT 5.330 44.885 37.335 44.935 ;
        RECT 5.330 42.155 1094.530 44.885 ;
        RECT 5.330 42.105 10.720 42.155 ;
        RECT 5.330 39.445 47.915 39.495 ;
        RECT 5.330 36.715 1094.530 39.445 ;
        RECT 5.330 36.665 36.020 36.715 ;
        RECT 5.330 34.005 344.155 34.055 ;
        RECT 5.330 31.275 1094.530 34.005 ;
        RECT 5.330 31.225 383.255 31.275 ;
        RECT 5.330 28.565 461.980 28.615 ;
        RECT 5.330 25.835 1094.530 28.565 ;
        RECT 5.330 25.785 648.675 25.835 ;
        RECT 5.330 20.345 1094.530 23.175 ;
        RECT 5.330 14.905 1094.530 17.735 ;
        RECT 5.330 10.690 1094.530 12.295 ;
      LAYER li1 ;
        RECT 5.520 10.795 1095.115 1387.285 ;
      LAYER met1 ;
        RECT 5.520 9.900 1095.175 1387.440 ;
      LAYER met2 ;
        RECT 7.090 1395.720 19.590 1396.000 ;
        RECT 20.430 1395.720 33.390 1396.000 ;
        RECT 34.230 1395.720 47.190 1396.000 ;
        RECT 48.030 1395.720 60.990 1396.000 ;
        RECT 61.830 1395.720 74.790 1396.000 ;
        RECT 75.630 1395.720 88.590 1396.000 ;
        RECT 89.430 1395.720 102.390 1396.000 ;
        RECT 103.230 1395.720 116.190 1396.000 ;
        RECT 117.030 1395.720 129.530 1396.000 ;
        RECT 130.370 1395.720 143.330 1396.000 ;
        RECT 144.170 1395.720 157.130 1396.000 ;
        RECT 157.970 1395.720 170.930 1396.000 ;
        RECT 171.770 1395.720 184.730 1396.000 ;
        RECT 185.570 1395.720 198.530 1396.000 ;
        RECT 199.370 1395.720 212.330 1396.000 ;
        RECT 213.170 1395.720 226.130 1396.000 ;
        RECT 226.970 1395.720 239.930 1396.000 ;
        RECT 240.770 1395.720 253.270 1396.000 ;
        RECT 254.110 1395.720 267.070 1396.000 ;
        RECT 267.910 1395.720 280.870 1396.000 ;
        RECT 281.710 1395.720 294.670 1396.000 ;
        RECT 295.510 1395.720 308.470 1396.000 ;
        RECT 309.310 1395.720 322.270 1396.000 ;
        RECT 323.110 1395.720 336.070 1396.000 ;
        RECT 336.910 1395.720 349.870 1396.000 ;
        RECT 350.710 1395.720 363.670 1396.000 ;
        RECT 364.510 1395.720 377.010 1396.000 ;
        RECT 377.850 1395.720 390.810 1396.000 ;
        RECT 391.650 1395.720 404.610 1396.000 ;
        RECT 405.450 1395.720 418.410 1396.000 ;
        RECT 419.250 1395.720 432.210 1396.000 ;
        RECT 433.050 1395.720 446.010 1396.000 ;
        RECT 446.850 1395.720 459.810 1396.000 ;
        RECT 460.650 1395.720 473.610 1396.000 ;
        RECT 474.450 1395.720 487.410 1396.000 ;
        RECT 488.250 1395.720 500.750 1396.000 ;
        RECT 501.590 1395.720 514.550 1396.000 ;
        RECT 515.390 1395.720 528.350 1396.000 ;
        RECT 529.190 1395.720 542.150 1396.000 ;
        RECT 542.990 1395.720 555.950 1396.000 ;
        RECT 556.790 1395.720 569.750 1396.000 ;
        RECT 570.590 1395.720 583.550 1396.000 ;
        RECT 584.390 1395.720 597.350 1396.000 ;
        RECT 598.190 1395.720 611.150 1396.000 ;
        RECT 611.990 1395.720 624.490 1396.000 ;
        RECT 625.330 1395.720 638.290 1396.000 ;
        RECT 639.130 1395.720 652.090 1396.000 ;
        RECT 652.930 1395.720 665.890 1396.000 ;
        RECT 666.730 1395.720 679.690 1396.000 ;
        RECT 680.530 1395.720 693.490 1396.000 ;
        RECT 694.330 1395.720 707.290 1396.000 ;
        RECT 708.130 1395.720 721.090 1396.000 ;
        RECT 721.930 1395.720 734.890 1396.000 ;
        RECT 735.730 1395.720 748.230 1396.000 ;
        RECT 749.070 1395.720 762.030 1396.000 ;
        RECT 762.870 1395.720 775.830 1396.000 ;
        RECT 776.670 1395.720 789.630 1396.000 ;
        RECT 790.470 1395.720 803.430 1396.000 ;
        RECT 804.270 1395.720 817.230 1396.000 ;
        RECT 818.070 1395.720 831.030 1396.000 ;
        RECT 831.870 1395.720 844.830 1396.000 ;
        RECT 845.670 1395.720 858.630 1396.000 ;
        RECT 859.470 1395.720 871.970 1396.000 ;
        RECT 872.810 1395.720 885.770 1396.000 ;
        RECT 886.610 1395.720 899.570 1396.000 ;
        RECT 900.410 1395.720 913.370 1396.000 ;
        RECT 914.210 1395.720 927.170 1396.000 ;
        RECT 928.010 1395.720 940.970 1396.000 ;
        RECT 941.810 1395.720 954.770 1396.000 ;
        RECT 955.610 1395.720 968.570 1396.000 ;
        RECT 969.410 1395.720 982.370 1396.000 ;
        RECT 983.210 1395.720 995.710 1396.000 ;
        RECT 996.550 1395.720 1009.510 1396.000 ;
        RECT 1010.350 1395.720 1023.310 1396.000 ;
        RECT 1024.150 1395.720 1037.110 1396.000 ;
        RECT 1037.950 1395.720 1050.910 1396.000 ;
        RECT 1051.750 1395.720 1064.710 1396.000 ;
        RECT 1065.550 1395.720 1078.510 1396.000 ;
        RECT 1079.350 1395.720 1092.310 1396.000 ;
        RECT 1093.150 1395.720 1093.330 1396.000 ;
        RECT 6.530 9.870 1093.330 1395.720 ;
      LAYER met3 ;
        RECT 6.505 10.715 1093.355 1387.365 ;
      LAYER met4 ;
        RECT 14.095 26.695 20.640 1380.905 ;
        RECT 23.040 26.695 97.440 1380.905 ;
        RECT 99.840 26.695 174.240 1380.905 ;
        RECT 176.640 26.695 251.040 1380.905 ;
        RECT 253.440 26.695 327.840 1380.905 ;
        RECT 330.240 26.695 404.640 1380.905 ;
        RECT 407.040 26.695 481.440 1380.905 ;
        RECT 483.840 26.695 558.240 1380.905 ;
        RECT 560.640 26.695 635.040 1380.905 ;
        RECT 637.440 26.695 711.840 1380.905 ;
        RECT 714.240 26.695 788.640 1380.905 ;
        RECT 791.040 26.695 865.440 1380.905 ;
        RECT 867.840 26.695 942.240 1380.905 ;
        RECT 944.640 26.695 1019.040 1380.905 ;
        RECT 1021.440 26.695 1064.145 1380.905 ;
  END
END DFFRAM_1Kx32
END LIBRARY

